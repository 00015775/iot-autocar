PK
     `+�[ީ���|  �|     cirkitFile.json{"raven_core_version":15,"hardware_version":0,"pin_to_graph":{"pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_0_0":[],"pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_0":["pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_24"],"pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_0_1":[],"pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_1":["pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_23"],"pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_0_2":[],"pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_2":["pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_27"],"pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_0_3":[],"pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_3":["pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_28"],"pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_0_4":[],"pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_4":["pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_10"],"pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_0_5":[],"pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_5":[],"pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_0_6":[],"pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_6":[],"pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_0_7":[],"pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_7":[],"pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_0_8":[],"pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_8":[],"pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_0_9":[],"pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_9":[],"pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_0_10":[],"pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_10":[],"pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_0_11":[],"pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_11":[],"pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_0_12":[],"pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_12":[],"pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_0_13":[],"pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_13":[],"pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_0_14":[],"pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_14":[],"pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_0_15":[],"pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_15":[],"pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_0_16":[],"pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_16":[],"pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_0":[],"pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_1":[],"pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_2":[],"pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_3":[],"pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_4":[],"pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_5":[],"pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_6":[],"pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_7":[],"pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_8":[],"pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_9":[],"pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_10":["pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_4"],"pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_11":[],"pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_12":[],"pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_13":[],"pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_14":[],"pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_15":[],"pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_16":[],"pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_17":[],"pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_18":[],"pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_19":[],"pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_20":[],"pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_21":[],"pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_22":[],"pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_23":["pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_1"],"pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_24":["pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_0"],"pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_25":[],"pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_26":[],"pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_27":["pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_2"],"pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_28":["pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_3"],"pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_29":[],"pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_30":[],"pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_31":[],"pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_32":[],"pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_33":[],"pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_34":[],"pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_35":[],"pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_36":[],"pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_37":[],"pin-type-component_0767d6d7-c92e-4635-8656-1d8c21f3772f_0":[],"pin-type-component_0767d6d7-c92e-4635-8656-1d8c21f3772f_1":[],"pin-type-component_0767d6d7-c92e-4635-8656-1d8c21f3772f_2":[],"pin-type-component_0767d6d7-c92e-4635-8656-1d8c21f3772f_3":[],"pin-type-component_0767d6d7-c92e-4635-8656-1d8c21f3772f_4":[]},"pin_to_color":{"pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_0_0":"#000000","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_0":"#010067","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_0_1":"#000000","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_1":"#ff2600","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_0_2":"#000000","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_2":"#0061ff","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_0_3":"#000000","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_3":"#77bb41","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_0_4":"#000000","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_4":"#a800ec","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_0_5":"#000000","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_5":"#000000","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_0_6":"#000000","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_6":"#000000","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_0_7":"#000000","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_7":"#000000","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_0_8":"#000000","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_8":"#000000","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_0_9":"#000000","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_9":"#000000","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_0_10":"#000000","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_10":"#000000","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_0_11":"#000000","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_11":"#000000","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_0_12":"#000000","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_12":"#000000","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_0_13":"#000000","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_13":"#000000","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_0_14":"#000000","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_14":"#000000","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_0_15":"#000000","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_15":"#000000","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_0_16":"#000000","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_16":"#000000","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_0":"#000000","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_1":"#000000","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_2":"#000000","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_3":"#000000","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_4":"#000000","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_5":"#000000","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_6":"#000000","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_7":"#000000","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_8":"#000000","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_9":"#000000","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_10":"#a800ec","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_11":"#000000","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_12":"#000000","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_13":"#000000","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_14":"#000000","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_15":"#000000","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_16":"#000000","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_17":"#000000","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_18":"#000000","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_19":"#000000","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_20":"#000000","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_21":"#000000","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_22":"#000000","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_23":"#ff2600","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_24":"#010067","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_25":"#000000","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_26":"#000000","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_27":"#0061ff","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_28":"#77bb41","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_29":"#000000","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_30":"#000000","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_31":"#000000","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_32":"#000000","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_33":"#000000","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_34":"#000000","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_35":"#000000","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_36":"#000000","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_37":"#000000","pin-type-component_0767d6d7-c92e-4635-8656-1d8c21f3772f_0":"#000000","pin-type-component_0767d6d7-c92e-4635-8656-1d8c21f3772f_1":"#000000","pin-type-component_0767d6d7-c92e-4635-8656-1d8c21f3772f_2":"#000000","pin-type-component_0767d6d7-c92e-4635-8656-1d8c21f3772f_3":"#000000","pin-type-component_0767d6d7-c92e-4635-8656-1d8c21f3772f_4":"#000000"},"pin_to_state":{"pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_0_0":"neutral","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_0":"neutral","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_0_1":"neutral","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_1":"neutral","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_0_2":"neutral","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_2":"neutral","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_0_3":"neutral","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_3":"neutral","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_0_4":"neutral","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_4":"neutral","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_0_5":"neutral","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_5":"neutral","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_0_6":"neutral","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_6":"neutral","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_0_7":"neutral","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_7":"neutral","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_0_8":"neutral","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_8":"neutral","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_0_9":"neutral","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_9":"neutral","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_0_10":"neutral","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_10":"neutral","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_0_11":"neutral","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_11":"neutral","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_0_12":"neutral","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_12":"neutral","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_0_13":"neutral","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_13":"neutral","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_0_14":"neutral","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_14":"neutral","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_0_15":"neutral","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_15":"neutral","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_0_16":"neutral","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_16":"neutral","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_0":"neutral","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_1":"neutral","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_2":"neutral","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_3":"neutral","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_4":"neutral","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_5":"neutral","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_6":"neutral","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_7":"neutral","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_8":"neutral","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_9":"neutral","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_10":"neutral","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_11":"neutral","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_12":"neutral","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_13":"neutral","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_14":"neutral","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_15":"neutral","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_16":"neutral","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_17":"neutral","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_18":"neutral","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_19":"neutral","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_20":"neutral","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_21":"neutral","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_22":"neutral","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_23":"neutral","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_24":"neutral","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_25":"neutral","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_26":"neutral","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_27":"neutral","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_28":"neutral","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_29":"neutral","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_30":"neutral","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_31":"neutral","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_32":"neutral","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_33":"neutral","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_34":"neutral","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_35":"neutral","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_36":"neutral","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_37":"neutral","pin-type-component_0767d6d7-c92e-4635-8656-1d8c21f3772f_0":"neutral","pin-type-component_0767d6d7-c92e-4635-8656-1d8c21f3772f_1":"neutral","pin-type-component_0767d6d7-c92e-4635-8656-1d8c21f3772f_2":"neutral","pin-type-component_0767d6d7-c92e-4635-8656-1d8c21f3772f_3":"neutral","pin-type-component_0767d6d7-c92e-4635-8656-1d8c21f3772f_4":"neutral"},"next_color_idx":5,"wires_placed_in_order":[["pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_0","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_24"],["pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_1","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_23"],["pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_2","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_27"],["pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_3","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_28"],["pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_4","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_10"]],"wires_removed_and_placed_in_order":[[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[["pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_0","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_24"]]],[[],[["pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_1","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_23"]]],[[],[["pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_2","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_27"]]],[[],[["pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_3","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_28"]]],[[],[["pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_4","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_10"]]]],"arduino_state":"arduino_off","pin_to_uid":{"pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_0_0":"_","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_0":"0000000000000000","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_0_1":"_","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_1":"0000000000000001","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_0_2":"_","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_2":"0000000000000002","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_0_3":"_","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_3":"0000000000000003","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_0_4":"_","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_4":"0000000000000004","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_0_5":"_","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_5":"_","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_0_6":"_","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_6":"_","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_0_7":"_","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_7":"_","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_0_8":"_","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_8":"_","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_0_9":"_","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_9":"_","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_0_10":"_","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_10":"_","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_0_11":"_","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_11":"_","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_0_12":"_","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_12":"_","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_0_13":"_","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_13":"_","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_0_14":"_","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_14":"_","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_0_15":"_","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_15":"_","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_0_16":"_","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_16":"_","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_0":"_","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_1":"_","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_2":"_","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_3":"_","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_4":"_","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_5":"_","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_6":"_","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_7":"_","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_8":"_","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_9":"_","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_10":"0000000000000004","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_11":"_","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_12":"_","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_13":"_","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_14":"_","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_15":"_","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_16":"_","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_17":"_","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_18":"_","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_19":"_","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_20":"_","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_21":"_","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_22":"_","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_23":"0000000000000001","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_24":"0000000000000000","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_25":"_","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_26":"_","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_27":"0000000000000002","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_28":"0000000000000003","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_29":"_","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_30":"_","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_31":"_","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_32":"_","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_33":"_","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_34":"_","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_35":"_","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_36":"_","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_37":"_","pin-type-component_0767d6d7-c92e-4635-8656-1d8c21f3772f_0":"_","pin-type-component_0767d6d7-c92e-4635-8656-1d8c21f3772f_1":"_","pin-type-component_0767d6d7-c92e-4635-8656-1d8c21f3772f_2":"_","pin-type-component_0767d6d7-c92e-4635-8656-1d8c21f3772f_3":"_","pin-type-component_0767d6d7-c92e-4635-8656-1d8c21f3772f_4":"_"},"component_id_to_pins":{"bc8378c5-ac3f-4da3-b662-1e1cdc615429":["0","1","2","3","4","5","6","7","8","9","10","11","12","13","14","15","16","17","18","19","20","21","22","23","24","25","26","27","28","29","30","31","32","33","34","35","36","37"],"0767d6d7-c92e-4635-8656-1d8c21f3772f":["0","1","2","3","4"],"b66c2a17-0752-4593-99ab-d606efa4d77d":[]},"uid_to_net":{"_":[],"0000000000000000":["pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_0","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_24"],"0000000000000001":["pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_1","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_23"],"0000000000000002":["pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_2","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_27"],"0000000000000003":["pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_3","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_28"],"0000000000000004":["pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_4","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_10"]},"uid_to_text_label":{"0000000000000000":"Net 0","0000000000000001":"Net 1","0000000000000002":"Net 2","0000000000000003":"Net 3","0000000000000004":"Net 4"},"all_breadboard_info_list":["0eae91f8-3d4b-4e59-8923-87a6d2900cd0_17_2_False_1195_280_up"],"breadboard_info_list":["0eae91f8-3d4b-4e59-8923-87a6d2900cd0_17_2_False_1195_280_up"],"componentsData":[{"compProperties":{"mpn":{"version":2,"id":"mpn","label":"mpn","description":"","units":"","type":"string","value":"DEV-13850","displayFormat":"input","showOnComp":false,"isVisibleToUser":false},"manufacturer":{"version":2,"id":"manufacturer","label":"manufacturer","description":"","units":"","type":"string","value":"SparkFun","displayFormat":"input","showOnComp":false,"isVisibleToUser":false}},"position":[800.38168,417.0763505],"typeId":"11b06032-2d2c-49c8-bde9-6a809e00e513","componentVersion":1,"instanceId":"bc8378c5-ac3f-4da3-b662-1e1cdc615429","orientation":"up","circleData":[[992.5,560],[727.8524695000001,274.3795805],[742.8200995,274.41025849999994],[757.8853374999999,274.390736],[772.8585444999999,274.40816599999994],[787.9349379999999,274.3935245],[802.9240585,274.4018915],[817.9511184999999,274.40747],[833.0032510000001,274.41025849999994],[848.046214,274.40747],[863.098444,274.413047],[887.289655,274.398008],[902.318638,274.39422199999996],[917.3476209999999,274.3935245],[932.3259009999999,274.39910299999997],[947.3580549999999,274.40747],[962.3991894999999,274.41025849999994],[977.4525715,274.41025849999994],[992.5043304999999,274.40747],[782.1481239999998,559.9470125],[797.1743185,559.9609565],[812.200513,559.991633],[827.2294975,559.991633],[842.2110700000001,559.980479],[857.2484199999999,560.0055785],[872.2506145,560.0055785],[887.2450329999999,559.9409315],[917.3755105,559.9619135],[932.4044935,559.9776889999999],[947.376694,559.9470125],[962.42128,559.9330685],[977.4518665,560],[993.340342,394.067633],[1008.3944259999998,394.0425335],[993.3375535,409.091039],[1008.400003,409.085462],[993.340342,424.12839049999997],[1008.3721150000001,424.1702225]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[1387.9405150000002,322.5251404999999],"typeId":"69390a6c-c81c-fde0-536a-a1b73720f902","componentVersion":1,"instanceId":"0767d6d7-c92e-4635-8656-1d8c21f3772f","orientation":"right","circleData":[[1292.5,290],[1292.5000060000002,304.8744019999999],[1292.5000060000002,319.7488025],[1292.5,334.62322849999987],[1292.5,349.4976244999998]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"Comment":{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"HW-504 2-Axis joystick:\n    GND - GND\n    5V+ - 5V\n    VRx - A0 (only analog pin)\n    VRy - A1 (only analog pin)\n    SW - digital pin 8","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"backgroundColor":{"version":2,"id":"backgroundColor","label":"Background Color","description":"","units":"","type":"string","value":"#d6d6d6","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"backgroundOpacity":{"version":2,"id":"backgroundOpacity","label":"Background Opacity","description":"","units":"","type":"decimal","value":"1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"textColor":{"version":2,"id":"textColor","label":"Text Color","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"fontSize":{"version":2,"id":"fontSize","label":"Font Size","description":"","units":"","type":"integer","value":"12","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"font":{"version":2,"id":"font","label":"Font","description":"","units":"","type":"string","value":"Arial","displayFormat":"input","showOnComp":false,"isVisibleToUser":true}},"position":[1465.994140625,488.4],"typeId":"9a5a4baa-44d4-4aa0-8d82-488487322b20","componentVersion":1,"instanceId":"b66c2a17-0752-4593-99ab-d606efa4d77d","orientation":"up","circleData":[],"cirkitStudioVersion":"1.3.3"}],"bounds":{"top":"242.97084","left":"569.23593","width":"987.76407","height":"341.87866","x":"569.23593","y":"242.97084"},"cachedBreadboardPrettyViewWires":["{\"color\":\"#010067\",\"startPinId\":\"pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_0\",\"endPinId\":\"pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_24\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_0_0\",\"rawEndPinId\":\"pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_24\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1262.5000000000_290.0000000000\\\",\\\"1262.5000000000_260.0000000000\\\",\\\"1097.5000000000_260.0000000000\\\",\\\"1097.5000000000_627.5000000000\\\",\\\"857.2484200000_627.5000000000\\\",\\\"857.2484200000_560.0055785000\\\"]}\"}","{\"color\":\"#ff2600\",\"startPinId\":\"pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_1\",\"endPinId\":\"pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_23\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_1_0\",\"rawEndPinId\":\"pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_23\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1262.5000000000_305.0000000000\\\",\\\"1255.0000000000_305.0000000000\\\",\\\"1255.0000000000_275.0000000000\\\",\\\"1112.5000000000_275.0000000000\\\",\\\"1112.5000000000_642.5000000000\\\",\\\"842.2110700000_642.5000000000\\\",\\\"842.2110700000_559.9804790000\\\"]}\"}","{\"color\":\"#0061ff\",\"startPinId\":\"pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_2\",\"endPinId\":\"pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_27\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_2_0\",\"rawEndPinId\":\"pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_27\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1262.5000000000_320.0000000000\\\",\\\"1240.0000000000_320.0000000000\\\",\\\"1240.0000000000_612.5000000000\\\",\\\"917.3755105000_612.5000000000\\\",\\\"917.3755105000_559.9619135000\\\"]}\"}","{\"color\":\"#77bb41\",\"startPinId\":\"pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_3\",\"endPinId\":\"pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_28\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_3_0\",\"rawEndPinId\":\"pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_28\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1262.5000000000_335.0000000000\\\",\\\"1255.0000000000_335.0000000000\\\",\\\"1255.0000000000_597.5000000000\\\",\\\"932.4044935000_597.5000000000\\\",\\\"932.4044935000_559.9776890000\\\"]}\"}","{\"color\":\"#a800ec\",\"startPinId\":\"pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_4\",\"endPinId\":\"pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_10\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_4_0\",\"rawEndPinId\":\"pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_10\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1262.5000000000_350.0000000000\\\",\\\"1270.0000000000_350.0000000000\\\",\\\"1270.0000000000_410.0000000000\\\",\\\"1517.5000000000_410.0000000000\\\",\\\"1517.5000000000_230.0000000000\\\",\\\"863.0984440000_230.0000000000\\\",\\\"863.0984440000_274.4130470000\\\"]}\"}"],"projectDescription":""}PK
     `+�[               jsons/PK
     `+�[�rՍ�  �     jsons/user_defined.json{"type":"user_defined","version":"0.0.1","subtypes":[{"subtypeName":"Arduino 101","category":["User Defined"],"userDefined":true,"id":"11b06032-2d2c-49c8-bde9-6a809e00e513","subtypeDescription":"","subtypePic":"c7631ad6-ed21-46e6-964c-e953ba5165ac.png","pinInfo":{"numDisplayCols":"29.48610","numDisplayRows":"21.03642","pins":[{"uniquePinIdString":"0","positionMil":"2755.09380,98.99667","isAnchorPin":true,"label":"A5/SCL"},{"uniquePinIdString":"1","positionMil":"990.77693,2003.13280","isAnchorPin":false,"label":"A5/SCL"},{"uniquePinIdString":"2","positionMil":"1090.56113,2002.92828","isAnchorPin":false,"label":"A4/SDA"},{"uniquePinIdString":"3","positionMil":"1190.99605,2003.05843","isAnchorPin":false,"label":"AREF"},{"uniquePinIdString":"4","positionMil":"1290.81743,2002.94223","isAnchorPin":false,"label":"GND"},{"uniquePinIdString":"5","positionMil":"1391.32672,2003.03984","isAnchorPin":false,"label":"D13/SCK"},{"uniquePinIdString":"6","positionMil":"1491.25419,2002.98406","isAnchorPin":false,"label":"D12/MISO"},{"uniquePinIdString":"7","positionMil":"1591.43459,2002.94687","isAnchorPin":false,"label":"D11 PWM/MOSI"},{"uniquePinIdString":"8","positionMil":"1691.78214,2002.92828","isAnchorPin":false,"label":"D10 PWM/SS"},{"uniquePinIdString":"9","positionMil":"1792.06856,2002.94687","isAnchorPin":false,"label":"D9 PWM"},{"uniquePinIdString":"10","positionMil":"1892.41676,2002.90969","isAnchorPin":false,"label":"D8"},{"uniquePinIdString":"11","positionMil":"2053.69150,2003.00995","isAnchorPin":false,"label":"D7"},{"uniquePinIdString":"12","positionMil":"2153.88472,2003.03519","isAnchorPin":false,"label":"D6 PWM"},{"uniquePinIdString":"13","positionMil":"2254.07794,2003.03984","isAnchorPin":false,"label":"D5 PWM"},{"uniquePinIdString":"14","positionMil":"2353.93314,2003.00265","isAnchorPin":false,"label":"D4"},{"uniquePinIdString":"15","positionMil":"2454.14750,2002.94687","isAnchorPin":false,"label":"D3 PWM"},{"uniquePinIdString":"16","positionMil":"2554.42173,2002.92828","isAnchorPin":false,"label":"D2"},{"uniquePinIdString":"17","positionMil":"2654.77761,2002.92828","isAnchorPin":false,"label":"D1/TX"},{"uniquePinIdString":"18","positionMil":"2755.12267,2002.94687","isAnchorPin":false,"label":"D0/RX"},{"uniquePinIdString":"19","positionMil":"1352.74796,99.34992","isAnchorPin":false,"label":"AIN"},{"uniquePinIdString":"20","positionMil":"1452.92259,99.25696","isAnchorPin":false,"label":"ioref"},{"uniquePinIdString":"21","positionMil":"1553.09722,99.05245","isAnchorPin":false,"label":"RESET"},{"uniquePinIdString":"22","positionMil":"1653.29045,99.05245","isAnchorPin":false,"label":"3V3"},{"uniquePinIdString":"23","positionMil":"1753.16760,99.12681","isAnchorPin":false,"label":"5V"},{"uniquePinIdString":"24","positionMil":"1853.41660,98.95948","isAnchorPin":false,"label":"GND"},{"uniquePinIdString":"25","positionMil":"1953.43123,98.95948","isAnchorPin":false,"label":"GND"},{"uniquePinIdString":"26","positionMil":"2053.39402,99.39046","isAnchorPin":false,"label":"VIN"},{"uniquePinIdString":"27","positionMil":"2254.26387,99.25058","isAnchorPin":false,"label":"A0"},{"uniquePinIdString":"28","positionMil":"2354.45709,99.14541","isAnchorPin":false,"label":"A1"},{"uniquePinIdString":"29","positionMil":"2454.27176,99.34992","isAnchorPin":false,"label":"A2"},{"uniquePinIdString":"30","positionMil":"2554.56900,99.44288","isAnchorPin":false,"label":"A3"},{"uniquePinIdString":"31","positionMil":"2654.77291,98.99667","isAnchorPin":false,"label":"A4/SDA"},{"uniquePinIdString":"32","positionMil":"2760.69608,1205.21245","isAnchorPin":false,"label":"ICSP MISO"},{"uniquePinIdString":"33","positionMil":"2861.05664,1205.37978","isAnchorPin":false,"label":"5V"},{"uniquePinIdString":"34","positionMil":"2760.67749,1105.05641","isAnchorPin":false,"label":"ICSP SCK"},{"uniquePinIdString":"35","positionMil":"2861.09382,1105.09359","isAnchorPin":false,"label":"ICSP MOSI"},{"uniquePinIdString":"36","positionMil":"2760.69608,1004.80740","isAnchorPin":false,"label":"RESET"},{"uniquePinIdString":"37","positionMil":"2860.90790,1004.52852","isAnchorPin":false,"label":"GND"}],"pinType":"wired"},"properties":[{"type":"string","name":"mpn","value":"DEV-13850","unit":"","showOnComp":false,"userVisible":false,"required":true},{"type":"string","name":"manufacturer","value":"SparkFun","unit":"","showOnComp":false,"userVisible":false,"required":true}],"iconPic":"97fe1122-b934-4e82-b9ff-450ac31bc7af.png","componentVersion":1,"imageLocation":"local_cache","hasComponentImageSvg":false,"componentImageSvgUrl":""},{"subtypeName":"KY-023 Dual Axis Joystick Module","category":["Input"],"userDefined":true,"id":"69390a6c-c81c-fde0-536a-a1b73720f902","subtypeDescription":"","subtypePic":"d5d3b89f-59ab-4c38-95f7-2948dd30f8f5.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"10.60724","numDisplayRows":"15.77946","pins":[{"uniquePinIdString":"0","positionMil":"313.52773,152.70290","isAnchorPin":true,"label":"GND"},{"uniquePinIdString":"1","positionMil":"412.69041,152.70294","isAnchorPin":false,"label":"+5V"},{"uniquePinIdString":"2","positionMil":"511.85308,152.70294","isAnchorPin":false,"label":"VRx"},{"uniquePinIdString":"3","positionMil":"611.01592,152.70290","isAnchorPin":false,"label":"VRy"},{"uniquePinIdString":"4","positionMil":"710.17856,152.70290","isAnchorPin":false,"label":"SW"}],"pinType":"wired"},"properties":[],"iconPic":"60da03ea-f7cc-456a-983c-41a209708cd9.png","componentVersion":1,"hasComponentImageSvg":false,"componentImageSvgUrl":""},{"subtypeName":"Comment V2","category":["User Defined"],"componentClass":"textbox","userDefined":true,"id":"9a5a4baa-44d4-4aa0-8d82-488487322b20","subtypeDescription":"","subtypePic":"c88b2895-5e8b-4a57-9f9a-b80dd50058b1.png","pinInfo":{"numPins":"0","polarity":[],"pinType":"movable"},"properties":[{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"text box (click to edit)","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"backgroundColor","label":"Background Color","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"backgroundOpacity","label":"Background Opacity","description":"","units":"","type":"decimal","value":"1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"textColor","label":"Text Color","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"fontSize","label":"Font Size","description":"","units":"","type":"integer","value":"10","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"font","label":"Font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true}],"iconPic":"d3694a2e-5bba-40c3-8069-8db85c4c9209.png","componentVersion":1,"imageLocation":"local_cache","propertiesV2":[],"hasComponentImageSvg":false,"componentImageSvgUrl":""}]}PK
     `+�[               images/PK
     `+�[�:��� �� /   images/c7631ad6-ed21-46e6-964c-e953ba5165ac.png�PNG

   IHDR  �  .   ���   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  ��IDATx���[Օ��{Ouf4�t{�q�b��`L3�w 		ٰ!��dI�)N6�KB�&�,��lXj�	�L�c6.���i*�ьFS,��+z:�D�F�<������s]@Y��m�uM��$I���K
Aa[6��+���<����{�ߞ\�� � �0��-Q�b��YC�;�+W���*.�%�F�`����@AAAA����z��֕�^ +��"+Hp'K��-������ � �]�O/��AAA�����pۓ%7�zޞ�n�"cHp'���;�en���w�o2A����NAA��H��e�٪o��Y������ ������� [��� � �� � � F�tB�H�{�7��l�3�wb ��63���( � �����	� � �ztX�ϖ_{�Mw]�İ��N�#�Il'� �A�5AAA#G��4�\zí���vcCB�;�K���&�����CA�(R� � � ,�e�3��o[�r�-@
	�g����e�Q �� � �N�AAA��]Q�)����^fpHp'8��߁H%� �B�;AAAB� �U=�l�����9D?Hp' t�(�_AA8M�$�C4��AAaG�cq\�?U��g�[��N z!�� ]�_I:(@X���Z�e�nlV��c��)C�˧��W�U���Žo�t4���$� ���s)&IR$�{�5?$�n �7�%),�J�R�����ݭ�q��X��J�rIh��+A�͐I�&� � B,:,�G�{í����. 8$�8���648�л:v��v�P(ZW�Xе���Y����/$_�z����zHW㉧j �Z{[��C��	�fH���|mri�g��e�O�Q�����X�Q$�a�8^�KN{ǚ���;�l_AEO�������AAQH��!�����+����BG�\����ͭ*�$�sh�~�K-r)q3�!�UT���~�.����Kmon�����z���StM�&���ޑ|�.A��Kj�k@L)��>U�}M�؝z�� vAI�}:ƷC"ڞ���c������G{;�KK^��Ӧ�?
��9q\Շw��A&{� � � l[l��Ï��\y!�\���B撇\y�ʥ3��^ב`{�ᢅ3���+�����]��c��]%�px��i��%�>�K'���dN�~�[��������ݮ���뮮���弸O� � � � �rV0\�x�w^ w]�u�c'A�{S6�౺���DT-yD��8n�1G�G�k�h�㳝�v�ܽ����1��ڪ57���p�2@wwĭi��|��펻�.5�ڊ�h^�Ǵ�~�OS\�.ĥ(zIQQ�
ĬY��P�1�'�$�
� L��=�k�OAA��pFȫ�ײr奰r�)�'�	���j�%)�s�FT-����)�1u�L� �X;(������Z��q+2�//��� ����s���rA[w�=�����Z����k!�$�N�5AAA&�K������\��B�Ip/`$I:�x\���bo���N�mHm�N�:N�2M��q�p��a����6l�����?��~H^m�!qH)�AAA������h�%}	�\�iw$�6c!ω��i)TgS�no��L����¹s'����#�Fy���X�ן�"q^�t'������ۡ+V��v�@�w� � � �D��/�����\y%�\YP�	��R@��^�wFՂj��q�-�w a)�$�(���·�fN ���.�<b�G�p�{�U��ޖv ��kz~�#� � "���K�p9��_/$ѝ�F��9lN{��v�11XD�F,���f��0��J�������ų��5���Ͻ���B8�3��3''� � ��ղpE���
#�%	����ռ=��=B�~ә1�n��DX2i�%��Q��#������W���A8]�S�Z�h�'� � �<G��B7�%�ܢ�S!��$�yMgL��(}�T�=t`��ࡧ�Z� ��bO�b5�^7����������� ���py�b'� � "Ϲ*t�]�-���;]t'���k±8	�w%�0&T�}�p��Q`7�ה���^�x�m�㕵@�LN��2AAA�#�u�����V^���$�yM{D�:L�%K�d	TM�í̲�up�e+���vŭ�<����*����;� � � � rG�겶r�y�ʫ�*��XY�����<��� ��.��=��&�xpɑ��?>*���O��A�ܟ����.aוu=:y�+� �5���t)?����O7EF���
yƦ�����yw߅���ARi�aA��Җܖ�tťk�˒s4م���y��V�L]Q�v�v��ӝx�<�'�qf�|����y����p���Icm�a%��Q �(d$�ƕ�R���*�tx�AVc��<l��h*�G>$�1I���5d�]}Қ�xؘ���l���>|�?U6nD|b���|=.w�\��U���w�	��y������L��w�|���A���m�-@"�nɌ�qM��fk9V��"�Ӌ<�*)��]����^Eq�e�_4�[��.Ev�k�h>�^�lqeG���y��󖂜g�.���'�� ���Ǡ^���t�w�,�0��m`'�'A ��OtI�w�f�e�_n�P�^ � �Ŀ~�y���|%8u��/�ʕ��ZN�{!#Ys��GV�E�#E\˧�j{+�ΛYp�\��z�1�ś����ų�W� y���2sT<q�p��Ǝ�Ewo������A�tt����s AA�5[���"���P�����;/�����C ���k$9_%<�bj��nQ$������RQt��/���q������E�h�KA����{wA�H|��P���s�^��֕�^+��@����̗H,�����+�y./�a�*���)~��&���.>����9]���N	P	� �0�p'� D���K�~fY8�x��^����f$�2�*	�H�$����R�`1T�����<|ng3�=^߶X3�Al�K�AA����Ys�tA�Ÿb��� +�e���y��8K	!�aB�,Q�;!M�D��<�S�å�aLH���v�ѿ�e�km�߻#�n � ��X���HA� �(\���i�u���BƢCSE�k:	�0t�|"�#Y���j�8�8e�xp*A���d���'G���R�� � ��s̹sA������4;,8B�#��0��$�"�(�=Gj�%�s��s��ܩ�Ҧ�Y�����w�MvR�ti|�3�'7e��K2!,O��ޟ�>���C�}.�}ݾd��R�c0�4Mg��z����XlS&e�v x�鷛^���g8[���J�<�_�+'��I��pm<Y.H�z6�ږZ������P����֖�^�2����3��l�}���J�����Pm��LD��-�p�s?2f��M�zD�������|�U���j���Dz�������2���|�ӹ]���$��SΖ�s�$Ґea[���Sǵ�����F�Õ��,;����_��d�yS�����k�s�\�E�w�d@�;�װ�"�c�	[���T�l�`l?>s	|(~r�x��]���uC���3y_WW'�����N�[����`�Lؤ2�A8�v���?u]l��.�&'��`E̜-�CGG;��'�M�gҮR6�6����3uC[��Z{ʡ��E��(�>A�^�����\m	�[{�U�a$h������\�mhmmU��A����C��SLЖp��wA�l3F��T�<JKC��������6��{�b�(;Rی���bq)�Plliifu,!:i�X�'��6�uM$I[�"�mɸ��֝7%k��އ�Z4�i��.��@��~���#��߸ �>QT�c޿���Vq�ݍi��ۂY6h����u\�H��M{oK��F�1����/�D"ݼ�!f�kɶ��PH�#�� b���
ڀ���ChK{{��u�J2>'���hOYYEf"����w��6��䄄0�0��~�1"揭�������+�ܹ����f�w�Lއ�P\4�"1c��4��"�P\.7[�yق>F���&����v;�8Hu�Ij$.|E��^������FӷHH��n�O�؎�->_���	£���`���f��YR�Q���uQ,6�����H�I��%\t7�/N����>�X�eYa�]j�-�k'�}�^�հ677�R.~���:fJ��`���4�"�v�?����7�>'�Xű~�n�8����⛙��@�؎`{A[P�6��1�aY'l1'eS�oC[D�9pN�e�t �:�E��^뮙�`?��+�&lq3[:�,��Ҍ׀�N�@�;a:��CSY'g��p4�$�7�9��X�C!qՒ�Y�lF�Q�N�Q��M�lOD�����]��0s�`�u\P����gf���^� (v���эfaD�Y�~nVC!vF����at�`0j���u����rA[�r�%�AC���m��؏a
�@�;�`u̲���f�LJ�CG_�Ab4X'Pt]'Ѧ!�1�#�wr^��b�3$Y.F��miQMs �ڈ>��}���W.��5��� �� 3H8,�9�
�'3m���([����T[Й�)�F�{&��Nd���㠮"���	D��L`�R��		��"ӎ�2sT�:c�M�m�x�1��K���~d�����!��D��:	N��q�QAF���0A�����u6�l��*�1ށ�u�(11����dL�E	�mID��M�Nr1ot{A[���`��-F�KR �ht�H��IYa�r1FlO��h���Dj��"%���YD �|S<47��O��2��v�)Pt7#`�W�lI��3�\#�%Y�r1VK�9���P����ѻkp���s�D�{�T�:p>+2��`�i����MSS���Cl+ٗ���܉��.-��\x"\t�L��OO@[�9޶�P��I��¥(�VЅ����	�A*8�\�h|����W��Y	�
o("��6~���$�02Z#�0��⤵m1��kT��t0�FU�u �F����0�Ō+\d�J����kdj���มр(J�L!5f�1��0��$�4��8��0���X����<�9A��b塩�n�O���F��8�0�N�·dt�Ѷ�-g�Kb��MbgC��)��;x�&��	��m1bWK:I�(��Qk'��fؒ���8[FX�$���Ip'
�xO#�[W�?w)|���j�x`�P{��]��a���v��B�r!���O��v�	�<�4X8�BQ���=B�
�K.��Pt1Ö�$����*������(P���E����QAmf}���x� ���h��F�^I��c�2j�z:}�F�K��\�I[��LԱ<;~�ژ�� q���W��t7J�E[���M�,<�	�� yX�hPp5����\���5�ɬ�9:y�$��]I,jT��t�bT�1#SpF2͓m?�r��_���/�`Hp'2ƛ��>��ϗ�����;dְE���#
��S�1ڹq��IP�5G�#5�Űh�hx�}��>�s'�<�'[f�;��K���7)%Yf�RfH�ۤ��,RQ���u�ۓ$��dvKFb{.�E�5�C�EG�b;yo&$�	���Ybd�D�^Hx�f�\̵%)�N%�}�Y�)���n�.���+��f	U���ٶ`�8����o�y8f��Jb��>�/�9F#�1H�#9�7cZ*F��6hƮ�T��xD:vr-�`=\��2D��s�UE���yS��n%���<*�:t��l��]�u� t��C���}ے"�' Oi)����x�h(�����i�.1'���ȒL_��p~�F�'9yڸ�wE�F�0�BI��#�I=F~y<n>�3s����(��^��$4M����r�"�}{s��H���GMYU.{��""�\�iQf?�����g��D=N��z=���n̮c����67������h��G���=�l��UUՀ$�C/45��������l�-(P��V���"H�b|j/#ȥ����GQm�P3Ό���+��ZmKWW���v�vr>��$Y67�"I�p�4PEE	�݊�(����2�V͟P���%�\p^i�YDÁ�`uVIii�%�A�ֱ�c���~,++ϭ\$��($��E����u��90���?o�DA&�$�j�~�Ax|�&h�~����D�����Z�U�h[+4|�?�����"P�89ۻ`�ƾq���P5o>T�_ �f���;x���G^WvEw'�HJ<�w:B�Jԫ(��r�$�#������c����S3A�G�{�Qq"�B�Ν� W���أ²	=
���rX'�0y�DKD��ݻ�I�2jT��[�8A�
뗈(���JfO5X.��o�!�Zc�Բ�u)%"l�%��#�G�b��i)X����f.~ǎ���Fc�l��Vڂ�([P,�ҖX,n�r�uwO����*��0a[��`�e��ɓ���ZfKwwD�-S�Nf�ǲ�Sss�0�شiSz�f����FaN�ɓ'��`XA&n�����ءC��\˥bᴶ������\+�h���'2O,R^�*��T#&]p�	���d����q�=�j���`�b���j�k���J�b18�f�{�5hX�]�b.��бo�x�i�����`̉'B���%����23�iy���Z揭�����u5�Vd�\i��.�Pp]��`6�`��eK�:y�_w����n�0���ň��Nj/V!�\�<@�аS�Hv�z�-��q���Ŋ�NID.:ڭ�Et�7�c�E�cԇ�D��U7�ϸ�a��3Ip'2��k��Y�[q|V��a׋/����������y�w<�T̞�>��t:���VDV;q4xƅ*�����[�e}�{��9�DO��Ωh���-ܝ#����rqV��X1Q_� J��A����^8i\s�-����S݇[i�H�ۜ4N��'��I2a9� 6h܉� �ۍ"�b?/� tU�]�?�{��c7�thܰ�?�g΄�����{w*��x�A�{�L�)"����
� zq��6��S����_�/q;L�����C\�X���hsJ{�]'�0tXlA�Z��Hj�DjѶȲ3l��be�8)���{B咿�u��=���l�Șh��sigC+��u7�U:���m��g�Q^E�&ɭ�4~�1l��C�{t1M7�;?Y	��ӿx9?x�i4v���]@� �������[i0�#ݓ�;qG�r�MdJE���	��c�P	���8i!o�nZ���na���:`�A�>'�b��@lJ	Hp�N�-�S��q'��7�9g� �`[G���»<'��xźS8 �o~�~��ܳ}y���}�WC��_�
j�YN��+:��څ̸r�9_FJEq�Q����+2��� 5��Hj���(sR���u�w{�Sz[b��R��Cͱ���
w��b�-"�/e�-�۪S�i]��2N�|��ߋ��y��#��Ș-�N�n��3뷂հy�c"����uw��{v���������D���+A�8#�OKW����	��s&Tt��MnF���>4MLUM�qK}h���] �������+��Iq�贐&�!�_�p�H�sEp
����V�m4Fc�:fB[S�]�Non��({=���M�Y,��:���G��wX��}��}u���n�	��U��4vGI�ʒ"��Jd�$�XՈK)#9**�))el4�Α���9u�Iy�D	"*c�,ll�D�F������]6�! �v�����i-֙�B�#�J���1xl�&������;�=���a��������o�w�w~�#X���C�����(��Y�V�#�� �9���@QY�W�a�&��hP��^�~�*�tK�bY:��.]'�z0tJ!��u�;����ܽ�h�4��Ael.>����C�H`"��7O�	~��h;��y]�w��l���o7�HK���?��7��'C���9#7��t�(�}*�|���)[8�5��E�S&�(ZmE��3� �X�,ѶX�D��A�҇9�bY�J9޻�~��qZ�-�i����)��w]'�4a,�����KZ�G��XI䈞�*�3��?��f���?��� �b�������� 0n�#�x��%���*h���-ґ���þG��;�.�A����G��I��s���r��B ��r��bm��:��H�$�;�\r�^%ꌱ ��}�H��s�m����j'�;2�m��^�b���Z��$�2]G0(iÌd؟�<��Hڰn|r�=�ۓ$E�E?�	���!߈�5���o�;J��P��u�7)���,���	��}P�{��D���:�j,��}�Ha��!�".�%�}+�Ly[B�b��G�z��#�9�C�=V��O"���-4��@r��F��/ZT�{}&� r ���� ̨���c��>������O����NeE>wG�0�ɞC �C4�$�k���������2���X�����!���Z^:o�Ef�loh=�{TY���%�Y-����`�X=�������mE�(am�h�kK����K)v�9;k�8�+w<�ۜ4N�-��hl3nE� �X$��d�x��s������ӻ{��*P�]ql��_P��IG��)c������q���:pUʣNT��u���:��={`��G����J��SIp�:`JU
�K~z��g[�+G�]l���&�V��"�5E�K���eu{���zE�N�0�6�n���[ם#R;'���2�{+�<��Md�=q�8�	�K�AX	��S� ��ՓB�������3�KR�L#�y� 8��>��>�8򅸦�}�n�l��'��BgWs��s84I��*{���頪b"���88e�k�CSE���շ l1������a��"YXǜ�<�I��bR��*��8ř����0�a�d'壷��[b'[�_�1�R�y�.f#�"K�b�T����$�#�m�l��Iy҉��M���j(�<� TΝ%c��\>�� �[�����ťx$������A�HjkED'Ei���I�����rqʶ{��I��D��9[b'[,��c;�V�>��P�;�c��N~r&�N;��Asc0Cp�%�}!$�2�D��4��Ue,���e�~���՞���H���`�]]��}�BB����?�����y�Z�Ȏ�v:�F&��=s�]�����Hpǎ;�8RmM-
�!�nBpw�#�]��w�Ejт;m�9퉭�E��18刓��vځ��g8��;X���8VC�=��-&�Ut%����w"g��"�T����p�w�G=6A��À����!���F�¾�_�ڥK�p&�~(�	Ձ"(T4��=�qG��Cd��%�R��'���]�1"�f������ G��>_���(@��$���#zp��T�Q��۬��vR��H�:�Bc�$�m��vHf���w"g&WW���:X�+�kOF���y3�j���/� ���G�Q����Ɖ`e�.���P���y��1��r'I2L�4���ϛ��:��:�:��׊�Gh/�Q55P2�=����o$m@+���*[�'���>������J��_ds|����������B$2�_��N�1�),�����KKK{�k��5�tM��])��W�"���Z�]�Ux�^������Nڑ�Mɴx<n(.��I���a��Q��ˊJڹX�Kᯥ����(a��.���c�H�2����-y�-�>m��Ta^�u��z=#�%�\<^k�c��ϖ���
����m�3[T�3�V��\�5}<��}u�dߢ���_�Jʘ=X���|�E[��v�X �1��}��_d����w�����$^��m)*�[Z.�@ ���z�@>�ݦڃ������l��\B�`���������^���/�l�؜���w�B!�&lL��DpH���9�_�������PΝ丆���b�ے��,�%����>y���7�!��abl��ڒk3�U�{o	)`�L9���������R����u���;M�=�h��|c]���UPwʩ`gIr��P�y��-�?�nKv �Q�v�1�GC�M�D�}yCsD��?�U4��";o��k�wvAK[�&(�%�-�z�Śr	�0��3�tvvBkk+�My0 ��p��롐X��ј�絏������ֱ��fV�̵��ƌ���ŝ�Q�-�v莘�^�-�bm��pK{tvu���-cGUä:q���h�f�t�xS׈@[ƌ���u�����KGWW���yh*.��T�ı��D4g}h��)LPL�cmu�8��4�\�:6&�v:eB��k�8���jz�1t9g�P�?aK��um�7k�P[:�8�c����q3[�g�5�Y������L��:�m�BKkx�@'�@���`���®�%�eD�ZSR��$��I����狠�����߾|�p��i�s�a��
0��)�6�fX0�}��נ����ؓN��[�\.�p�"9�j��M+��\�ݔ�߰isl$���)�#8�,ASktu�'���\�MI��/F[�w��x�S #�+�ˠ�����ybUQQq]<�ML�VZ�l�DB�˃����\fQ,�(R1��U��Cc3�c��:A܂w��\
�ǂ����Yp[�bmQ*�u}���Z�s���dٛ.E�����]���fQ��I#l�v��z�x��V|KM�A�`s��#
y�ll�oj6M���V�.�ZhKMejl1Ux�6���Hp|�r9��l�񴲬Txt=�RS����ڂsѶ��%�9�M�<��pn�uL�-|� ��[Q�;f9�q=Pn�-^�Uy�Z�,G���1�u����R���0Z����%�)����ph*:��	�If�V�t�U��̲`��/��C�FJ��иaTΛv�#�TP#$�&�����|�1Ph`tkWvb�r,��CB��������DU��,0��~���o�-m��X�ș�A����IpttfU�-��7h�-�����r.�].(�K��m��<Q�̈��7:�� �X��6���l�]-~�q۱����nn���*2�,w�;����Q��g���#��p[�����c����GiglK�%.J��d�p��(碻Ѯ�L�L�s��DͰ�|Fق�mAǢˠCF�h:�>���	؜ӨT6�w�-�o�����Q�p���fF0I9�E1�\�k'�ot��Ta`� e�^�q'W���J�e�"�	"[�l���#$�0���uM����
D�=��dk��%I$�����\�r�B���I$�h���Y��.+1Ȣ��d��-N�αY�=o���r9c4(������(��F�`��Q`H���`P����Hw�:,7��a=��ڳ��l/e:A�`�..���c��r�()T7��rbDX���]���������:*��(t�T�~��@[P���˿�#��2�c�d����/���0�|.Tc�;����--6��$l	A}K+?��(pזi��r1nYbc���s���똱���A�JjIQ�hG��Ω$���Ƶ�E�Pi�x[X����D���q�g¹(��N�炒	��P�;����=*�|����J�����1ϭi��C���}��ԯ[��Np�3�K�)�{Էw�=on�o�0
���~
���t)��E|![0(&�c��`�}���7����f΅�S1zW4|+4+٤Ԃ�@�GU��m��s������F�t�:��R�&7�8ec���$��>d�-!�c���Ŋ&���,x���,�#��� ڂ�̈�,ܙ���9�y�0$Uֱ�PȴrI8�1���s +s��Y
">�Ǵ�����<�h��c������M-��b䮭t��� jD�,�!d���lL�����ؙ!T���,0h�FD���L[�X��g9Q.E&��<$6#ǎ	íK��D�޶=���V�����/H�<Ҷ����k��C�Š���0���`G<
E���-/��=�~kOp7��������j�+㺆9TE�;>�=k��hW��@mn�F��$X�P-�H#s� ����Ao���WQQ��3���8�oo'"&�%dzÅ�|"���
����"��$�]���J��N9�����������nK��������n/(~�m�cAL�6|�law�Q��{��ߵ�
��������]�l5c7]*8%�]�9�ѹSn�-r�y�Q��`ښ
S
Oc��S�%"���3Ԍ�A�$�#@[�
ո�(3�\)�Xkjz&��bv� �]�݂˥<d�.�T�W����w ��+��N�l�;�Rl���ͮ֭�?���XpW(�=G�:��Ͻ�:�p:�}�=��<2QJ�3�1�N���Ol$��: ���?Y��k:?�S�D�"K�89�v,����Q6���ك[}1�zDЄ'�n���?�����s�ʆ��e�-�KL��2ء��+��ae�v�!&h\a��x���{O�色��Q���PQ�F�>�u��
ݿ�$������~���Q����gڥ���Ol��E=y�_jK�3�;�p<����6v���i�bs����a{��Q�(��g�J��f��>@���H[D�e(�s�����z��}��3Nkܩ����o�$v��u%��0��2q��gJ{���M-bw?D9��灒����>��Z��2"����˱����C�A��)�2H��=�s�ّjK��1��&�@�Z@2���/����`�Ĳ9cH��@�w:���B�M�8�#*�\N/�[k��m�����ظ6\�7Ep�(�;AX
��]-�������d/�h�hCb%)ٯ�tS�����pтip��Q�T>�����#����d4���2�3��6�/}�e4�I��O�5�	~r�`&��?\��]�ђCJ6,���_�Bc$��:���Uv ���!+�@��#)|;.SE8+�Mk{'������-��bU]ôa���_6�L,+�+��X����>l����V�<�s���`��IVق~fbK6�@��T��%۹��c������Э�����lɴ�XU6����X���NGtیm���2蓇b�9�PL�U�Sw��I1/qZ�n��@"���y� ����)��p�r�/�+������Dw,_��Y��p���x�΀��D��@|M>���9����z��r��ƝT.���?�m����LJFC;�A�'��|�Aw��5���L�9j_f�QN�|g�D�D��e�28��'O�����
o|�b�1MR0��,	����~�͖��[��6�ZƖ�f�����.[N���_�Mr۽���y?y � "$���A���c�g�q�p'
�1}���p݉G�/�{~��~��t�X��ajUY�k[5Ê�=͝��oH�O�Ȁ�@Nx�.��8�����6����pͲ�~��:��;�|���Pu#� �@�.�bn[n&� �M1^p�"܉�����ӎ�����~<w�d��I;oju����p�=O	�	$s�nΐ��F ���!�#.Eɯ=ry�����	��yS �yr�6f��B���<y�'� ��H���CSU��j�C]	� ��Du��:V�Hp'
���p�){O܏���?}q�؞dŬ	�h�hxg�~ѷ�g�0�f��I��<W918�6�e�Ip�s������v�> _yj�6��gA��T���R� � �B���e�WEx$� ��.�wP�@)e��ٓ�	���	�������3�;����9ue���ӌ���]�C`b����(�d(�m�tFȲD����_�����W���gO�|��5�_~Y�9��&�� � ÉxIp'� ���!th*QH�]��ŧ��nPd	�l����O���b�t������sP�$˝����u����X{;ؑ�w�ژ���W������p�I!���~�]���������gG���e�S���.�Q��QUK$]g�׊$M3!y �Hd�$)��>�3��i��˒�zX�j�ʪZ
6ۇ$ɝ:޿��J���g��X{q��b�C�	�Td��-"�qP\]ɗ�x�i^�ڊ�ݾ܏��A������ZZ�x�@j�?W4�x��wE8ǋp�H4�4Yf�d7.��=�����D��N$��t�\.v�.P����~J�Ȁ���O2�������>1`�ras���<䞟�#�+V&�(��,�����-��+���<��w,'f���>K��q��["���C�x$�~��C��\_�`��՛�v��a6�������ǵS�ޙx�
�"�X��Ñ�"܉¤��������a�Ժ�~ϛ����o/<���1!c�7��bYUU �5b��7�"�gv�@0�O��&l�o�__�����+�Z��^�U[vr�nieGQh��ob�����{�&�:�� �q�M:�]Q��&G.5�J�(責+�eQ���n��&�^P\Ŭ3/c`�@.�(�y��;Aךe]C<ީG#Q)ՠ�]�;�\P%��6�T=.��.K�������&�9_[s�u]�� ^�M���:�N�d˃Ƈ�������1ţxb�8Q��.M��ĺQϑp���QY�x�rit�ף�]If+E.ao	�w��\6+A�}@+�ԍW�Y���c�������:�Z�$I�cJ_���s]XN���RO�I�{��%�^b���I�!��"�n�\n?k?Iq{v�yRH93Eof�ڢkZX��:!�q[�a:�3Z=�W��$lq�G3�5.�/)���Ud����+��=K��t<j�BYV�(�C���ڊ���"p�J$I��_�q���8*��̎f��ì�v��%.G�l�a�M$�V%��{6wd����-"��e�H�pt�-�$E�%^�Ou`�������&�p�8��߹h��?�w|��U�M�GI<�"�p��<�8���H:k\�ˍ�Y�U�%t�}�	�K��������d}*�F��B����uHά�{�
yd~�4L�d;h���^��3v���ј2+Q �;C�QJ�pX���tEq��'�Q$��l�+�=b���"6]L���63[��G��[T"����?���zH3�w���I"�v_��B���;+�b��1�2�r���2��Ⱥ�
�ݷGu�R���(\��O|X;��g����[�rA[JV��˹�zR?�3+��H�����^g�,{D�'�sl{*+?I�z�S���{��sA�~!�~{�O��\�Y�y�xO�|t��:��X���=/iq�&T9!���y��}�p1Q�E�D}J���������'5�}kv��=�Вƕ�|�,K�
��T��wH�����H��_���c}][	v���M[͝�u+�ޒ�-3O�l�m��)Z�G6�i]�>=+Z-{�l�J���P%��z���
��Sc��1@��h�ҷ'T��<cϞ�V�z�7�M�3��~�}ztSH�j��QͭiAI�GR�z�'� �\��1�����Rj����J-[�5��]��H�q/["��u}��xq]��T�+�g�.8��*mrѴX�l�6D�0Ķ���}Ek�I�"�^���F�Z`9��t����]���}�Vf�5҈�+���G6�`�3��݂�m����
4K�ЊQ�Ey��#�*�c�����8��#Z�Y��5h��A9�EE��0[Bܖ..��JR��p�J�-n?�E7A{t�r� /�ܜ_�+�q�I�l|8�C�\mJ�4�O)�w@P���s .)e���J<X�g5_G�Skc����0����m�­�{��?��s��:"��K�B���g[D�p'
�ww��_]Z��rH�Gڻ��y���@&U�ezi�6&��u�Q�v���pQ��Ƨ���;�^:n>�(�A���Mm�ӧ߂G�m�x����.y�+����Dr�b�}z��M,U6mUp�'`�б��$G5���d�F"��D$w�<t	���L�y�RV4�_�.�3�=/��]��}��x�O�Ep��^S0����&}��)�����2D$���1�=Qy"{�D0v���J��枠|�T�>>cm���n��in��%�wD��O�1ܙ��Z\�c�%Ee�'�{ʺde[� �p ���r@	��
�6�l���f���PU�7Tt��MMO�/Z��
llQ�����ʈ��cm�(0:%/t��E??�FX�	^{����]�L0���ĈN�y�"�K��]7t�\���K�J���R��"V�\(,�Z�?��a7�C�y*��
�=��*�S�T�{M�z�磇�-��-l�EZ4a�؂w�Y��F"��5&���=�p;z~W%s�K��`���k�0[$<��LD����z�jOw�Gt���Gˎ���km��&W�?��*R#�c�ڡ'�l9%�^�?��=.ɽ":
�	q�q�n��a���2�Y+��H��j��!��,K���\����#�9�2��!]˓܉�ye�nh���"TWaʈ��{��c@�l;��/����6C�K���v"�cQ<^{:%$�w�s �\�><��f���G�����}���g��o^|�Gދ<��6�&�cڨ%����W�l!X�	�Y��)"��[�*l�4)�I<3F��L�N#AɫJ��ݺ�l8��3(ʠH��0
F[%?�;QpATvA�?(���E}��q���X�C��I��T(�K%�k]܉����O��=mр�|��yl�������'���c?�,K��C�$J82\E6�t�!� t7���㕵�����e�̂��؅:�q����m�����mA��� AA�?��Nd�m/���gM��c�{_�o{��>N�=�e<JB�~ՠ]�b��T���٬�A���	���5[U��S�����gϾg1	Ν;N�9A�᪸���G�����`{c+�H�  � � �BA�4�y	�F�fӋ�iw='N3kʡ���ڰ����D�*���+�cg����}�@�$[)���+/���z ⯪;��F{[���G�Cf֨
XPW��anm�����y����`ws�?6쫇���w�n{e�""34 �p'� � �BA��D�y�_ظ�?�}�m�#�m�{�_YE��UW�a�:�;t��}͇{����{]�$�
AU����[Lk��zkW�;�� �yˁ � � �B!�nHp'�;�BM��O�H`��#���C������ � �$;�AAA�.�}@$	�D�����J˦N���^b �	������:A}�Nt����QAAD!���N�5�S�{�0����1&W�P�1�-4m:qC`��#��N�� �8c<�m�&����`z��������aNm%\���=_�CsW7��}7l:� ;�[��R �����JX2~ԅJ�|�$��NA� 0�d{$]y>�EYѩ1"�>�2}<<���g&Ua���?�|�i�P��܉����3�kK������a_|����u��
�^~:�a��
��Ν7�|��O�7�7�^�}�6T܋G�O  �p�>�g�
�~�h�:z� ����D�j���'agc+�Ձ"8yz��1�M�� �&����|�R���- ���p.����YC�nj'�ʶ���W߂�����,�.8e���)��҉�r�<	���UÁ�N���>��ƄJ����l��;���5��\�(�3:�ǎ{=p�����o���v ;1kt,�Xs�T�C��1@w�ԇ;� {|���o}��ϩ#q�ױrVo&U������v��M������s&C�����~H�k4k�G�r��5X�ytD�y����c���[a3�� �OU]�`[=j�(���+ۺ#���I�-a󞫖΃G�l�=͇_w�H�>/�!�Z�!��9��W_��_��ęO6ĥ�p�:xc��A�ǥ�헟�U�?����i�q,�n<�������.��5{2|�ԣ�Y6g�[ZӱlM�l�X8��f�*�����z16om��!6��x��^ۺ��y�С�D^��:6�c�6b| o���Y��?���'������D{Re�M�y����\�Sp�PǅGQZ�4*����u��#�0�"��D�W�/����z�.���0�G�/�1�]1�=�ق�޷�=Cc��J��g�����ކ;^x�����b��y'������|�lgP ���'��u�d���l�����9�^v#ݤK�����<�?x�u��O�-��#/�7n:�h.�"-lqr�C/�S���_^
'N��Ж�fX��-�,�6��|�l9Ԝ��{m�~vች����ǶܧՔ�]������C��9k�$�Ŀz��}vcrM\�p&�0mL�.�=؆�l��X_����݆;��am�'-�����ᣯ@G�}�Hq�����z��F�~��'^��3(tn8�(�ފE\�yp�&x�����a'K:����;.f���??�����O��/>�ב���[_Zw���-"��Y������ˎ�+��;��m��WW?;9~T�k��xq�s����OM���k���}��˯_x�V�+J��/�G���w?�?|�%8���O���MK'���՟�۟}��̱���糹���J��`Ֆ�����ö��N:�8l�o�|�9��wp屳�Xm�~~���X�"�qB�RiŬ	�gw\��z�C��3o�?�D��~�	�L�)e��!1�DOF�#(����$�θ�+���A �;{Q����|�^���$6Tuؕ����N%=�;2gl5�U	�4��Pd	�f���N���N�Q��þ�Ͽgy�h���.6c�����������������HlO���~�?���S�`��}_9�G."w}������aOK�L����u�"J !�����_��'�o;��/�[
�3�_����5����"n:��#)��y�#?��A���o]̣˲�[/:	���ӧ��pղ�p��E�}V�i�*�泏��-�?j5��}D��/:�WlGN�5���������p��)�g.�Y*���?�n��YX�q'2%1U�`*|��}_���~s��� �_>v6\��M��gܗM��?~�A,l�?auf7=�
���S&�����q��ˀ9�rV����3��!��Ue���O�Y���K�98��tጌ�{+�)U}�~7�vwr~���"�݊�]v:ۑc&��G��<����lN��W��E�T�N��k�?����8e�8��/��wp&��������ހg?�>�op^����{�38>/�:�9�;8���7/�9�UY���ջkO<�;��p��A�)s����^�d��4��+/=�d������'V����Ta��qMs��S?Э��-R�Y�1}�7�Hk��i0���s�S*(���Ip'
L�ʒ�cm#���iupp��	PV�L�t��G�YMzP���n[�������ߪ�/�Qt�p�t8nBd�bϛAA3=b�o~��<e�q��>g�?I��LSg7X�.]�S���B<B\�`|��������:�x����v����<k�=��O:
^ټ{Ш[�Y2e,��i��өí_8�x���յ`5c�K�ۧ/��x�n��?] [5��1�C�=������rD��H-�-E0���.�r�>����`3O3dg��ط����<恶��h�/�]:d�h���>�խ������zJ
���`	�4c<<���B���/_1@lO�['�v�g>�� |֒���s��o��p����ڔ9�,?�9�ll��%�3&��Y;X��}�q|��묝ע�{ߕgZ������z6ܿf#���U��-a��d�:�qn���DK��<@�k[��Q��ccs�b{*�͜ _?n.��u{8u��=�J�����s��h��?ض��2�?�*)��6�f�Ԧx3��I6=�#��,;>{�	  �N�Gt�PD5J)C���bUE����y��6�=m�8(Isd��g޲E�n�7�p�T$��Y�:cI�ƍ���̄#j���ok^ܲ��ɀ��o��.���h��3&�o(�'��o��.9r����LlO��Q�?vb-��ث�eҞ��Z���F�c�d*�TPdx{��3��}�n�ue�0kLSv�b=���m!�_���M0�#�x���8�O�w���O��7-��'^���^|=]l�42;Z`��J�#��ק͞_g�S�
dy���F�Uw
�<k	O��_o�t��H�i���d*�œj{S�%������~����,����)c��;��[>w
:S���y�m����������sfi�k�/�O���ϭ����{��'�{0N�3�������X.�����u� _8j&�c��M�=	�{*(���~Ĥ~��e㶕�;���d�H���<�&���9����������ݥ�w)���z��%�R����R�����#���+��$dBy�ʀ��9����3��n[�b�g��g�-����(|�Pu�`g�q�ڙA�Lz���c����/.瑄������Eo[W7LU9@<yc�>x�{n�O�%)�B�_���0"��K΁sfM��+΅��X���QX�g_�뫶��g��J��SǤ~�z�C���?[���?�߼�����:�������`N�2�0��EG���r�����]��O�3	~~��Y��g�ft��ъ�: ���4|V�<��`ځs�O�_]��W[>s<�Z,<ج�����	ѱxza5|�m'w)Μ4.8i	�8�l�%~�ܓ���ӎ�7�>V�畜2k"�k��{�AsS3x�^�:u2�I啍;��ǝ�<m��g&�9x�j�
�n;1�(�n~l����a�F��[�����Y���ys�ҽ����_�ѻF��/�ɣz�V��0�6g�^��,��9�0-��R_cc�6vϩ�;�����۴ߺ�jgFyg���6�ϐ8����GG}��]0#EIs����\�Ǿ�-+�j�j�&ZwM,"
?L���5�E���mi��N�7<�sGN�ߢs<�Z�S�?yLoj@d����C/�G��ީ��޿�x6|g�Q����yc��*%X�a���K�t�Rx������@��[lPpǃ%RN�Y�ɒ}�=�A��8���*(dƟ~���݈���]�0�ⴈ�6��X���ހC=ۃg���ˎ�s�?���x��2���l�cfÁ���`z��`��QC�BY��ꋰ�w����ġ_������Y�*�g��mu�+���*7�2��"���j��k����	��Ϋ���m�x��w]�s�c>��R��&��篽�G��G�� �N)��΃9�_�G��S����w������P�T]����vN�0eZ�X�i:�bJM����{�G[w��8�G�]�4�R��/��G�ON9Xu��jfKlo�F��ZS�+|577��W_��77{}��	��wD��c֎�养��ȋ�ܷ/�����hP�M��Ir��}͗�O�A����3��������s������oW��9)�/Mq���{{�vdӁ&.�?���{_þ�J�ݝ���>*��P(�ޙ�(���êM;M�w4'��;��u���o�?����iu���7^�t���/q粕�������������<�L:x���}��|���b�e��0oL���yܡ�iUN�>�;�S�!���o^���q6��?s��](F���c�\��VFMO���'V+�#��y/��'�>�wGɄ�R��wbD̬�]r1<����+/��o�@�A��b�5[+�Ͽ ���F�F�{��`ܩ��E�EIZJ�pľ}��)�8�����жv׃m��O)�>hI6��΂�Ȫ�;�؞M��'�%���l���kC](K�Jឺ@�:���	?{�->o� m��"KRl��I]8��+���,(T`^��7��<�����L�?\���~(�09��w����-0��z'�RJ�}������'���a5���6wڎ�-��xρ4}�}|��ז���x��Z������--J4���`osZ���������Mm�<B�Jp�:WO�F��m/���x_��=�~����~c�_�<���AR�a�w�z��I^ݲ{��v5�W>����߉$���-+�)�~v��;�l��_|�?�d�7!M�3��}��������9�� ܁���x@/������E�����y �x����/���6�����i�<��~����}�zRlG�J�;Cdɺq�4�~��gնD���0%�䅽�q���5������Y\���g�wD��V�=i6���ѱa_���Z����%�g� ��Ș����#�t�ֲ|����;V���v�WW��3΄���}�y��v2�	qM/�U��`�ѕ0F��~�s�;�`	�}<�R�"D�����;1PPOO)yCw<�o����ç`I��S���������5{�] }oM��	�|���, G�D�aʕ�);&�Y}K�f�Z �g������̝|��/�_���l���ň��<� �[;Ep�z����4���͙��_�_�:�u}�csƄ:�{�����}y��l�|�������o0�B!���olKy�L�YV޿�M�*�Z��k��6:T�z�t���d+�~&��IP|��������p����|��c��bj���(�Z�dǨt�jO����m{���x��#i��������	WZNf��?�8}��ｅ͕�}>����cL��mt�,��~�锣�_N>������惉s�{hͮ0*�_(�]ivۑ�ÑD?�j������)N�_=�z�؎T��P��:R�Od��*.\'A;1�ރk7��/X�w�!(���oGQ��Ow�GL��ZV����?S�|��L����?�fϳ6�	d�s���G�i����n{�E�}�_�H��g�,ࣸ�6��n6�F��$X�ݥ-P(������ʽ��:mo�)JE��[p����7�Iv���Mv6�Svd73;�3�<�}��r)���%$��������2��U���f�Y>�R��
��3 ׳�����<-�P��Gw�c+v�N��S���qt��a�ՙ�c���6���*�Z05Z]�%�pOOu��\p��V&�D&3[[�l����^�wV��8��Mرh6���f�Y�3LK,���e	Ƨ� %%���N$f`�����=�11R��)�}��DܫV�+������Z�:�¼Tk����=��Њ�pB*�wG{���,��?b.`��D��q�½lPxEcLd�@F�\�,�F\��c"���`L�^p�����q���Ȱ��[���i�� ��$Ꮎ]T�<-'��  ��P$���;�N����R�����A3����o���R2���O�&Lγ���H���Rp׶e!�~�뱋Xs#�k��a��h�=�\+�}48���Q�� w,���A�!���8�lg������9�hY+m����UgY�p?�t>Nc=7�l��ٖ��(���ێb�٫�|�h��g���7Rm�'������w���5`Y�&\�����/,��MJ�>�d��VlA?�3��\�vO=E�	�7�؊�,{䓻F�)#������#����	τ��j��V��ya#��V��������7�j���5�oks#]c��!�Y�ͩ�,�I��0!���1�s{,�;�k�K��ﾭ���E�����Ÿ[���6���\�N�	n�RD=��%�Dq8-��v{��S��bJ�0���$�{:;�}��N���waڷ둘WK��N��>.�0��йr�ן	doc٦ZEu�uA����lCDg�L�E磠�t��ƌw/$����Y�1S+:����ހO܉��X�A��׹T��Q1�7�f��Dq#Y������Մm�����#q�µQ��b�r����F�C��o�9�����sqx���ﶡ�3�[8����bTT�r�=��V�=��4��X�7���{�]3t_ҫ��q4��rf�뚂���2[�Jʰ��uL�/�����&C�Ĳ'��S�Nqn�Y��I�/RE��O3|�.E��D�$dS1Ry�8\+#�%G/`��O#;�����^g;�3�����M�t)7-��Y#���u�dS=��&,�ڼ��-y�O�j5��ܨ�x{�fsG��Y��)���f��,�6�������;�r�,|�K3C�E��IX2��F�;V�6��fcPV	�+���/���&�H����u����d�M΄4��U��V��W�n����v���.MY�4ҫ~ �
Ծ4�!j�7���:���
���sn.�s��Jfk�4��)��1��PQ��i��h���={p;>c&\;��Z�5���T� ��:��8�&jO��Ԩ0��Ԥ�"Y����tL�f=Ro�� �Y6��\Mp'�$߀h����}
+L�f�5�*�wo�Hd�I������V�Xy�k�n$�X�1�t�I�<a �/i�u�_X�q��xw�0U�Z�:�����S��k���A����;�C�lR�X�(�Ż��	���¨MA�����^��&u���Z��>��|�+���q)v�>Gn>��!�:��-�S����\p'v��$��&>���G�ocv��|�kD�N����lƒ�'�������}�46F�HL_s��r�̨�1��=����'.cߵx:ٳ�3ch�]�g���~>��&cH��N~�fۉl���v-ҵl\�4����<6�iI��tC����j���۲�|CЀ��`�c3T�d�"�"joP=����TYr4iRG���J8�2E-j$R�A�|�-*��>�jXz��xKx��~t�N�(��V�P���}��(��QH�B�k.�s��*��J_�Z���;�{?�/]FI���Gs��5w��c=x6!��6��[�e6�6��3{��TPW��d���1���z(���V���k-EQ��R�-����-G�5�Y�_X�7X���f�YX�C"�>�s�����5���2K���q,
��Z~�_�2>*̧׸�1���v!3��@k���ps��z6�D�e�����,ۂo�j0�x�A�: e��x,>�;��yz/�����"q�߶��������XǄ�y�D���&<W�����)Do��?c.���ۙSIu�)T849�4�������W�Ok�İ$T�c����ͳ������@�T�[�G���%8����-e����S}Qo�&p�Ϡ���=Q���������� ��+����'.�'�'����<w���[�!]�h��)���D�Wk@Y}O������=}�|F��������g����gi~8tV���d����2�3$�� =������1Q�=W�D���s5
ϵo��Ҝ{�'��R0-�8���pn��*d-���#���QU"�(s`��1KkB���9�����5�g]�W:�:���5��(�fHX &F�bB��LdWghx ���e1�a)(��ZQ�[��M��ܛ�n�G<�>�~��:��r >_�=��?�AC�A"��%���黚�pWg��k�t��SD�N�~,�i��o"��7����Tt��bޥi��8#�вz�?:�'+f�T�A���m;�m�}NL�N���/W��	1�k��Ϝ��i��a�I�t]�}o�����ܒ
���3n������=S�'g�P�v�ӿmA��f���]����������G��v��f��<pB�Z$��W%t?����G/`R�06��-���*k(�]����c7����x��-�ޙ�̺"�98(��/v�E=c��+N�����R��~��}B�j�W�{�+�vbh��l�u�8�ug�pQطE�� �ݸ�%�C2��LtO-��A�)�a�٥���]'�ӽ�MY�J�~t*i^�8�e}�!�g�?
����9(��n��w�U#�$$
+�S8��s�����Em�8:�����}^xv��6��Ҷu28��B��c�h���)�}5�M/�"�=1�kFwF�P?&l=<(ʢ�;	T�|�mJo�ݣ�AGo���$d�p*��Bw$0��V�MLP�؄/W�x�6���i���*��X����ט����I��pNE�R�N��;ݝ�����h���������\�=!V��
���ۘ缿����0��Ƭ�
��$&�Gygl��ˍ�|���8��e�ޫI�r1m�����e6�.����F(Sm�����BT�7��X��tcdo'��M���Il\���3�2�=�58Ux��ի��wϲZ0����5����.�����<�r'��v�(�@7g��ۢ���~P�7��8y�_�ʇ�DH$
����wN�����~���Y��bJ6�d���z9;`l�06һN��ܭ �X���g׮���c����PԊ#R�V��ڢ�?��KH���'��X)��yl�l�i&l�Ǩ���^�O�F_�9�N��}Z����=+M���戵q�7�$&�k�^�/�"�AS!���,�D�rZ�������i�p,	X�๱�8��2�9pb�2[���4�Y��%��[�oB9��\p����}�HL���.G�i���ߧ��JF��Dv���p�n��
�<��F��S��:;gÆAjc�s_i��������<#��Zq����C����Il�mG�p8kg�ն�|��P1Y�p8�@~���=���|jΧY߾����1�'�+��.��?(�M��E�ssf"���Y�i���ZXmo�o� �w�믠���<u�NN�Fƽ��R�L�Yn�w��C�e��ɶ�*����ʤ�8��6z��c�
��Ԩ0���(8��������]�a�P�fj;]o��;�erwaY�$���Q��0w��O��0�[|1gf��Kk����`�v���4�g����"XWmN����N�)*ĕ��N~����p
0�3^���R�c�Pu�/��i��t�	�޳��;p ����e����na�5}��!X�8*&=%t��:u��]��5p����J��1�4�;v���]R�����W��g�N��v�jn>ʅ�/�S`3��\c^.���V���\��X?\�l���*T�N&��I�*D\�pz�p|;o<{��U�}���(tŃS���]Xef�ֆjFl_4�3�����J��N����Оg�FR^!��� +|ɱ<4@���ss�=?o����#>�k+.�d�].z��;�v�
%{i
��e(*�@�w�E2?�~W3r[d�m��E���~�/F����lׯ?��Jm�8ډ�g��4��T��L��.!�,2�#Q&4�^�8�	'3�]�l�Ч};���4fMf*v4�k(�^�T�'�mé$qxy��������8t5Yc���������\\�~n��B�����ƣ��"&>�%��HX�"V�M�XP�����t�89�,�K,s��eR�{���:0;/��cK��Z���|�:��±P��G�a�P��K�=�
�R��ߎ]d�Ь�o�apq�������u�����v�ߓaӅ��Q��6��i����捇��-~:|��ɤLVX���'�xx:ϭ���ki�d�go{OW,�o2��ˏ_�rP����f�sB��`
�
���ker�0�sub��Upop��c4](U��R��?Vnǥ�|}�dD���}�Bh�-�S
o���/���7��&��Z��6"�آ⨝���Ж�r�����΃����N���Q_d�{��б�9?m��,tW?q�I�Cj ��.���F�A��HL��<4�7�1y{���9�H�S����5��y;0"��-��L{OX�]±�y�0�=��?��lYƅ	��q�������#�sB�5_G6���Ú����8��q�	�@�������ݬ3O7Ϗ�Ƣ?w�ñvh��ZV:��ćw�`6}�O_�5B�Ս�������Fb���Ξ�]�|�:�֓=�ޟ9�͋)��v��6�zd:��+��?���߬���X#���l��k)�7�1o�H÷�>��I���[��a��9��i���=u�o>Ԣ5�
Xw�W�\�Ns��7:��ũ����C������mO{9�r�j�?7�o�ޛ^/�㺆b@�?�Y8����Y���AQ��̟���GJ~,��c�ٮA������Ι�T������8_YY	��
�T��H����Q8���%�co�s��ۿG0�}
����x�,��[٩?�$R��͆�\ԑJ��X��y0	ؒ���;Y��̞���}(���p8����iL|�{��G��ߵ�����1����Ij��Kǲ�>}�	�-�tno�;���V>4��$ц�I����_V���
�V�&#�e��h��U�=t�4<�r�+��FA��'.�����j�����Gt���>@��]�_�����ɻ����{��mw;��W�8�[$���nΪy�@J3VgJT������R%�ո�S�J�:"B�⌠���F�-G &�#�;�y�پ�VEf�)z�kWUe]y	�r��$8�r��8��\OF��"��Ҫ*쿑���B���R&G��LE"q[��b��.	�J��Xܵ2G$�>/�j��\K�'f`��k��o&E�y�Tr&8k���4,� �0�Һ��F�X(j_8ן�~r
����u��{+C�:K�a���subV3$�g�*Y��m$n)c9���1�z���V!t�l0Pw�	��b���۽�0&��r�~!��m��ۊZ�u�� ���~�x��m[��c;*��[u���>����##���N�����)κ;��X����YƲD�i=u-GN���{�a��T��@7G<3$ue��J&t�`q�]�R�A`��**.�j6ł|�5櫫�wy�e�:w��d�64 ���#H/.�>H��h�p<ѯG����5f��n��gh��2�L~+݃Ll��P�--�w��b�J�EtmH���O���롱N͔��cHǠf��ө!��
�vv��1X5���wN� �]�9MEG�S4v�(��jO��,-{^L�5�����L`��(��Ve�ѳ���N�z�U�����5�]!���P�p��c4v�7�A��Mg}ay�*v|T��#�pc*&�A-=t��%ÜH�6����#l�Lt�:��c��s'�\���<ީ����=��p�`#���ɤ5��+����r2��1E<��]i)zj	�_��n>�z�I-(ſ6���t��wl�-�(�:�%����til]�5o12-K���5�k�{=m!�/�*��'���v���� 2��G��8c鬉1@b��Qͳ`RG�n�v^Xd�c���n/t���B{/W<m��b!�CÃT�8��Ĝ>�5�%�������aWU��z��Mpg��̒6�&6>�c$�BS�WZ�]�1�����B��(�)8����a��k��:M�dgc��KQ�t���ok���i�؂���NIi��������z7uTnv�&y�T���˪����k۸஄"��bSEArΜF��Sȋ�EUɭ�89���3��EG��K�6D�l�v���í|�p͗�e���jӽ8I��U��ߋ5��)��,��$WK��a�E�]L��b�ԝ(���=����^l�DWg�e�nF�:��.�Q�nZ���jN�)Fv��3k��	qp&=�6���D�"��/�/�7{�a���9���c�e��KK���,$�"����D��<�����#urK,��pn�nW����F�lO�*S��^����E�֘�}^r�yi-^��R��Wb��1�cC��L*œ+��Z1��R�?,�o�/٨7�5�L�NE��;�+���'3�u�u�
��Rb����ā/g��y1-w	�E5����9F�p�)h[��3A���>��㓽a��,*:��;77��&�,'E7Q�����BT�R��J����EUi	�\�������>�p���s@ \��a�µab�=#�m�@��\*����Vxl�C?�U5�����Ns.5�5�(e���u���3��@F�Ƈi�d�ϲ4ʴg0xa�q��<�:r/�ꡊr�quU�� W��j��.��C�u
rJ%R&�UJ,?�WV��<��O����p&���=�h�Ӳai.
��l��$4�Aؽ�i��[��M���^��9R̵L���Ԉ��K��{4Dҽ�bz8kgX��%ԁ�XkP8E��H�Nlz.8���-������Kk0/�+^�0P5Os����w[����n��M�����P�7c8^\�����e�]��Sg�G_I|s�a�m�}B�TO�h��>l�A	Ygݻds���.���HL���E�}���h	�
˫��ۇM����4��*�K%��>�p���TdIY܋��q�ݧK�<z=7�
�vd].4����'�������$�^�F��x:-7�*`,B�tj.�����6�Z�%���h�ɱ�xu�n�su�X��V7�Y#�b�̱��E�U@��r�DQ3?���WwBN�n+E�SD���z�����iF���N)���C�vj��R�{|v>�PZ������Rr��Wַ�2ˆsq:�{VQ)J+΍����7������Yu�.75��²
U�:�ʤM�i��S�I�S�C8���cS��X#]�4k��|�
E�ɦ����,p,K{O�vj�﹚N�2�S0>�=Z��l��܀k�:
��2y}��C��i+���{tH$�ዽ�`	(�l�c��Y��+���,�h��K��
��Q2�h��Q�xc�`�|��"���z��^����J�;��;�hV9���Y�*u�_m+���J(��yYe5�Kʅx)=�h��CMm�m/�s�CEe������X��9���]a__&�pbd6$*R������o�t�97aI�S���� ��{P)tB�J+�+L���`yuJ�gL�p\eUu�՟Kr�e�Z�Ϟާ.�d�W�h3;�J.�3�C�����$)Jm�Qlc��qS���c~Y������rwTg�5f��\�kL��J*�^YS[Yݵr�F:��zM����m��U͋@�fHIy������3K0��nO��Q����	�VlTQ��3XgeǑ:|�?Z�<U��q+�������le��E�F��ޚ4X��W�?k��l�h�G�z$ �TV�c-{4�[�`3�:[+$쪳�\�Ŭ08�_c��+I�:�aB[���&�����R��o[Z�����<�w�f|5w,f���}$��rfv�'K@V|w~��������������W_/��8%ꭣ�B������?jk����H/д)�q��8�"^�@ě��R�P��GTSS�R�Y����uY������n=���ѻ�x�HDm(��?����V?6��zC����h�+3������1�w���C��n���PXQ�Wl'(3b��+lj;[v~:i�	KABCj~�J�6V�U��$�"v�e�5K�R��g�G��o��9����HM�����xdH6��p?kJl'�ӥ	�Iڂ{�{��7������H�
����tm��-�~*9�y�[+����݁��X��������̲��������vK�^h�*�V�Q�ƣ˷1�)�I��q���ߟB[�2�dC4��X��L� �/�M��/V!.��F���>���)PA�H�	�ل����g�u��α~$
�Td�X5U����p�Jk���Q�H�Z��.�5ձ���I"���0$��nP�[���C\��7©9�t�ғ���"��B��3����>�>���}"q��]'���ql^"�c�P/�S��:��PP�9"�Cav?�P�QSP�¢�w�W�#L�L���M�I����5SV�0v!ͺ���]Hϱx&#��b�A|z&��N�@�o�e��K��c��X�g��G,=v��c�9};c��S0��,�<�����mŲSX`�|x��$U��#K�t\��t��Y[� ���u~��$\p��!�*�tN$f�pWX֬�Ӗ���jy~�f1�҄Z� ��E��w;aoc��t�����޲I\��=�a*�N~o�a�9u�uJJ**aEj�c�2�}-�oG/�Jf.|�5,���P\
K_�:cR��ԇR���2?[cPF���!�WS�/1���e$� ���.F[8�t�Y���!zKu�m�kǚ��#wֿ�n�kF�g7/�
�	�-N�C�EY��DP�8C�K[�"���z�Q�*�j��Ƃ������l�ڒ���{��羾{S�½ݱ���,*UmC���;��}������ڃ-��Ӳp��vFb�����g.�r̃�iw�c�P��='Y���{aJT�������eu5ʘ�Ei�)*Ѭ�R�6~�'����LzOEU�^��l�F��Sp�t0=!�<�����l6�E(w���(����-E�'j�5�����"������k��䗜YX�����|T�#9-MVa	6��k�{�:���L��b��}�Y�5�=�s������78%�>��ā�5�ST�ڐϳ�I�)`��=]Y����`l��e�A��ə��������ٍ�h'*�2�J�lSc��<q�ݫޙ6��	d�Jf��������=�R�4��	�9VOmm-I9fA���*!��YV��pnJ~a�^6��8���+(y�$E�xo��2��%�ESI�p���B6��������)�ˍ�\P�rq�f$]���e2�"q�.��-�zEjJ'���
��U$�G������������ o칚��9�����Q��ـ�� �`�|��>�=���c₻8�t�IfGB���2^��g��i�X��w�Nxvt_6�0�.�����9p�ց��F�*��{�s̆Տ�r8�d���Ϛ��iY��>;�����T,&�N+�g��A������ .�s�/�ߏ�g����"��Zp_~<s��`P� ���q��b��ԭ���cyʪ�wq)�-���d��tӻ��ێ���'�i=���iu�4(��]r̂D®'p8GH�R>��j��ߪ]���E��78��o���Z,��G��!��y?od�2�c0�w��S���"���Y]�|�ؓܮ�4|�9Vj�F�����������ю��.\p�X;��w�Y�Ie�C�w�cV��G�7K����EM��An�Eak�u��*�
���z�I�X<e8���ښ=xdpp8m��i���r)j/<��^ȸ1����������傻X�kj�w��Ȑ���Tp,GFa���u+θ�A�ǖo�����"�B浍��i}��αn
�~��T¯'��"�J����1���0��vϏ�Ǌ��� 9�ol:��g�Altj�y}�ࣝ���(ұ<7&�";��͙��φ�,EWL��K���ѐ�JCPgwٱXV�V��y�?4(
�F�a��r,���=�q$1�{Dg��o~á�-%��3ƛ�w�^R��3$��p�8��Ql+�6P\jEo3�(��΂��Yu��F�u[\�M�K7cÓw���4��� ��Ta�Y�\p�:
��l��'ȫ�q̆�F�K�s��ߝ>!��x�-XwV��`�@�xp*ݝU����t�D������O뉷�e��;bt���e�ֱ�y�aق)xa�^�,�cy}��ߨ>:�)���)�������ˬ�Q���dpw,ه((�K�܆���IV�����mj�h�MHl�������p�2
n��*PpE��#�����)x�Z�~I�2U�vǡ�T���)�3�]+�#�e��&뙸웸�����;Ǫ�E��N��Nn[�ʘ��=0E�rS3�=��k�	OG{���{ޟ9�3p.5�fjT8ޛ1����E��ӡ�X<�±������D������ƾ�6恁�XØ<�i���$����C�U�A[�L�v�����9(����\n�ߗH����p8�ù5�/f���x�q�l`j��{�A��#�}\�P�8a �l���o��N�TӁ�:�x ��i��αj$�p��c6l�r_��*(R��;Fh����	�v62,_0E��Nޑ$��H�xm� ���oX:�7�V�S:�z�4	�K��Wl/�š�X(���`i֓�c���>�����	!�����yE߱>j��'�˫�y��Τ�/���p8�����R���hļ|?����w��ké���$п0�:��d�>�vb�.�>}���>��E�＜ؤ��� �6y0����e1�V]�B�p��c	��V[[���QTYUU�%�e6R8H$R��N���Dg�pq;��i%���#أ��%���j�/O�H/��Q��q�X00�͏�ܞY���4��li��0�%ڍ��G�FT����� �����z�_�:��+�y�$�O������9?n��� <2����!ʫk��`i��h~��F%ߛ8
7�o�fy��/��`�5�y7U��7�Lܛ�>�c8�v!�����p8�a^�p��������}�aݙk�p{�������!̖SIVQ)�;pb�Y$��%�^�C2��$��}����f]����xu� ��|JJ*���֣�\p�:7�+�;/^c�Ϻ�{P��Q��ᘃ���%䗄�᣺��i��t��PF����҄D��VlS��EI�ի���,E7M1]]p'[����y��˶bz���{w�;l@��:���V5O6?��3������v�xa���?�f,݂�I��4՚��c�w�w����S	�ͱ�i��N�k��ù]Xs�^���1Llz��O��òg���=;���X����צƠ�@��1˙���XX.��~�?;���.!l:���Ow�`��/O�l;��"���F�X�Q+�z�.�s�G��es�9m���2�B/9�l�針Z��(,�z�8��&�a����Wc�z�%p��<�r5������o�y�1��~��n˻��oM�#���2�&�����~'�y�fk�u<���,GMp_g'���Z��Y�%���i�|y��IiR)7q�p8��ᘇw6At�t`�d��`pw�;��A������3W!6(Hg�7k�hD�2q 䲺���v��4E��t�<8-�9V�����G�8�@��n�Uպ�ñ"�K�5�S�ؿ��9>�����i�l�	��]�3���,IqE�Ƽ2�}N��,RC���|�I���Q�XB=-{,�Ʈ�4-H���ضp�jYM��<�w�hx�[�^��eUU,�G҄N����ENI�j�����_"1]oW����p8G<��o[�빹�uih���i[迲`pSP�3�Ot�F:��?A�.��6�g{N��-�J�5��;Ǫ��Iy��c*kj����α*b34�Z�
J���A���jD~ڏ���e���ய�jk��N��n����a:�R��S+w����^�Xl-ۼ��)�D��QLi�40B����j2�����
߯��<��Z��̞��+�m�[�7b��4���^�B*����p8��1�ť����!�����{�"&� յ��^c�;ه���8��9V����9桰�� ��q&%Kh0���ف�����`A�gW�f1%.v��,�Ix659±x�I��L����ζ��?�k���y7���L�j�dw��ģCz����lmd,Z�m/���	YAU���:�%�8�ޫ�,"�R8�m���>�`oC�|텫��%���c"B����1!�&�^��-W�Y��:����o��oN�{c�~�TV�(&�߀5SP^��Һl��c����e�8�'48Wc ����V'���=+��A�0�II���
S���Z&ͅ�w�>.����[ӆaHx`�۽9m(��
q0.b����=>���'��ĥ�\�q�2D����k�Zɱj�2poW�Y�-�,�ceP���#��������%G/`��8�eNZQ��r`I�X~����u�b�S~��k�x�Ѷ�9a�b���e��:PB��!~z�E��#���$����gc���0.I�ڷGO���w��,A�����_�=���XF���j ��2k���1�c(��j������b�鋍nCY�	{}�����{��[��%X~�"6^����Y�+սF������09⮨�x}�f��ck�`��+���Xƿ��ǿ��m0����瓍nSQ]�w��R�鼹�ٲ�G��`�1F�-��������]±b��Ϩ��Tj���ẗ́z�!����|1�S8F��7����ُH)(T���8#���?�~Z��)��:����磪�&3�lڅ>�~�}�tt��4�3\O��k	������v͝z�AX�%�p8c�)�����JhO(�j��A}�����߭c֜b$��k��Wl'�Q�,f��f�8�����%pZ.�s����.9f!�����X%��=�y��L<������Y�U�t�
}���6|,�����:��#�)��*�6����r��JHL��;1���(�4=�"��3vH���DҼ�����+�Y�Y!_�O-(�ѤT�<S�F<�c(^3�:�7�9�Fd��7^����²�Kt�!|��X��D䌢b6M��������@7u(#�V?SI�f���QXQ���VUi�8�����bt�����l�y�,���i˕|��(�<=���Q��Cw`����3�T�n&
��s�Z��N��g�� A�K�������5qײ��V��z�����p8⇂?>�k�F��K����;�����#���a=Y����:K��	���sĕOY�K�?W'�2���|>�u�Yv.���V	�t���jL�&>;K�R�����αj������(�c��TT��6`��w��X�PCj��UH�PC�ѶAp�|1��$��WTbΏ��D��,�߯�5)��E-��cp����R3ڠT�X^p'�fǣ�0����*6޲���+��D��q��ژ�R���v��n�����Q�ӆ�[E����7w�Zl�S���o�����!_��`̵�.�p�>u�7]�ǽ���#n��1g���:L��.��{�O4�D׮1�����
�hՑP���;��U�Y� �<�����i���}���p8�3�o�x����,�p.�l>��B����7�O����ذ^Lp�(��ǔ/W���d.���uY��L[}�*>�sW�jc}w�,~���cCz��Q}ر����s�b�Gˍ
��R�ñ,Rp�D�y�-���ñRb�s1t��xy� L��,J�Ǉ~ۊ�b��I%���J������X _�a±<?&��c�r�Gb^!X����ڸ�YtPd�K����x8��;�R$�;1�} �?��߸����*Z������w'�Dd���X!Q"�������/�����{c"�mj��N�;fܵv׼�{�̬�����6�
�[�ˊ����1U�5����׮���v����=#U��==t>�g]��5�
���Kx�U�ݧ�5rk�����2���F�|��A���j|r �ñN�ދ=/�>���E\V����ۛc������јۯ+�C�0'�V�����7�/ˆ]�
�R�Id��ٞ����y<>�'��� 7g�6y0^X��������Ϋ�q�*Jv+�,W�!Ѡ��g�
�P����Ϧ���o�e��17�!��������Q'Gl����	�͝�7��g/���$V,�</۹8���/&w������*J�<K�?�	o}o�H<5��

����`��=�:o�:���"�K���un*jj��_�c�A~�Ay��I_/�sͅ+����F@��;�ͅ⽖���������;��~nOw�l�@�J��^T�z�:!n,�Y8�ri]���\�+A�}d�l'��1�G[�}R�_ɬ����TP�&G;v����8�����Ƴ-�^��2�lS74�!��������wV��w�pJL�#k��rv�����د)�{y�lC6Bڂ�v��;�G��dG����5(*k�o�����Z���¾�z�<��Cgݏ1g�V�;���p8���L���p�N�Mɂ1$�ᅿ��������^x|XO�y�(����bYL,��w�������<��N��G��`���g���
�RM����n��;綁�/7�*� q�����jW�2,]败!���=-�T*S����<("��({D���z�ek�'!Qg[�
��`>�6^c�_�����A�~�<�����g�}Ԩ}��e�^�����ofNdQ��P�A|n>��N+,�+88i��Ϝ��Jl�zCg�ѧ������:}l�f$��
�	/>���ư��n�	|�E%t��^M`Ec9�v�c'�u��cOޏ?���tMу��k�Ա��)WՆ���5��OĻ�aN�����%Ȫ4�Y��ͯ�;��ߗm������%(��c��|`���p�ORn!f}��Y��E�����,A?�pB��e�Q������X����{�s8�PRRZRPXXP\\Z^RZ���;9:������f���:I$�}uj���U�{�յ5�EEL��$7WW��L&���8;ɤ2����+�7+���1q8뇄`S��%�����7��1�]6R�G)E�oZ0�Z���:�/=y�O�!ȵ[���Jv��r/G�<k�^1��0:�x��T�o����[�N��]���?�8��|m�U.��"ڙ%v2���Zu�Lt��'묋�9���n�{Q����殃�߯���C�F ����m�Z����fT��w�Ⱦ>r
��Z�D��'�[�X�����X�,��p8-�9lIxoKPfcR�H��wǲXk�29%5y��݉{�DZz�GiY��B����Z/4�D")������]\�J���B��l;m�$7G�a��<�[�fE�����������Ds8� ��㺄bbd\H��;[��vE"m�z�2���5����5���Ug�Ͳr����:����:��+t���&�R��!+��jr5�7u>#�EA�3 8c"Bu��c���w�~�>v6��^��W$��),ohw�;س�%�WW�W���/!�M��W0b� �:�@��n������{�� [~YC4�{{����=�� z�/̫3�S�]M�1�M��ث���vv����]�ѭ��eչ�Xq��Ȥ�p8N��n� Ϻn���\$�p�]p��o��6 oyrLBh�V��'��cg�.�6DV�J%����ń�I�u&UͪeA�
���+�k gX��%E?/]q���������(,
��"�n�{UuM()-EFF6N�>�V~-�<�����]j��KF7���R/[{g����\�a#�� �Xl\�˪kTҢ�}X�I[���?vb���p8��"��S��c�0�j�P^�yE2�
�V2k���O�A��_�6GSZEpߗ��w��Ȏ-��G��̹P4#�i��k:�F���¾�P1���I��9��#��aSѱ�ib�cF׎:��v"YXi�j�2���-.EmW_A��/.6RvGQ.U���%煶��z��{���b��X$��Tm;�ow
�Ф�N64O�ߊc��{q�nV�x~�(<>�7T��=X�~�\I�[ㆃ��p8�����70���j�q|�F�Z�=\����!�i7r�?.���!�f����"�X�T��y����\p�� ���rL�Glml#������-vJ������l������n�W�j���mk҂�J��`EU��յ�f�����J
*�����LϨ,-�����R�PZrDQZZ�(+��-+U(*ʥ��	*�m�P[YaGA䨮���o�ښ�?_QK&V���	=�j� թ�E��nH/��iWb���ld�^���v2i��ܦ�A���FR�bk[e+���P(���WU�0e�R8g%¹S��/�T��eU��U�
��[���r���^&�t��X�M��w�Ihq\C
1Ef�:q �9�����������O7�Ě]Wq;#�5/½N�3�]a�HdR�p��{lv6Z���Wh�l%z�����l)�ِxݜ�u����Q�!�tG;g'dk�Z{�J�����\�]O²S�����oMK�TfAw=Q��^������S����q�oWg߅X�ׇ��j]\���ښ(��l�R�p��&�g,]�Z�Ɂ<>����n+�]�#5��{�nܡWlW���W��Ż{aAt<38ZU��>�w��9Ȋ��箨.�p8N�)�j�uu0)FT�P���'�D�g�CnG_�����ELb:�<u�/$`l�&�Gx����t�E"�2�ۋ�G&�����H���2����������ǳ��`8�A��᎖è�}�*O),k��j�����^:�j��V��p� 	:�!~u"{TB�&��m�+�TZ�^���p9�^����(��YT�wy������[�`�;��h�I��XF��2�}@� f#��:a���Z�;km.ef�ǣ'��nh�X�F~[7�syZ�\���/�_cE�����ܥs����I����
��5���W���V��1=2CB�p�F
�'��I?��QC��@���&�4���s�����rPq_��ᜒ-ҝݺ��#'� �dr�p��p8��c/o�psK������~b�:�L�ϦO����rfĊ����k�~~�_�n2E��T�]9�P(B*++��r����55�b��q��9��mu1=��H`�D�)Qah�j\i��b���nw��nb��$;OVŕ-_d*�L��� 7��~5;��bx��j8�K�����ֈ�Ӡ��H,eH<�~���Hj�r��sJJq�F2F�Y^�6�~e!��� q�25b�rX1���\�����ͤ��v��=��s{t����5�U��o��ݍ�5���_a2*��_�����ǡߗKT���b���������5&�S�������)�����x��l@���g��0QqVuhww^��&u��^<u�ڲ48�8�5�Pd��C��t�X�YX�Ҫjt�j� f���F��5����z8�Π��vZ�����B;�2���u�1/���><MC˾�#L9�i�eR��I";>�01����g����-A-z�)��X�zGu<[!2��@Q��
��V���W���Y���B�鏀RG*m�wS×�_�c'�&���>�M����T�������N~�]0Ζ�|̿�>^g9YʨC�u��{�tz�8tBc��g0g���?�zO��ߴ��������a��Ѿc:�^�<���zt��`	�3�1($O�Yݻh�}}�0�:z�.��kt��^�d�4t�����pn5��[�ޝ5Jg�Ҋ*�^�_��v>g�2!z�­������[c��)���&�~�>ŧ")����[�p��"�;:(D�﨩�m���p.5C�����ƨ��ؾx�	p8��t��Ċ�\O�'3rY25���q��Y��%� �fF��*�W���˽�w���#Z7{�����N��TK��
�r#�˖j��\S"��+p���C��3�
�����I%:�.�ᳩc���Z��ct��{K�G��;����3a�:�"��f�r����S�"��+�ƪ�o:��ǎ�'�ߵ��3�(�櫪��2zw�ILcYJ���s��k�1$��䢇�'����R�ӝQ�ٔ"\��O_��ث8����κ�x�������pnu�vW'UUcI�-���-��j싽�Ub;��B����c,���G;��{O���n)ù��ADFmm�9f'��on>�&�c}�	�'����n��I�����ŻO�Z�M����`{>�u\Y9�S{�|x�>���G�oCa����ۍ�f��*��4���w]��>��4sA�r9�xV��d�u��"��r#��z��@��t9^oT��;����řy��w��=$��dQ����6�&��k�T�?�N���.oj߽������g��םl��q��*j��;���������l�Jirs����P&�8��CT8�L��*�X�t?���l<�jV���VΛ{[vC�C4d)C�}G�/S����FbSvI).e�=����p8��V�JD6@�Υ!��T��@���T�}��xn��C�pK�Uc|��I�ȓI�7W��\�����p8�6I� lzr��G��+����?o�i-��"��d����6��&�PB*Fvf�Ѣ�}��֣��!����oNg��@�*��|%^���-�@Q�%�i��
,��o1�]"^K���5�>���.�/�p)�$�]"�;�Զ�H�puA���btD��7��B�)��|F��:��MHbES��;�e4|�d�J�`���y�=���3�]�wO��Lp7ܗw��Ū�w0�y�4Q�lɩ�2�~��89§C{p8��8��q+��]`���觧N�s}�fY��tK�^ �����m��2�r���5n:K����p8���g��{M˾�7}�_���m)lx%��"	N���_�},��?:�|�9B+Ej��+mFgȐ���o�+�w�tGt�?Z���'�����I�%��p��p����k)C��mW��V�p9/�N�1$4K�L���<�8��<�T����dv�o��l�H��kJ�����E���z{�B��66HE5*��[ʨ�,>�$оNpW�/�K~�p8�!*�� ��e�~�!��\XWQ��s!65bBݟ����8~I��E���#��J��3�G���}q97� ���_�7sP�Vq�	p��c���bC�Ē�|
���p8NTi@�a�� 7g���}�RВ*ND�'�L�;b��_�H?/�<a ��"/I�~L4��n?8�Lb�s��MmK�|f�vl��w���{6K�o����[���%�����q|�5�Ġ��̸ﲵV��[�w;E���3�KXFBcMJE�����8-�vAW;�^_vSQ�q?����%�`ǵ�()1�S��u��&=|������������5}�����ES9�c�,mhG�O�ī����Q�b��P>2��P�샃��/��_���ȦQ��5�ߒ��xA&�ũQpw�큷\ReZ�o�P(��;���p�M�2:�b*�1�g��_6aj�0L�� �WC�丮�lj�B���g��W�����"��U�#�<���}'�#e�!�va��:��:�����y�e:�H���/�<��=B�����!ۆ{y`|�0l����9i�E��R,�3���"��	�����??���:����
U��pb*��`�F[W�3G��gN���0�}i�N&������ENKN�;{a�%��GH�|%�v�Y��>�v�XR��yR��]+�y��~���Gsu���D{��<.\�J�}@p ���SR�!s=I�����ac�p+���p�Ƈ�{�Z��W�H�C�8�IN'e�w���َ����ljHy�T�Uc|����-�ah$�y��p8FVQ����1�U���x�9�}�|1�M$���̞��=�E�7��/�V���T�:��?��c�_V�dj퇓G눭���q8�h\��Ͳr�:wIg��� �]�7i @_�F�G~���C1�GWd��鳓���������+xS���
�Ʋ��l��ߗҦd@p 6�?������ަ*���9������ZP��<�cfd.�� a��z�g�4\�t���IU<Uu��.w�9Q�{1�%���qR-�]��n�ñ
�]J�C�z��)mBpo�@"K!�J��αf��p���`$�%-e���é�������>���?���˙y��O$���Ʀ���G?O��ё	��y|��}����gp!-�7��1dRӛ���u?W�O���}{�_o�搡�����爁x���)�bW�6�C.��P�!�ؔ�0����Y9����Y>2��^����Q���ƴ_W�B��l�z��հ��ݠ�@a��/��4�6CO�Wp�pӘ'[�ϭ���	�vn)��p8���kI�IHE��@��[��~0>�����\�m�ve�m���b���?hyK���n�L��6���p8��Z������Jf>,�K�^��������c�����%��#	�/��{�l�mM3<�me�o	��Gch��4����4f���	��z�kM�������`1՘������+��0�����ѧ�ǌ�������J�O¤�a�<��`�]t��qrԘ���{{Ga��˃�]4�pjEsw{9��?ӝ��pn;虴h�6�x|&Rr�_p���9p��ok��pڷ�̕� \p�p8�
����z���1��3+�əX6�Y���k����/_�;���cb��� w�/;:�������������:�xaTx�v����|��-��wZ���3�mߏ�WX��>�l���!���>�Bu�i��[�m���]���q̯�1ڻ����������呓*K��ႻuA��`77$�if:�ws�����\P�}	�l�~;����x�J�e)C8��PX\���Xم%���U��=q"Q�w�UcJ�;����\�YL��H$\p�p8��^�J2�����j콖�&���
�f��4�ނ��M�F|�I@���|�e8�ڲe����'��]�.����yw�
�����yw?_���O��#]�8�����+���w�&�x�7}ޛ8Ҥ�+��DU3;�o����XF�`����5 ��N����>޸�[G�n,4���Աxz`�8��I),�]�����P�AAy{��	�i�����e�?~/*j��w���h�+��ox�����e��x%��v��m�I�8��|�_���D�o���ۣ� ���"�v����s8����)0����Ýc��^�P��bWpK���AȻ���S+�t���,e�\���4%�� o��)�9;�5�h��"��AVK�ϝq����'^;���0��rsEK��c�L�y�"�dSn��;gO[t0P̵���#��>h��p8Nk0��u9�����ۃ�Z�?{�'E}����z�\�8��{��Q��51�$�1!M�ƨ�h�&6����{=�qp�������(p[n������g�c���������yL�s�ʦ�j�ڽ��#5��Gñx"""""�R3Ý��^�2�cI�DDDd��n���
�Yp1����1SR��������p'���M����:�3܉��,�nV/i�7`�;�r�����%`:�]�_�j�Z�V��� """��WV�g��'�r�Z""g��k�y99ށ����Rp'/Qg�z���*���W�����DDD���|��0�����H�4z�p'��`�N�K�h��ZmMe�>DDDDDDDDD�\z��j�f��.�N���k��Tׁ���������M�60�Nޡ�1j���htY��V�U�hp'""""""""R:f����7�m��OT�o���������H�T`�T����u�e��������j��d�z��\P�ew??��԰� """""""""ecw"���z__��԰�S """""""""EcI�*��h�i��%MS�ה+M)�!~ """""""""E����N�Am>��w�<�"%�קcT�o�Ś�X�2���gQK����b�S��T��@���S�����t:��+�0^vü%�R�R����d��HW�I�����0i���^�S�b��#�Zw�w"""""""""�RyB��K/��^ 88�d@@@;x��K�_,�����
� �Z�1P��O��/O�)��l���������O��[�D��Jzaeҟ�e�Z��WK���F��I��		����a�Ƿ�����~��j*}4*��;P���jT��hk|4j�� u�����A���F+��U�|�7��P?�Fe�[��4��5���N��V�?�o�tz���u����gf����y(�����{����4�ml0U��F#��:��t>�:��SY�2\hj0|jA """""""��xH�{ox�NW/y�M$�7ɧq8��>�J��H9)�˕@��lhh�r��'NDJ�h�*g���FΥ�`u�g���A2hPo��/��BA-�֨u��;4�Z3�j�*���FZ��T�V��5M���O]@@����_�/M�+���s��8i��""""""""+�PϦ�J����z�H��	"�$�#]��2HT[[����k�t֨+t�c�DDDDDDDD^A�ew����L8&"���P���������ț��*��J�&�n4@D�FT��%"""""""r�V�w�6�j�:DD�@�w"""""""�+T,)�(�!�w"rr�w��������H�we���/�j��-�Өa�DDDDDDDD$Q�5�E��5���M�Xŝ��������'�:��J�*�������w��G���������2�
@� �	���aw"""""""�Kj�,)�(�!DDn¨Ri@DDDDDDDD2����KxU�]�
DDn�h42Ý��������2����
`4�T*K�����p'""""r��@$�A�Q�bU-�ʪD�G���3�]iC�F�a���\N�w""""���a�12=	����*$�ۋ�k��ޓ��}��ׁ��Z����w�1��&DD.fTA��F����܋F�B��PąIS b��s�o��*�P�ף����ոPV�s���XUj� i�&G� E�����+O���֡��E�2Ε�uNI�-�I�_��/�TH�^u�ե�z�N�нU$���'����D^y���e��< �=))�tY/M��o4�zi�5q=L]��hZ$�/=�ALM��������鴥��C�����������*�J"7!��z��J�W����L׻�G�_j�4�KG�ML|5ͯ�'��O��`nv��Ǯ3�8UT
�Ix���MD�V���	Q��.K��l��ʻ��9Ҕ���P�༬r�ш�@�&o�a��4�w�DRD(~;�����%f��Z���N��Z��/`4O���",,,��ǧ7��\̈���5��V��3R�)c:� *(�!��������C���׉l����b�4�8rƩawաU$n���;��{b�<�a/�Z���0y�ܵ�|]�N/��;�E�p�bɚ���gϡ��9TT�b@�^��=g/���Z�Z�Q�H�ה�Q�؜������H�z&�➾�0�g:��Z�9Ãq_�y��k�����v�1�>z��&N�����u�����"�)Rnj�(O�'�|��{_�:���Z��o0X���9�	�bC���ODD�Q�(~�5w��^١������HD����5�z%�r�k���k���r|�-�o�����}[��AiYO���Z�欉�[L�? s���� ��E��g� ɥ����4�̀;QKSU3� �p'"�b4r �����	"�~���xvd/����I���&�s�z�m����}�Wp�ͱ�Z㥛��[b܍hx+�0��_��k+w����fϧA��K]i�۔nұ�|.R�c�3�ND��ԁ��+�7�W""""""�Q���=��I��w'�ޟ��9��k����J!���a�@n�w'֍)���5�EY��/���A���j$G���=#5�)�h-��Q����z��Pܕ�5܉������WǸH���������ώ�{�e��K��;���K�����<S����J"^��;`B�4�m�N�{�~��-���R�wᶑC���'�r�v�DDd�<��i�R�F�[�Ǉv����n��b��Ό��ѫ�����J�n���	�2���P����y�`9���V���2���t2�ӓ��b�A����`���y�@_$G#2�a�r#nq裕&�h��Hۉ�K���:t�K1���(����T�Vס������T�����.V(~��5w�%e�Ƚ�l�LDDD�M��s�XKO�'�.����a>�r�-���a�x���1��j<6��<�`=��}��}�J+�x�qL������+ļ=GP\�9q��Ix���F�A��� $��\�;X�;��N{np?[R�3�ҥ��q��E�&�'+D��^�>�����JD
��!"""�U��X|q�x���'�9_��&ܜ����Y�.l�*ʯ�7s����D-��9Z^�~�h��LԦ���Fym=�to��h�s�\!V�F���@D7g��E��kB��E�������"��;�����](����"��)���<��:��� �V�R%�(%"�`3܉���;M��s���2��!럝�{?[���[��E���ů��S\�v[<:�:�E��O��AuSvd�aO���
����u8WR�������xn���I���*RpS���@iJ���g����{� O�ǏG��/�,c%����]����$"""""r����o&7���!�X��T��`>۞�"���+g}O�orS�D���4����9�@d��*,q�s�zhj���&]=H�����kp�~����:� ՞?h�J����&C�$`h�t�����C?�R���ѽp��
?ffc��l�?���g(�����5�-;��PI�)~7BDDDd�'����&��{b�W�j4x��H�
����,Ƅ�`�x2:�E�uM���'o��9�[Z��ykk+�[Smu9|���#��#]����Z�?o���. u�ahE}�t.]��j>1+2�o�H�M��vu�0Jk�P^S�u窆4��� _�Ӳ��Â0k`gy�+���v�w���
x�ΙF̅�i�ju��`𖀻Nz� """"���l>��^��M�^�� ����o�:���_��5j�ٌ@�9h2F!����a-��F�}?�Ĳ�1m�r��A��^����*���.�*����K�J}�o�z�9\Z�-��oG��7�������]c�ָ�ZG��G� -*�Ll,zl&����L��JٱP�&	��y�++���s�'�.$d������I]�0>��������8_Q%]���ty�����r?���z���(=uej���C��B�}��nR"B����K���*!,H�znTO�;���ߏ5'΁�A�5��=��^_��������Y�9,�5"�� ~d�+o%��h��x�VƋR	%a	�M��繵G:ޞ1�E���T���*�V���F����<�#�v����j]��5�O�j��W84��9>�,��q�M.�yQe-*j�m��e�/�R"C�L���&:����Z�쀚):� 9�����c�ƞJ���1Y���bs�x���ɼpYEe�..�.��bN_,G�{2��v�/&!�Bq���[�%D�S��Vк��T�9D����$y�y6��ڍU�r��f�^Z³�d^p'"r'F�cHDD.����_e1����g4�]s}qQ!��1�D���9z��¿f�rzY P�x2N�����w���櫊�h�H�G��hi�Š6	��"S�����x��	��I��܇'!<�-�VZ��O���\쑖���B�Tך}�(��~�q�6C�&8=?#>
�33?��������rZ4�����]O���K�=�:bBF�������e�"��)���"��-@n���^q�s���43[�������r6�Ęf��J�ӹ�&`��^Z���\�gR)>Dk4�j+ �_������{�x8L�u:�m_�����5Q:�����9Y�"�p�|��V9#gU7���{<�X���}\�N��q�Z�Y���LӺ���0�|����!2�["�^YW���0�ql:�'r4�x���O����c�u=�cq{����#�i���;��᷋7�5Ce9�s��Q����>A�]��
��}w���wG$G[�8QfSV6J�qy��J'Ww�͗����#m�0�K�ѳ���Y}��[�n���T|�#�q��L{r���^�=#o�!!"""""r6����AG���m�E����]c� ���K��]�0g�~�w����g�3�)=&���g �Gg��3��|��`�����`����� ��}�.Ӱ7�@�f��w�n���셶��p4ѰwKV�>m�<�Ņ�1��,���A_Q��[��Q"��޾1�}�UY�b@o��\l8����w�x~	<]AE>�zX�ҢBqw���&&��~W,���N�H�oo���'�!<"v+��&�NDDDDDD�u06�C���������޸�]"MdX���-r����(,��ně�w��G�tsJ��SҼsJ*����z\|X�� ��5�%�ӏ��á,��(_�8�/w�3�EF��3�ߞ1{�(�Ul����G��șD�!C��m!2������� ��?[\��G�bYf66e����Jԝ��x}��ڽ���2�"->N,����m���x�2t'�VÝ�F"rF0=����ܓ�rMq��l���c�☾}Mg����7��R&-���Z����<e�\��^�29%���p�U�������u�k)����m�thSWk��3_�:���N㥛���A]����wf���.���ƪ
40�E�T�<?;��N�"��M�p[�vk�:fa��38|�"�Z�T�W���=�1�k~5�:����8���9>
�}�ʫ�`����;T�YIDDDDތ��d��R�Ci�!�t��o�In�(��³�ֺ�N�����rMp�ud�T���q�����B#<���s�Xt�"����7 �ܵ��k�����)|x�X�e��N���Ts�+Рn�RT�W���&�/���R�^�/�wNI߻,�(,Y&�z,��ǋ�����w7���9����Ǻ����W`WN>�3;��J��������ș�����ExxpW�i��!��>7�\jĝ�:zC����}&tv\�f-���x�~{�\bƔ?M�q��H��x���Σp'⌆���->�k��'9d��N*}�9r���0TWA��8n,�<��jq)n虃܃������n�lXVQ9��=�OyE=vg�w���P�0�?f�lvp�Uh ><w|���Z��0��ح����Y""""""�J�o��� 3,�/�uL)�����;*���=�.�#���p�c���n��?�����GMJ���O���$����x�����>��{3G㶞�v�O�����xu��f=Ψ��|�/�L2/�O��Pi=ke5��:e0��Mh�vq�w�O��='�����~�&Uux~�&�x�>�9������`���åؖ}
�k�We��o�4y��")��I������ܒ�J��f�����^f� �A��s�P^ܙ&����\���n��;B��h�u�<���k���7��#�:{w~�T@pg�l�G�\���Z�,
{=yS|��̷���z����s�s�/G��u�pu�_���zC�0��aձ|��8�9#� '�Y--�Q�~�/�'��7%�G���	s�%}�e1Ý�����Q�!%*�=��������F��?����nv?���`w�7��xƽ� s����`��sF��ؖ��O���-�����6��ç��W4�I�DiQ�F�Ra֠.v�Kd�>3�'~�x�Տ�:��+�d��p9�^_'�hP�ԨP||�h�L��������]G��cJoҩ8�Ҳ����r{��X����"0?�.��q�*2�p'""""jB�����qX��$^Y�D�B��L3FhDֱȨ��yF���Rl;����G.\Ĥ9��iHsL��o�n��["/�7n�Ԩ08������W��J���7���,FuH�k>���k+w�Z�!�z�5��gq���_>3�ji.��MBL�u^d�/9|��8��r9��B�l�[>\�E�LB����&����?_���K���J��s=�4�������A����S��#gBz4#+��n�n�g��h_Ʊ��r��Re_,�K�,y��N��D]����/��t�.�BdͿ��z(5X&��<��2�v�D�>��{�g�_��Y��A/�X��q6 ����˨����qQr07"�G�K���#�f�	Wׂ�CEm=f|�˥}NZT�����h��zw��v��3�MS�h4zćFDB%�ǭ�����C�`���Aw"+�U�ܧvk+�����g�ջ�tYEe���"���4�عL�-�+5���=���W|f�h����V`�S��jX��.xo�>��Cd�˗zB��/@r��׍P_̙9Kg���;���Sae-��|9V=u�ٳ��8q V=#ߟ�O�MY��{e>Y�A�~*U�ǀ;y�妩�����OG��O�v�:�F�'8�_�i��E�MET��AwGY�yO|��c��ޜ�c�n�8�����0�k�����߱�23J_��d�'|��������/��2/ㅅ�����M�G44aT���&�3XÝ�����#�H��&�7��2ܙ�B�g�ZpO
��v�v=��V�@NI<I���r��ŏOsh�S[m=���X&�cq�{�v�3�{����:�����:���k��:�o�ۋ�Ŏ���\�wI�/�C[����r���w�(��2zDL���hT~�M4D%e�b&tNń�T����G��q�S��cK�(��(ơ������̋��D�/3�ɋ��W�cB�4��8�X�`��� <��3��6��G��u�V��ϖ��pg�CzL���|���S�<���_�mǜ��m���m����2�Z�U*1��5�j&V3&g�H�� _��7�0���E�12=I��_����[�nK�w""����@""wu��
���"Y�x�b}g&���ߋ��%l<�g�3�%!�����q�g�PXYO�������^�i��Eٟ�ɱ�m�N��� j�Q��Br�����̑��o@��]���K�t򿷜>�������G��`�ٖ�F���3�v��C�ug��TbΦ�xvDO��������e;�6 � ���DDDDD����ސ�Hi��	�p?��I����*k�ծc�t��~:�����-^\�{r<���L�x�!�v�M6�ct����4r���p��O�)�뭯�.��Gd���v�&l>�r<(�gP6��Cgh:�mt�|n,K�i�T�;��A]d��Px��tM÷{N��G��h�&�]4�Q��c������+��6T�cH�"�	&��`;��w�wβsH�������;�b������b�x�o��&��l1���i��2ܙ�Nf�s�����l��0?�s�2N'ʵ��4����4}lZR]�/v�cC�����npw��f�Y\�������+�`�G�'�6�h>Bзu+��k�,x����׫0��-R���b�����e5uXr�4n�n��{&�@�V�^���RK���8�� ���R�J�84�(��c��vd���j�$7�=0ܐG��,)CDDDDt����Z�p��?Y�x}�X�d{��|Y%����R'�[{���� �ͩ�#�=��jw�8ͺ�gm���"=6B�h�J����%e�wNkUrέ�b��f�,��l�l��~��J�G�K�?�����]�&�����ᆔ��6�Uwiâ��\Ol{�=""rS+�������U���M���Y�?������lŰ�$������|;���ۈu���cIR�6ѡ�**��:%osߜ>	a�&oO����۰��R�$}�%U�a/�<c2�.�Omŀ�i�j�G�"""""G)�����>j��{4'E�ud���s(��HԬ��UX��t�jl�oʶ�yxg�^x#q����r�ظ^�E�@bI����2�T�_���Sy7ܕ��`��7�6l7ʪkq��E��45��p��-�מ�ŋ�{���[��`<�O�e%e�W$""""�j�:��������������}�k���[4�K+A�	�Vf���A [�+��>�k�MA��:'}�_^��a�;�[�w���/G��#�`��߬1]��3z�c|FZ����A~Z$��X����탋Uuf��ʊ8QP
{d]�=��m.���o�7�Q��\�~�F���ƣud^Z���
^w-�vw/�cˮJw�q_�O��4>��^�h��Ps2�� ��ew""""�k��l"�t9�(�J���c��~�H9wff�%*뚦F��4'�`��]ۘ&8R�b��ı�|}�.�ң���j�Ud�rm,#.
Ӻ��{>C�&Z��������)�=�7��:��<��Y��S\$�?4�a��`�AT�7�p���r�;�S�)�VΜ���Ǹ�Q��˖>��b����m�8C�ɔ�A_��k��1�3Y7�ț�9Z��k�u��f"���������O�Y��.����ǆ�[8cC��gxD<��E��e��M�3�C�uXd5��t����s�yR"K��RC9e�&�!Һ"��asm�� ��m5��"""""�"�Z�L��3�=�Dl%�"5�:�˨��5�s�`�	��#ݮ��������׻]�ŉ�[�XW"I��}�K�÷�& �r��׻�#����n��R�����.9����|��0i�W`�>df�]����^xD�N�A�^�lD����}�n��O���R	vekj��L6@�2�#����_�W�5�O˶�Y��f�_�Fg~ ���-����AZI��h<�4��������L��N�=�t�4�,���~�����=���6	���9�vv����P�)1<�=<�?��zs��W��J��@_-jt)[biw���I��L�c$<��+�±����-T.Hq�t��N��<<�i*��W�Y"rk�!""�Q�T5������� ��m��V�ƴ�Q�T��&bf�v�G��xg���\�<h�g�c�>q���i��C�����q�	�z]ni%�l8 s~9�'&wI5y��~܉5'�5y��C�at�d���KS�债|4��Ax�?"��_��w�u�D�+��-�����X�=ks�)�>��D=��ok���B�@�L쒆�qQM���Won���;���������/�Y���#p'""""""Of����*�M	��;�d"`��m����G�t�{�Û%���ؒ�:+��� R�צE���k�{���r6�9I���Gb����M7�N����d�B磂�[b4����u��x[&^[�۪}�Vm~c�#)���	(����1�G;�h̗���^����𶴽}k�^����W��o�<�~�ע<b��z��DDDD�͘�I�����z�U�5ZK�
�;K(y}~nT��	w�<;~ ~8tg��0Q4!-��)(�ոk�_YB�����j��Ǩ������鸯�k�ے���N�=�����a=pK�v���Rd�/6{����0�C
޻}�5g
XKd�4�/F�O����Rڟ��~�"�f��:4���(gҪ��º+����"��<$"""��2��.���_�&Fc���>�^�J�-1?�����>�7n�-v�`�_W�'sD�������-���p���"m~lA��@FʓkD��)���NdW��p�bW��`,}l*&�{��h�~�2ܛkJ�4|x��Y�H���N��9QXiz ����A�	0y�ْ
�#���J�BQ�L�\OO�ʥLl�%���)�(%3g�(�Ă3�uŇ��D�Uh�]g/(�ݜY}k�0�_D}o�����2�ʝ0�����з�,/���1[;$�~E��0|z�L�`�\7�)�>7��8���((�;RyJ�ݛ2�/� �)���t������v�r ��?����I���������r��L3٢��.��6	v=�p�c��D� �DC��ΗU��U����э7�iQ���
kM4m�8(�]��edl�bPZ���;��n_���t��Xi}1'3�m�w6��^s����!19��s��{;����	18�[o1�}�����9�~���Q��;���	�D���T�+j/p� )�Vul��ā7\�ʊ�r�QkYzi���.>t'K��@D�!"����ҥ5��z&ǚ	��q�8yu W��˥����S�ʥy�ٝ����8���QTU�V!A��OG̔&s�QϏ�϶����-��.֗��7�ݞ�r���#n"�����DDD��v���}J�6^pe �uǨ�u�������d�ӟ�lC�}1YZ�l�����?8A�O�B�Ij��k��(,�׻�7k>j'n�V=��w1y��G���{ǡwJl������������/�ɥ�����ם%p���܉7V�&X���N�aөsxGڎ�Z����t�?��+k��� Ӄ
b vwNܓ�v)vcw""""""j��OD�{��+����.�-�������"Yخ$J|r�8ć���>3�'�`���N}�2��\��jos_a���Z��sl�Ml?~9��׿�f����Z;ʨ���D��2�|iJ�X�=,��1p��G�6;�������ʝ&o�v�q����z���m=ڹ<���P�gRm8�g�sp-�g�5�����Y���^�}sVF�7�)" }G����LV�'xe�n����+~��3c$�����"�=���#�|�#���5�u�p'Gq����H
����|g�@��R�ڎ��#�F%����7��q[������q����u�L��)�!Mޞ��`�T^s����J�	��O���i�1���������P�Y,��]��ms�]xzDO|��(����}���v�Cv���냯fM��Ε�t�`U ɉ�}:�C�H�J,�]g/��T,$!v٢��>ߖiS	$�5Y�NfnS ���Gqum�'\,0}��;�6�(��E�P^[Kj�uxy�&|v�x����:9%�q���K�����z���l�-��ܙ�MD��!"""g�ˏ�O�S���I�����]���i����ߧw��@rD�\����A͕ѯ���k�2�=v��Z�ʁ��Iې.	Q7\?w�	��gOIG}C,�S[�6p�������d�]g�妫�Z*��v�� o��9>
�\ʫ)��%b��^����*���OD���9�'�-�����\�hdP�+����r1Ď�)/� ��~���"#>
�<8�6ַw4Q������׫,6l�O�g�=�7V�5�~=���6��}�k<Id�#��w��p�u��q,�Ħ�i-45WR��Xkߵ��5A~>M���X�oSW,>x
�b��N/=aE]�� 5����׸�x�ɀ{ZT��Yz��&v���צ�x���[S��J�b���܇G�D�����Yw��ծ�v�C�}��-Cq�?���	�w�L�k�����M��v�C��D�-�-�%�]O�i�<��*��d.��A_-_�S�ߘ�������()c~���۱`E)�vѦ��a� 8R��04����W&D����Sy�~���gyD�D˒2DDDDD^���d�5A+# �yߟ&�k��jR�6xjX��~�,1<���ؐ@��O4��d�a�˦\qWߎ��������^B�}��;G[ Z���L��!�4�}R��ԥv4�4�����+�m�ݤ�w3��� ?���--2-iZ�6�5������b��+�xUI����؉	5:|����Ǯ��~�@��-�F�f�`���ME���-"8��+���9���9�O8�:�g�?;o�"��"p��}��Ɔ,��juzy0��Z ӌ*�|�F5ь�����r2��Bsk��|]G��Q�x���__�� ����3QA��Jw��^��h�=}���-�
۲�����W��X�fO!���YIDDDDD�x���P���=�!�q�x���ޜ(I�V����$��7���r�]xn�ztO�F��(8���3�`�s���ef����1�}���#��Ǹ9��7���+�+K]oT�w�9�@\m���ZZJD�5wK�m�XS�B1w��,�9�u�xy�VPˑ�g�^p'"""""�S34# �"�noMmq����'cʜ�q�|�`h�D|v���پ��Y�c�����o���-���f1�b���g 1,|�\ȸ;���שCqo�Nv�Kd��c��^��+A�^���X�{oN�]�I��̷���&��[X�����T���-%"{���y�3��in���� ̛5�!����ۑWVe��Li�����]��Ϧ���}s�n��?�~v�Q�x�Sp�'K����=2��2e����(����W�n�d=QX�Ǥ������c�1k~q��?r�"ܕ����m#p�����\i���/�8��)�����o�쉥@�����~��75�"}�tpYk&����V~��Ոr+�]�����OS�zT�7�N_۠���ז���X�9a��`,|h2�D[._��d.>ݞ	�;3܉�\�#v"DD�@<��fi�!KiM�Z��'��������ixn�:�o�Q�Ѵ�����;t�e�2���kJ4���i��z����K���ʧ����b��p7b ����`t���O,��g���	M��m*��Kգ̕�X����`�0�T`���|������H8UX����&oOă_�3�Z�p�V�VX��D�5Y�oAE��Vq�:��jM��w��������lÈ;Ybl�Ok�k�~�ֳ=��5��V�w��I�����rYw0�}2ޞ1Rn��H"(��+�Lvs^Y�]n���`�h�����J�]�|�Z䗻G���ɱ���q��u�����յ���Ȱ�c����D���ʦ�U�3�5����گ������WY���+)#�9W`2�> 5#ғ��r�gY��XSRfDz">�{�\z���������8��R2���DDDDDDt���AQ�����[L���\�*�>y�5ؒ�W�	�+S�`z�t�����o��#g,�O���vZG��_j�C_ø������˲��|{���$��0����b �96���W���	��ZG5=�Thg����|������~�L�h��o=}w��|nd/��M$\ai��!]��*_&��<=wv�͇�HKA�m�DDDDD^������/۳��u����5Pm,-*L.13o�	��b�\缥�����C�ə���;���e��x)V>s�D�9��D����1k`���mXu�L�&uߜ���N�ЬvA�c~���x/܎�i��Y�2���ƾ����l��������6����-:t�Mbr op��ҭ-�;p
�`�������~�������{;��G,��n¼}'�D*��Q%7�U�Tޔ�2��/"r���j\R��C�W�m���I�G�3z�Ǵm���L��a?N;1���u����������;��8Qe��K����v7�m�(�탓p0�o�ً%��,�l%>��S�ܨ>rG��/�e�Tr{� zX4�W�A����`im����5U�<4:�'��m��r:�2�K���c9���j�>�O"��9Sly;���=�1�k��n/�[p�X��n�Y��&���%�Āɳ6����>��<�V���NDDD�h�O��Z��^N�2^�����3IkeV��q�S��i�P��J����"��!_��A�
���2���mrƴ#�EQff֠.X"�n;�G�:�)�h�9�kL랎a�+�c��=���m~�������ݣ��LHg����+��I�W4Vݓ��l������}: =6���U���~�d|���̱s���5Y6$�W��:۳�/��o�j�;��K��zSw�����8UT�,ij*@�����)�6�b_���[��;0w�����F�Ӻ��-�ۢO�Oq�f��e?ٖi����̟��71�b�9� ^�_��2+ʒ������I+��ӧ�`,)CDDD��ϓ�J+�`�,��J���~H��\
��tU�!���~�AUh�aQP�B�o�AÀ��bĝ���3�������܇'[Uw��D0|D�$y���'s����>����-f��KJD(�$Da@Z��G����֦,�wO|��lV�5v���;>Z�y�r���Y�`�#C�ɓ�]{<۳/�@n�Y��S[ISnJOD���p�y��d���8GnG�y�}D���h���pw�ע�Dm�^�=�2�銲�:d�I��EWk���-�K��ڽ��������I��W�Qe���5h!g�7E�ޘv����l����Ԣ���dY2���m���\i%��|���<��hxL����2�9MDDD���됴���i�B/�T��ґ�^ ]���hI���p�4c���Rz*�z��Tj�.״���*�t��\"��n�J��E»Z����U@SV
M�ih�ש��Am�C���6�Pg]�I"r�~�;q/~�A�	�L���N��IA���8[R!�=.����`��!�䇎�"�lRWI9��j&�f�3>\��fMtZ�{c����G�<]QPQ--oi�W��Q�
���#���V!Ah�¶�s��W+���o''2W�9���չ�J���_�u&^ú9�v�ڳ�¤�cQ����=�p#�����I����6	��xY��_z^_�����6hk������M�-ܗ9�'�]+���)�P=�������s
� Q�ݛ��DD�Q3�V�Y��Q(�F��C@�W]��ue�d_?�KOW_��c[P���(�aO#��	��'[#2( ���?Z�ʈf��n(�s6��K�69|Qo:��i�/�܇&��(O}R�Dv�h,[�RC���$r<s�۷����"��[Z%gA�0�[C�����T�9������=�7��DVyc�윇�Z�E�L���|�U[�ҭ>��y"��z��؍��%4ٸ�TwS��b�&�l9䉇v*�J����ُVC��-Ý���Hy�
(�������l܉H�ƪ]���ّ��DP����z��"��L|o!��5A�(�VG.\�-,F~y�Z������z9��Ti���H����o��G'�Gs��-���9~�pz%��Z[C��Zݍn;�\��/��簆��m}��~�x3*j��^Y�z-��1����SRfk�y<5w������VW�}�ۿ���3�ӭۉD��7�Y��JDDD�r�e ��]��d�\��t�\����ۈ,�'�Y%�w6l��y�⁛10����b߹���p�B�E�q;J�#��U���"��쀀��3�������7�	�7�o�i���}��㐦���ǽ;���1�R->UM��d|�\L��=�Hˡk|4�!��͢-ؖ}��}J��S��x��!�{�z�%eD�ۿ�ڍ�wi��כ���;e0>)�dBA�����(8@����z�D�B��`�[k�ȧ��~�0��O�}�w}�o)"�|�����iC�����[�r1��&3LBŀ;9�,7p�h_`����r0�͹xad/�ۯ���*z��3��-�y�"��x1Fuh��삑�S�M��o�9��m���������7&�"h�ΆXs�l���/¸�������#1<��`�xQ>��͇�ƚ�V5��$*#���;ڒ7��*)�5��/XDDD�(fGAD�@�?�5G��%�1rD����L�,*�g��CTP <ي#g��W�\�ЮN�ǳ��aÉsx��+��D#ZѠW�og[Q��I	D����7��k���Hd�/��9
*j�������}xaTo�ݧ�٬��ϡ�� ��V���MV�ANi�\:��竬3$��V=#O�z���	vZt�ܘ92��������d5�?�v}S�0�K��n��	��.�/���)Ė�yXt(��l/Y%��ܽ'��P6��d��<�>��<��2�-�eT����ީ/}���R��^WÝ����(��w�������O�b�?�⃻G{d�QB淋7��]�)�n�I��)�{3GbP�Dx���������92�@f��Г��i���p�B4R����׆(7�=�43[�����p�z�;�\�'{��M�v�qy>�k���9��XYc���=j���[������N���0OF��ߒ�ُa�l��u%e�F��#"""�Q��z%���~3�+���9��Q����Sbf��<<������8S\.-����M�����M�`P��y�x��p<�qHӌ��O�<r�L�6�W��z���N��~"�oiM�<�{�3�+"U��g?��Aw�+)�R��o$"""�Q]�xC�����
��r���[�C��8(�������ri����L�|û��a��,�:u&tN�R���פ����{Ѡo����{s
��uS�Z��0n��M��@�
/�A�G�9�.2ܽiO�~G<DDDD�Ph�]���ND�Eۚ��p�p_��zl�&�+���q?��f�s�u:���r���R�ꐌ�M�n�1P
����)�^�E��o�'���iDc�}�
�3����χ�d����J���L���5�.�!�w""""%Rj�6�^4�R�'�V�'���O���='���xtH7���]�@�7{����;�[Z	�Y},k��`j��rI��&�4�Ѵ�e۱�}����]�y���	�M�GuHA��8��v�w��uf�WD�]���p7h4�������3(4��j9"R7(;TYW�W��˟�l@g<:��.��*���Cr阋U5P2�q/�J����'��Ĉ�IP����!�O�u{��\��_���=~�<�_����m��������TyqvWYM�tz�E��+��2�[�]�94KD���LD�%~Y)p�at�x5��gB���J"ʳ��n/��a�tl���wƨ���uA����x��u�fAgp���vG�"�]L)����O����Qa.y=G/��ZL�6�{q��y���ErY�IMg��J���7uÿ��)_tp ���;�=��%�˫@�P�,�"ҿ��o���n3J�u� """R �e1�{"�qü QjfYf�<�3�;�bb�6�6ѩ%g�����9�:z�d)>��Z����V�'Q�}b�4��HE��hh���� ��#g0o�q�+��r�oy�O��?on������mԡ�� e�	�3�{��A�ࣕ�S�1�+I��ΰ�|U����b�l܀�܉���I�}�UL�v;<Ɋ�N�j���c�$���c1 -N�����p�h�?�'2ֳ/�#�|�\#|�|��������ʓ(�#7�ţj<�&D�kb���mk��z8�R�i9�;~N.��m;�o�2o�I�q�@���Z�|`<F��@n�Jʑ�'�vǽ�:"����x��|*g�UD�]���XR��0����Z��9:D
���L"�]k�t�V�FRDR"��`pdP }��V�7Ie�uh0PTY��U8_^��2�^8�&;��ip�X����N��w�� �߾�u�F5�:����t������b���"βy{�>�|s��߿o������k��Q2Q"��a�1�[[y�nal#�����ٳ�qu��J�]�g)7�Rw�D�y�="�fQ����A	"�Q���R�z�<��@��ܹ�C������l8��vF��������cS1�?�Y������uJ����.���y�l;i�|���ݮ�k/_�n/,-CDDD䮔Z]�m'S*���""��kq�v�Lst9����l'޻c���u����ǧa���SRr=q��}�;��H�i=#�"���wic�7��p�^�����%1E�Hy����,���,'�|��(n��c:�6{�6ѡX���x�۵X}�,�婥�Xz"���	��������[��A�J9��.W��ADDDD�I�Gj,)C�DJ��9Q��'d��}���[����@��Y�sgM����K�z}�疒��=�1�O�������=�Wљ  ��IDAT�"RU���w�GZ������^����GD�LJ\���5�ި8hFt=~-�Dm�Ǿ^�//�7G���^���x<���<�r<QWr�4��3}RZ9l�j>;�m�!uh�{��DDDD䶔���Y�x%�~�1Ý�pf9�G��O˶a���Vݿ[b4V<u+�g���-ބ��r�}��C0�k*�uk���[�%d���Z+2��l���Ւ2���Y�DDD�L
=�72�K�h*��Bt#��go7��vR#�����3.�5FtH��ێ�ߛ�TQ�:�l��ɱۡ5�tJA���?'������R����o�;��9���NDDDD��_D�sM,��DM`���h�<��l��F���v��1�����uƪ�g����X{"��GMh$7>�!#:$#�B�|G���1w�IUՂ�A5)��K�~{����W�^��V��!"���m������W���˚,i��e�;�e?m;y$O�Z��� �˟��:����ԬǊ(c;������Xx �8�=9�V	a��.��0�M�ń���W�5��G�����-�9��0?Ղ��߾ՙAw�j�*��������؋H����N���Ȝ�I7A�_�[�3��x���6�f�D���=��Lq�efc݉s�t*�u��DA~>rY�^ɱ�)]�f��!.y-��h�a|�������RTF�g�倻Z���w#��DDD�PJ������gB��w"Y�p�md^ˮ�X���J���#��k�|ZG���!]�Id��9[�-Y�;�@�Η)+�Z�^�S\:��@�Hd�E#=6\�͕��l>���O�N�!Y�#�}�]��On��9|��JI�-����ܙ2���a&�5J�T1Ý�	ܷ�i��n.:���E���1r涽��{�'OW\(���sE8r����8*]����p�������F�"5"�ҥ4������B�̒k��:�r=�hg|xE�\g4R������LD���D�l
��ss�~���%����p�ѻ��m�� _-}}�� ��ǾZ���2���Ҹ��

@Ym�<?��E�Z��KY���BYM�*kp4��.�Da�U���gG�Dy��`R�� ��=WV���er J���=?��5׉�_\U�?/�n�q�S�1�����Β�!^�[�]]>�zmծ2]��iQ�7�W����n���)�N�5������ZD�����"g��D��z�^�jp �O�b��S��u\yF���v���1�_��=������j�Hq�A����o���^�/�נ����ٻ�6�����v���qb'q�ك�f()�P�@Kݔ���JiKK�e�2 !{�A�r�#���%}�_bǲ�%[�u��W�w�i8>�=�����b���M�Ҷ�������/���[��יo�b��!5*���@#}�c�&���'�|�1/��@_D�KSL�?�<(P���s�݃g���L���H�e!>XU��7nvg��W�����u���{�l���^���"���-��c����c���9��[����`��lQ%>:|��9�23:�����+�&oN!>=v����s@�?�=5�j�8Q���ힳ�l��Ru�����)åp���~�j��1�]%l{��S�����oMJ��T��+:�o5��$�Z�^!�8�#ZG,7��|�t�g�1�c�a4��`7�d��[q����5V���o���C�{�1ŉ����.m���J]#>;�%�G�KA�Ma�u!u�+��{ݠ�DDDD�$Ӕ�C�ɜ��C���M�S\
�M]<9,&�[2�MK��V��Ƴ�p����+M?�7?�d;6���~��m��/r{�}�}"�����M��J���~8{4�8p�5�+������%��Ȝ�N�^��^;��q�Ww�ڝ=��Y�˖YR�^�s���'�����ըo���K��p�:�㖓{�{��{UK���L�4p��&�v�z���Rs�������م!���!1,�{��y��Ӎ���.��Vn�{OۼMWۼػ�� ߝ'?��������ӕ;m.W�����9�\
�ۛ����7���Ϯ<Oџ��;9�R���Kwl��ǜg?��qC�Y��r���fl:{���ºӹR�N�%B����U��������h���JD��{�D��ۛ��E$;��O7�����ݙG��'��ݱ]��b.�>����Y�M��!���=s�,�U�bs�E��*�oK�]U��we�Ļ'��{N"�����������n2�cfJ<���O�f�t�֓O*�D�(<�HBlK>�:>������Q�a�;P�*�K.U�I�����ؕU`�J$�'��"w��-e�z�*oy�DDD�����H�O�3q���g�T�9i`�S�Mc���E�;���0 �Q���4���J_S��*��Ŭ�xl;�g��ק`^���D��k���O<ޓ7����}`�秴��C���� �����v@Q<��!��eu{q���Sٖ�6�^���p"@���&�[oo�Z�J��㋦H'I:zu�Y��5Bס�T����aV��ќ�.��+)�f�N�Pzh�-�+kNfKSjtn���C%�D����Bl����s�8YX�]�~��{렩,=""""�`�y����P�-����%#���A���}-��F"5:�+:]��͋������e5�]�@��j���.��N�Kӳ[�"�W�������N����$����ž�B��*;{:�"��٫�}r���u�d�����r�᫽p�3[�e������r�,�;N�=��-�Zs�*l����G�E"9"��5p�B��R��#
총+��c_��o��m�6���1Cpèd���ۉ�u1�������n����t7t���2<�#"""y��^���"���a��*ܗ�[���8�_-�dU�,O}zc灻=��p?�a���c�;�{�p��=��ok����2f����v�������u��=�{;�Ӳ�X��*��%
'O)�7�fu{���f�.����HfI@v�i�B���Z�����m���Ӊ����풘~��.LM�������'�pR*d[���z|}�D:��<�/e�N)t���<�'��)��?mp���Rƫ^+y.n���e�N�«�S�MUv?l�!B��y������h������v�^��z���P�-m�*��m�ƈ�t�R��GZ-�[:��s���
w{���^�~jbb��H��v�j��D hK~���}���l0���N�7�����A�'���L����Vh}!'"|�s�P��P?L+�{0}p�c#\��x���x�����e�W��19��1)���U	.��^U�΀�����J��7D$k
ׂh[��l5���Nj�;��*p���pdw���n��UBAu�K�ᨏ���b��{jT�`���������V���x�ޠ��}ǀ'aݙܶAa�}��"mοXS��y�u����W)|�V��-�Kޣ��P��9۪��r�I�T�	Ǩ����H�k�}=g\�� ]�58WZ���)���WV�SWt%t��
w""""y���Ox%�	��q7������/\�猳Z.����������I*�E���D�ltp���r������� T]���[Oc�����k�X� x�P�l�C]�����4����'D�{���W������U����k��:����Zi�O�-8|�D�ڋ�3�}�!>41A~�	DT�?B�}.O~b�5���F_��� 4R���fi�Қ�f��7����<����?7"���Uu(����C�n���^��x�,yn���e2�n������A���c�0.!�j��s�w1(��*��c��:i+cg��1���k��nI"l<�gu���QN���8Â��3��mڍ�l�}Զ{���]���o��m���(�� �J�Ǯ����d�A�\�x���
��ZǹG��v"t�2(�j�㵀�.�R�~�\� \L��?I*ޣ��x�J�W�5�ۮ�!�"t�S�>O��?n�,t�������H��[�,�g�oqϟ\�
������L���B��;��Kߋj��Ee7��6C�¤��g�\�r���pLO���Q��-�j�6�s���j�z�Q��ePn���T��
QWצ��K^j���̖�x��������F�[�8�G�e���";���U��p�ń28��B9"*�U� ���@��ZD򡸶N�y�������<�@DDD�%�
w�/!��+��!��I��տ]R'Z�ڝUh�׏�0p�WU��y���Y/�8Wt�9nv�߽c���κ�|�D���=�B<�7���C�G"%2�b�g����2�Z��Amuz�����v���^���D�;?ר�_�:2D�_u�{U��˯�[^+�#lEE��6?�����f��!��H�n���N���K��L�\���x=i_v!6f�t����@���
�e��h',=��W���`��tv,>�D���������-��h�肉N�����J;�u�z�OP(C������)`�:��;Q��8t���2WTy:����dG!׊:w�<�W��Sw��&���B��X8| �*�^������&����@tL� F�������,����]._@��@��#�ƙWn�Z��%<��a�{=�Z���J������U'�����0!ѲE�7�uj��v��u'���99�J�6��R+���cJ�
_Q'�����%�������
܉���d��A����h}�I���,��NF�%M�X�>/�<����7����91����p�
���N�Nh��U<�܊Z�ybP@[D����6���D������J�/�߮ه5߽�b�J�\�/޻J]������ ��Mbs~Vy�B��Y�1y �D�-��Lگ<������v&W
ܕJ�W�<�@DDD�%Ӗ2l�C$?M�+3E����n�G��q5p/�m�#�lC�V��F��]�����X�zY4|��e;�_���۫�S�.�I�����i9�s��z��L�=�EX&���t��ű�2��`5R� �#�N�����뼒.=uS=�1�4 "o����kY�>t�w������<�l�����	�Ad��' �5kh�|�_�9-9��~����w[V���h�w?܌A�A�`;�}l�$|v�ݶ-v9خ�?mB�|l.���^}s���j��xD2�=p����<Fi�k'=����W�_�����.�e9�o;p����� \��OB����jOv�����1Cpl�/��*w�Ϩf�N�},Cw5������+�Gb��y���u'����kIz2�A���<��}J�/��"H������ȭ�Q���'ǫ{N���:FԢ�v�yZ6���.����ÙV��I��j�E�[-����ؐ@V[��"_0�˓t���,�_g�I���ز#3��k5_�R��o�ĭom��� �A>�a��AY��s��~lQ)��[������	o��	�cdK"/����5��2KZwo�p���IDN��O"r�l{�s{�I�^�\����^���# �90�[���.1�j��^oc5��W+�}�P�.o'VL��l�o��������]�j���u��g;��]m������C�5;_�,N������03%�;\���_ۭ�ߛ]h3p�U�p��{�_U+Uw�T���%8~��f/��
��{��~<w���]���Z�y� �W���@��i^j"�>��F�7�����E����<�������П7��)�ӸV��;� �5���ѳ}nJ<r3�2�./�ך�;5n3)�7�8+]��w�R̺R]��7��իQq�(�laK"/��L���C���NDDD$Wr��M]h@=������[n]��BQz`�l������}������ןε{?��
��%J�g]��~��j��V���Od�Q���QA�xh�(�s�a8K�Cyi�<�o�;� ��9ew�����SFH'*lI���#_5��v�'�|4j<2w\!�������'��o��ۂ�ڴ���Ү����I��xj�!�s�l��E��G;�����w8�?}󬶰��K}7<�tW�5*�0�l�@0�vAJ��e����I��*i��߉�C*�M��n���DA��Ź��ޢ�7�/�������8���*-y$ADDD�$�@�^ A}�Di-�IC����e�����sǏBa�|�E�tv�0�0t^-�4�F.G!&�J
�<���e7m�P�n�j��̾�=�Š�"t��J�yi	������{�7Z��Ū��34�6���h��������+���o���6�Ta���k�|A�a�=⽱�v��ٽ��[����U��zwM����[{��i�}��C�-���w?܂Rc�"Z�,�j5p\~�����7��2�=���o �������!"""�%��&�p�=���>�-|x� ��E���K�ՉCQd
��,9���9�{f���H~1&&�X-[62�*p���������͇�ǥS����+?�5O�?w���o?.��!og��x >|o����#�x���v�7�ȝ��� ���3���[��/�Os�������6���)#\�omc3�`6�ͅ�ĉ{�g�1>��f�GDDޡ��;�Sȴ>������7ᥣyH����ϔՁ�]D/�l����I����\���}шAЪTh6\{�UO��7ڜ���kbR�����f��+{NY��qE}���L�Tm^��|{���/vagV>����꼭OfI%�X���������Шw%p�������x��t$G��������Xs2�[<#�":���'��5�PP���N����q�5�������""��x�/�ȵ���a�'j6q��D�&���um?�7�-)�.�|��7���Z��⣱��z���'<YPn���w��N�T����Q�k-��UJ�n��F��}ĦY��5�ȯ�s��ݑ��r��t����ُ���� iP�����un�d^����?�{w}��b�Tq���۱�g�1|z��ż�f��WGb���oƘ�ȶyUW��T�:o�)#O��'Fa~Z�y= �$��/�W�@N1֝�E����U�\�g�+�8=F�	{.`�L�;7p,yo�p���ID�d2ɱ3�%��Ű�;�W�XY+M]%*�Ws�
Y�ή�*��&g�˛�N���]��br��'�k��U���u�~G�K��;_,���"���w�qi"""rM%"""������
w���W3A�uF��������h�5/-	iQ���AnE֜�����m�~vj"��C�~ί����#��J<4{,�uM�lhDFQΗT��K�����<�<�v�A�QoJ
�s��Ǭ!	V��1�3��w׵���[SGa�蔶�[���w�߮]��V�ǗNo���='��g�@�J
�M&��sr�DϨa�NDDDD�g`x0�~9bC��f~Z>~�,}�3��;v��U����lh�磶xZ����3��]�T2q'"""�T2.�0�����|�¶�]T�����ffJ<R���n;1)?�7Oo<�p���O�+;��x����w#w��m��y
nx����*�T�b4�`��� """"�w݈dL��sVi%~�j���R��S7���G�-�ެ�x~��7饟mE�b�ﮟ��/~&�lU�Σ{�-e������,�<
�<|����Oq��DDDDD=��)�?g�^��4�L���ݸk��i.k�烹C���d����Nm�5)�?|6��a�;uF��2DDDD�N��iQ��%�1����I��G�@DDDD�n��}f�� �E5u?7�[p0��b0ՙC��wS�+K�#4*����K����\hU�����{���Pt+��B�{u(q�D��7�be-
����X�NDDD����~?st|$�����zBBX|4�D��Jju?'G��}߱Z��}'q�4�b"�b�p�+�u�8�1}p<��I��@-�Q�kĩ�r�-¶̋ؗ]�&����DDDDO��ퟹ�F""""�� ��t������B�}����1cH�^l���M�/>�bqV�;G�O��&`ńaX4"����a��׌�xi��6�[��t>��,6g�JW%��֖2 """"%�M��;��KYDDDDD=�`��g��ҫ�=�eH���h�?�~?^�{��stp ~8o��m����a�1�N���@��_��i�i*�k�w��
]#��DD��ǜ�\`RkP8j>4�uP7Ԛ��J�k�0���ڷ�yk�)Q�����159Dr���w�ŝGAD�GQM�ռ���[�u�E_�VM5LXs�<�a|R�4oҠXP�D��G�ǃ3���=��~xl��q_�{�tUM�m�-e�[6EDDD�ϙ�;��������P77Bi����&(��al1�k�R��Eo��7���%�
�Wv���+�?
%*u��&�F��&���m��*-��2��ܤ����:T~��J��l.������z�y����U�H�o�
���v�O��S[u,�3���E�������h�q�Rƒx;n��?.�.���U?�=�O���ߏ����yDOa�;�����E�_�_����k��-��MB�|Шoqz�1q�(�5"��Υ�3�̙��E��p&})1,Ȣ:�����/�=���f�i�9��@�>jU��"L_}���������a��|��{G�⽙(y��b~Z<AD��~��6>��`#rʫ{�q9h*�U�����ȫ.�)P��Wqv��5�
���#�10"��}"���A���V�pnV�DM�KU5*%���N�?��g�1����|Q��Yc� C1�ُ]~���m�z�j���MGBX0t�z��h�^Lz��5HӅ�J�.(�[���9�Kr�%���F�;���j�C�����3���%�k�a�%ѻ��i���1!2��� U[�)ټo�j��l�*�U���x��п|�k~x�U<c�ˮ5�b"����fʠX���7���ᡳ=�x܉���<ؤ(�H�!C��r8�����Ve�/9�Wcu��Q+��TJ��j�r0b뚭���7�H��:���&��}�y�ilF�� ���c�[[��Pk^M^� >�V��
dT�#%G�ⅻcx\d���h�q�u�p<�����^�~F�	eu��D�>
wLHë{N���[T��0����cΐ�f�������I���د�:���MЬ�$�u����3#\�]z��]���.nu�K��ŕ���ɂ�-�(=���f���:���Uxv���ŵ�������GVؼm�y�����e1Ϫ�L��#y��p:�ғ;܇��wg����tx|��DO��y-�&D�7_���3�ї���DDDD�(�W�I���uP'���Px����Ư�~� �a�'��h��*���.��M���7o�y�`qɱ=���c˦#5&?�h��?��(�:Z�
��y��X��Wȫ���1x��k �����s.=�E#I�A	�;�a�6�\�,����C1:1
K��tMWO�|~<�*�,U�����`�{�a����;b���Ҳ�6A}�g�KDDD��������e�6�X�7V#��q��Cf��ڽ�ּ/־o�ҋ�v��c�\�=%r!Z%���w�:��U�p'"�&��^"����	�K<����`�����w=Ŏ����ˣ���7�aRr�����ΗTJ�Y��,�R(�b2�RU=>>rwNL�n?,:�{�=x?�;��2�ǳ��-�
��H5� /��_�ۼ]��X\
��tƈ˩C�{�'E��[�җ۵�?�l>��o_�6���MEI��-��6Y����w�	y
����mR?�����c�B���_�������}G���Rp�5�ud���G1<6U�� q������1�hq�͉� 7�ӓ�޽�p��{$t�w�R	""""��xu1��;���F����g*Ez��o{�S����'o�gb/x�]\���#��v�OHm���X0��6/�t-�awܕ������O��pW�����F�75c@p��/��ƥ��fLR��:>;���,����jqn{/�8EK""""O��l�4	A�Z��Lg��rH��C�64�H��>�bVL�_��J���=Kp�k,z���DDDD$[��q�0#b��1ĕ��*�!�B������[fK�a\�YZ�/Of��Q�m.ߜ���eN�O��-}/.o��a��{ǋÃq��X�5��t*[��}�&Ł�+��K���"*���dDDDD�Ι�������:lo�p� ���xt���������{�����
�� m�+
@�2!�I��r8�N�N.��㎧I���-u�%��7�#�l�����\z?�3����%#O�Ԟ��/!<H
����ɖ}6ϗT�\�[�N��NF���j��;�H�;y�;'�O�MD���18[\�7��t���G
V��a�z�!����J-�m@���c@��>�҄����B��{���}	��}����74�b���r�t��g���i7���8�C�'�v�-L������FX,�u.��jD��Xߝ9�b��_���	""""��a1���-s��<y�,��.ę�r��������8h4�0��0Z�拽;������q��U�NջV�����-:�9�� �������V�{UCL&8�q���j��� �_�������oBD0f�%��$1Hj{����\ۃ�
���U�5jxy6�W�3���q�b�k#�*�ϊ�X��'n�������O���ǰ�T�������S�V��oh]���k�s�u���03%;���r��]�LQq���x`ڎ���S�q�̱6o��L���'|�~T��|��h�x<�AÈ����£�H�����h���l?��u��S�`�z"""�O}��4�%��
*�=��Ե
�Y)�V��_4	�^�<p2 �b��E�����p�Ri����Yv�MM�ElH��e�_3
ϙH�k�ADDDD���<<k,���/������(��
w��DDDD2c4)����	�Kh�h@�b4�^�.����l����Ha��̋�sǤ�m�{N�����w���X6v(��FZ��LA����5y��e���O�M��V� ��jз�d��_��\T54����:���k*h�*i<���0j=�D����������y���<[j)�߅�������5����:B#""""�5�4R��I��V*`p��P!�R��2��_��R1:�j������A�m�[4�a�.~�����NF�}j�~��o�g�W^��X��~t"�,��J�Bvi��:�}��i�ж��-���Y�;mdۼoO�o=�'N��ڦf�ϻ�]9�;7��/b�w����Dx��U5���9l���×��U^i��b�904bqcz*��P?��uz=��bwNvg_�~�h.~8cJ�='dx�Q�����)�����l?�������;�L5=�ʱJ�(�`����v�!�=O�UwǴ*~9b��ŕ��'ې�߻I��&&Fcᰁ�p6��zfI@|��.�jJ����x"��V������*���[�_?(_9g����R���l�y{-6��A����&�L�`�8��� �5�؝�9`7=RPdu��S�))ï�mŗg�Y�l�xi9�U��ɉ3R��7Ǥ�fbH���խmj�Km��.����""���M�7��߹f�Ӆ.��V��񸇈��ȫ5+|�ijuS����o#�Z�0���p���H
��ϫ���o��Z[�+��-�]��ݷ�+��h6f��VF�lo=wo�;����XPS~%��c��K����{����m�s��v2�-���jl9�'���O�"*������gJ:������[#!�D����v![��`������-xb�N<�}�����7������)|g�8<�t���>���;Ϳ�m��r>'����y���DD�n�y?q��xqE��7�>g��-e�����&"�4zx^����I
��(r�X�Z�8،����'}���|��(��:����,{����E: c�"�tD2V�ʶZ���R�[Q��[�RծU�{��M���}�W�]��QatM��ۈ��&$EKml���Zlo����|��}�c>n���F�����]�"�G���럞8��g2q��
rV�k��7?���|��W�Di��ؖ��O�u+ң��+(��'Ϳ���p�R�l�, ""�}�Q�F��d���X�a��YR�T����DDDD�M<��]����ag\9F2���"����MR�{��j�{���9��5{���6[E�-�Č~�������N�W�s,��#������.W����(�#C U�ט�w{�g���>Ɵo��%c�`Lb4��� ��RO�ិ��j���3}��;��'o�����sێ���|���xa	^�w+Oe�����]Q�E���̲�{�����7���;05���v��u�������{ɭ�����%"�l�~>�a�x�[ǥu/p7�L��#"""�����t��E�
8��� ������ͧ[��mVY5F��]i�QGD+�n=�vÌ�q��iT� ,|��Wպ�|_�~���T74��Ŕ=�R�V�:�|i%~�fw���n>��)�������8UX"wx|�6|y&���u�:�UJf'��ä
���i@���F��p�R6eeccf�T)o�8����p���������g��.^�BD��KO����V��]�#w��M%"""�+�絔�I�#V�h�?h����zl��s���Z|�V��x@�����g]��YTٿ������O�\( ��H����r�/��s��>�I��	���u�h�,����B1!>V��^߬�+��o;���N�eC#n{�3���R��.2�@DD�aI�`x�`_-&&�`o����4����H��j?x��
���1F9�����y�SťRE�#Z�
#c`\\��EcHD��!<ѫc���˂}}�;n�����'E���)R�~�'_H��m9RP�W̏�����O���o#��I�ǘ���S4[�	��J@DD�!N��MM���2(���]a�+܉���dJ����������a`��z��U�v*�ADd��˫D�|�%�Y�		��h�|���Tw��S�Js������vL�Хu����;nş6���6m�y�ط����^��G����'=�D�c|B�y�5�^⤐=����?m��܈��s����ڞ{�	��t?�p'"�
��$"7���맀��:�� `#�G�>��{��T����b����k���q�1H	�\����iJ�u6��q��]�[���f�����u�j��������kg����͏͟)��͓ەN�b�
���ͤA1  -�kc��V������Hf}����LQ!.�]Bj��bWRi��Q���!"G��(}MT�������;������u�1�N[��u�<>o����]q}z�4�C""�5<ڽ�n����`�������!"""��P��܏�_Dsc1b�41@c���/�X�ND^ൃG�N;�����u�c��U��9���O����U�<sέ�+�։�d')<t�}Zd�?�k�]�M%"""�!�I�0�^\�B%��q��� "��D�nˊ��H
q��ݔ����@��Y-{�ȉ�ܙ6�NR�V��c�.�l)CDDD$/uF�>�;"6�.!H�rx;G=ܛ���$��-��gJ�l.�o�yLq��ui)x��1�e[�r�b4B��^[��`w""�	�〩�B�|\�[��P��o����J�׈R�F����f�H��ID����ٜ��I=��S�l������+�R��H~�4j�e�.|�I��d�' ���}��j��x]�+܉���~!������{��|JR��e;���&p�&��HvD�r��+��^��]�����A�7�Bjt<LM9o㰇���DԿ+,�9r��@�F�D�W�FcK�ղ�Ŷ[��4O���Q�3""o'���|�&oP����}��]�Tz�'``5?�Ɂ��]
��ЛLhlQ�� ��YP��i�]c�M-}7i�Veq��Va��Z� ��6������5H���J�[ՍMȫ���lB|L�>�����E�V�N��/��lɎ�,�
�5]ܽ)�V�z6"""���F1�ߏ1\�<C}��碰󕈨�ʭ��[==0,��?52�f��QZ��`0�~3xlND乪tM��J�t.���ZʘX�NDDDDDD=�����|�B������6��57_n���FV��NAu(�ա������.p'"����C�*���� t�!�v�������*��&#��H^.U1p�ʪ�r7��+��Z.oz�DDD$s�>&̉7b_�:������:�&j(�- "�D�mK|HP�<~T@��ee:]���i�^K""�\��f�mOs�bI���u�
6�#"�x�%9��u�ϨQ���jT�`R��(3/k��.,D�.P�b���s�R�X�6
!�>��V��Q#�G_�>j���+�ֻ>A>Z���w��-]����!�G���$=1��Gv��H����'"r���z�����z���r��k������7m{����ܙA�'	(����=�MA�MX"O�~7m`�	���<]jiB`�D�����9��Cp����O#�3p'���^K�J�+�`?p7{��K_<&u�٢
T74!���J�/�q>�K�U_^��w>���`K""��^�Dm��EīK`*]��C�:x*b���}���}���DD�QI��
����.8
�}Pm�
w""�i1����Q)�V�
�P\S����J����<�ˈ�r�� vkRT��egc�f"����V�;��#��	�i� "�Ꚛm���]�TviYOa�ND$O��xu��剬.�׫z��L&���;yn�P0q'j�tbk�l��>�9q0c�ЗL�\����KS���k��B��Z�8
Ճ}z�k䠩DD�������ͳ�Q�}v�\���u�"ty6��!j�P8TD����/��l(F�NG��/�Bg�[���p'���^���K�������_{���DD����kN^��q��6{�p�����o���-�u
w""��`!QE"	�f�,3���0%�/.u�G�a�;�_�Z�4�[z��+쏑��R��;�ze����uw��+�Jo	��(CD$<0#j�ʞ�J�D@�IBXD��Ġ/�:���e�;�_~����t��^y�ʆ�˂�"pgK""�:|���05�o[V�&Q��թ�Z�����9�o(���������Ug��Z�A����x�FG!Q={����E����D$?�>�O*����ۮp��h�d��AS����Ok�b����-�ڰ��'������hT�zitx""�̈�t�r���I:�pW�4�t�!��ӢQo@s��z4��6v�%D�����
z��M�÷W�\$�T��p�j���N�c�њ
�(��ټ�J�@��/��\:���A�������V���F��Uc�Z�Є���8x~D�(��vyo�*l���}�`䕋DDr��B֟�������X��G3���
�E���BD���"Gz#pg�O2�٠���������w��2�p��X<8{��e�&=*u��T^�CAu
�j����6��)���{�X�{u�q�r�v���ń�h|������GR��^�����`��_��=oeq��/��	���Cay%~���8-2�N6�������I'	�q��/o;�U�3�i%2��9����W�\Y�����C��a��gED�~�j;f�����g�J���sw\��:h������2�gS�����AS�]8?l!cr0�޼�������S|X����%�|:�n��ґ��.9��\����\>��oN�����X.*�۳���'F#2�r��ؤG���z
��<�55#�����a�����1o� �����L^�^�]��I���v;����������p'"�?qU�S��˦��zn��+����p^U��We{��""Y�QG;i���i�)OZT��}gL��ٗu	�2r��l�J+�~qz��<ѲfBR��ީ��z�AV����{�
u]s��5�_��fǁ���2�샍xz��ǱE������oDRx�˪@�͆D���	6������Uy'�Jl.����pDD���ۏ`nj�yJDs4�Y��m�k�p���]�
w""�m5�H&��i4j!7"wQ)��� �ߛb�,���3F����`�˖�Lq*pf��WmY!��Jѷ=����M���T�����wr^��#�p2�?[<ғ��0��̋����6J+��3$2��#E=�/,�;h�Ԥx����DD��8���6`�OoGT�?�1�ѽ�C�� wi�p��Q����Cw""�fR�����, yp�/�Z�� {�&�������q�뫥�S]�t�`�ˮ��߯�m5_��	�^�����[�tl���X�klw� X�7u��E���o����'���m�G�-ەy+�� YK	GT` J��L�/�=F��c��γ9_�OJ�C_0�Q�QR�Ê׾Ě�o�������W�u���R�[^+�l�z�<0�H��\��S;c2�e����_}���]Xv�������0>)ߟ5N�@���H�*,�����~�\��>	�q�RF��*�F���uqoXT������]j"������D|z�ղ��.��co�α9rb�Ǎ��`!�,��+��o޽�j�SN�>�C�ױ�|���-}��F��;.`u;yn�0�z�Hm,
��3�92�3��{���8�Wl������u��/)<#b#�?����V:�����(�k��8%��;�����.[�X��q�z\���R^�C��6;y����|yΕU �0�mjƺ�,��n5DDD���|�����]�d�����6b��Y��+�g�Y��Q2t'"�l&w"�(=����5ɯ�]DLK���V�5�R�~$��?������0�ru���B����c��uS�I����6췸_�Z��Z��ol��@Wu����[i�����.J�N9�t�<��z��ܽu���p��s�ɳVW�����Q�@DD�N�����	�ܱ�v�#�f�T�/N���AS�w*�u�ȏa;��T���&�iFT�Y��S?���E#K���ظ���������M-�55�G�'���e.�]������b�z"#�C�^�a׎{�A�~m��ua<���l)C����0�<[�r���~�~?64*��x����sDB����������Y�ᥕx��e��+���o�Ƒ�%=�8���7�1�%x�k%"�H�/q�P��׌�M�9��pZ���#9H�������c��'�G�Ƀb�����ჰ�L����$D\= }����p��M--�e��ve���� U�B�,O�t�j5tx�����l^o}�w˟Y�BԹ�&���������i��X�
�������i ""�)s�0��⵻ajr���m�������{J렩ސl�� ��������S�QQ߈J]#*t������'[��I���$�pԺC���tQ)m�a��L>9tF��Z��6��Y��%�V��5$��zU�z����'���b�����l�e�.�����
�o�7&!
��B��e;!�]m�h��_���]z��*ܹ	%��-#�!:0 �u�V�~�q;n���s����W��y2stl������'T���W�g&��'Z�7ԗj��{�ڞ�v������v"��s$���&J!R� Ixn�ad�^��
V��q��=�½���*KP^]
��
��2�ٻ��ہ��
�>v����KK��YT��8z���NL�A\H�t�Ҫ���b;��	i��{�
���j��[�}�C����9�]{�;ދ'-�:�Q�g�Ͼ�ZV�k���|��߹��]?y*��}�{r�m.��u�x����z�h���ʼ���-s0���G}A����h&�r�4�Roj�p���`�8A����<�Wn��:蓖��C��D�m,|5}W�^ר���� Bی`- �a)v�u�[ʈ�tW�MM����钑�������]��Ř�m?�<&_ϒ�:�'
J-~6t�pW���6m�i}P�Ԍ��&�66������)�Dny�����w�AS��s��qx~�!/��:�_�Y/�����B\^�h%��U_᭯��\~��t,f�DQO�(���/~&�T����02.�W_�n<��'���G�-���7�Je>l)CD�w��+�����a�p'���_��O��Nlǰ�f��g2�'����|�>("D���EP��s8�W��� �t�$�0�j��f�}�.n�$}p��b����������΁SRO�V�噢r��`0YV��'����?�wϮ�mwy�_���;�S��-��~!������E��QϾ�?,�������F��:�z�f��O�lDFi��ۈV6Ϛ��������4gh"�9��Z�s��b�����˻�I�_���������ZiJ��5q��j+xP�7���p0jj�o��:ī�t_���_���sS۾�z�"]����������|��o_�o�O��]38�������c�X�>��Km����6R�Z������֪��c���F��M~il)C=eթ���j����_��7>tx�/Z���eMJ�Çw܌2��;޲��rqՉ���m7n=ˆ���X)4o%Ƌ8QT������S8Yd�b/@�����@T��wWI]=����n�U���Ъ�Eo�v�~��]��K��ǳ��7f���<��TL�p��T,9X��uG�.Bv�n�:f��l���s��	�MWFzby;Q�zz������D���KW[4>��ڼ�I��I���d��U�o���,8�u	���5�(F2�u��*S3|�z�Қ�Uڏ�����&wѿ�����b���o��3}t�L3l���E���d�w�L���߀�����qH��l7!&V;/ e�'���8@����Us��zJ��o����$mG=ލ�inyZ8��ux��Q��)��ᅽ��I=��||��Ij��^|t�rLJ��;5��CeC�[ש�륩+<!P!""���5��]ǤI�����Ic0>1C�¬�y�H\q�WQ+��9q�L�O�:�H<�Ӵ�ް�̖2DD���q��#b#�S^-Ue��)�h1Q�"MDt9�n�hԠ��_b�c���@O�`���]^U_���JT�UA�X���Z��P��������̺}xn�A��F}�Ӂ�Ҽ�y���I��H����x��r�]|}�	���$R�b�0i��u:�/q��Ķ��} U���m���UCu�������s}v����k󁎑A�(Ok95%�=��8}u�R�j��m����=���,���s��yZ��'&���WUM��D�4��ը�(��j������>oqm�t��\xM��R�l�C`�ND��D�.&"�\E�_� $l�#H��P�d��B�޽����vtD[��No��;Uk�6���$Ч�$�y7S	u����&ȼ���yx:�7�t���S�����u��4���8�RE�۞C�8�Ѕ���U�'Żm]b�����bVr���+�VV�m�3�������3W�鍮�ӌˉ����}��
����&��&"�D��>��Ď�Q�w�t�&z�
��]���s�xo:�'��ANe�ÅQ1Q����X1:=y!wK?�p'""�)^��J�I�B��������Hv�F���)�|�Vw��\�9j7��F_������������P��Je~��q�ı�~!��f⫳�YV���&&�bQj�y�ɉ�荎�b`��N�����+����͛w��!"""""�`S���[hTJ,�,M�^�Pj�u���U�4���"%"�!!R��ޖ�o�DDD�9��9h*y� �Fj#&"""����]$�&����֖2��5QQ�K��*�vX!""""""""""7��]�T�����9D��x�Q?�5�{��v�\DDDDDDDDDD�v^����Qj��I�~�t�ĝi;�]k��`�ѿ����DDDDDDDDDD�n
�	�
�DDDDDDDDDDD=D
܍Fc�?��!"O�my,��_g|�/"�4�U+�7�P�܂��&4x��������Ȟ�
�~���;�cj��ą`F\0���C����g�uX�[��f��������Rk�C�����;��"�Q^߈��f�1,CC���V�P`td ����P��Н��.{}�I�?�"GT*%}4�G�K@DD���������
���DDDWD�_�ga�����M-T�P��]��<5�A߂�&��\o0��];��b�p��
�
�p��ƶɈ��}|8DDDDt%p���l)CDD�%�1n(�z�t������Q���銚�f)H������gqM=�;��w�@Y]����������777{�h܉�ȫ�j�o����-�7��-3��
p�R)�J�PTcy�[T�?�a\� LI����D���H�D��O��׌����='��w"""""��IƄB��:���j���U�F��#
�Ң�(}�|<�]^��}Â�
?��58[Ta���Qq�U+a0�P����vWZ����������;y���^5d@޻�:�F���;c�!y~�q|~�j�h����`n1^�s�������;$Q�������34|�	�W����=4g<�v2���ѤoA^y��-ā����Gqu��m�����I��ԑ�R���P^^�q�?/�-�����	Q�����S��R���_<��Z��`DQM=2K+q0�/�8"]��]R�����ϙL��*~�\DD�UF�E`�w�!2�򀨗�����=Xu"�˕�b�d��\i���?-��iɱҲ�#����WWKUDDDDDD$_=��w��h�3{�U�HNJj,�vq���o����������W�'�l��̋m˞�~�?{������G�� m nxi%��m�;�|^E�TY/��E����&ań4,~�S)�����t�hx�DD�5��;1_<x}[��ugr��7��ҹCy�X���j:��l��;XS�c��p�lV%��V����>Ó����A�6o�QX��^Y��Z��2�R���Y����|#w�>�gf��{_���l��l6ɒ)$��H�(�������?��w�@ !!�����I6�[�7ۻ�޻�.��;^ے�ʖdi���K�6imy��|�a{ek�����N�[�ZP��kEMGo@�����O��6��u��gb٦��l2@�d$�Zp��w�s�ֵ���>��w,���\�����K2R��[7�?��P�|>�{v��
�9Y�gB�z""�!�r��
�����=�VDpQ)�����]ӌ�|�:�&���J��+�W��������.~��:pۯ�DEn:6�.��n�8t�8��~ḭ]��Xs>���_�m�a��q{�����%C����˟B�z�*�x�m�����(���8���ux��;��(�~a��/�2�{��f��P/7#�I�d7�L5��,E϶��=��p�f�&j�Ee���|;�����p�o��K��	�ғ�+��C�8��	""""""�"x���Auk׸��Ph�a<��PЯ�� kh^R��I"d�@Һ��l�2���ܲ߻~�����,)��k��b�tmmm'�f�~I�\��Q�#��%ix%��D��C���z��=���N�><�SWI9�:fu^42��(RQ�'�֮��:�����w���-VI}��~�I}��ϥ�=h��H�A��8��M,���-~Aa�~����0���{A���;ԋQ�&�s������ns�����u�����Wo3���NJV/Ũ��.�����y��<_�o������n����U�Շ<�<���کy��e#���gADDDDDD�cd=���Ό�X�F�<3u���G�'�Z�V�i���h�m������8m�}>x��w�Wtd�.�r��P�.�	��Dnݑ���3��(�&�i�d�'I,H����Wx]�������냗Jp_̢�7D ~��uk����m��O�:�m��=�����s������l���ψ������l^^8�豦�I��g{�~����s�����Ճ#����+���l�ϕ���]Ϩ�G�z���U�M3-�S�I�(Q���(B>�t6������v<shr�Ჿ����KO�=�.b�NDDDDDG<#z������ow*8=m`���s8q��>�G>q=6Uݞ������م��{�WvbdK��*�S�pӒٸy���j:zp�yrF�^��OTQ��-�#""�F��b����	j �H�0�q��Qܯ[P��d��ކ���c1�q��2�g���j�NӮ��Q,��iwy0q&� ��@��Q��������ŗ�\���yL~�������xyg���_&�b�._��+�r1����v�<���j����f��Ϙ~$ADD�����yQ5�ԡ���K�A�����r�<1�
6�.��O���.l~^&��u�M������u��[����(�F���n�!wV�eT+�`_�g����N�YI�K4�7]E���r�*<w�
��[�|��J�i��5M��cxl�q�Jw�wx��yQ&��B��lš���0�u��γM�;��.Iz�ꛆ�o(g�ND�$�aT�.���߼~=�7�c{e�����j�G�����'���K���^8�2{��/����
�,ia�'�.�W��e������mx��9�e�	�����d��_va��$9�i����P~r����M�&��n���[=+DDta���;*l����s�Qԍ�p�h���g�cw"�dЮhż�wA9���`ۡ��l�"�(D����}{u=~���n@�́H�܋1Ȳ|F��""�8�y~�T��5���Ce�%Tut��rà�i=܉�hb�ӆ-��k2��jݪ1�hԃ���(�F�p����aS��u��|�v}�b\��o����=~��Aˋr�����v�h��V��o�y^Y��쬡���8�[���m�n�?��A$i������D<Q�܉�(Ne$���O�u!�D��� �o�Bin&�MFE�-ODDc�!��6�]���׾�C��������-�n�=n���<.�^7$�C������޲�5�9^���n�Wѫ��1�}������Eɧ�<����.Xn��� "�����"'�gbMY֔�����}-���賡���������C������`���I����Q�g���EU[7��}���Nu���k:z���q�rܬ>wPg���[������5+Q�?|F��@ݿ���m@�`h��$I3f�{�^?3�,ь$F\T�
w	F�==Z�.6����0""-��,�ڼ�q��~��o�����.[�T���wv���=���v��{���hU�3�&çn�ԯ���tх-+�ŏ�
9�o�'k� �N����[�,������]V��g���s��{���y�=<�����l�f1�����i����s�>�iבq�q:��4�X,�e9DDDq*#a������m�L?���߶��yޠ�J��h,k2+��������?�ި~�z!�]�2�@D����̓�Ѱ����<"�9p�	���/XQ�����P����́�2N�;��=�618醟�_�j%�Z�@�u�x�H��zf��ƀ��iF}wr�,���b��T�QkGӠ޾��n;�����^S����ns�^�pl)Ӈ@Q���DDDq*�4P��P7l�},]�/��&�""
$��9��U�+�Q�␩��u'�]8DDta.�;��i$��ju�^�k ��7�ֿ��6��K�Q�����-4mdF�:��}}��}�c�b:�ڃ@��U��p'"��e�T���"����o(u[mC7��DD�\�߃��I;ġ�~S�v���tL�V?�ߩ��U�*^���[b� >Y�G������`�Y�-��b���j��5nc��h�z*�_$ ��M�O���]�כADDǌ��@��~�9���ep���H��>�_��a�L�b0BgI�>1���y�� ��]���e OqG�k5$hg�9N8��`��n[?|�)��}�"$�|/���B$��鑤��Y&�r�^�?�Ni�{\���3�{~�C[��u���2��IQ���dP��<��hR��+�Mz�����w�U���t�}W{�mrtu���%,f,�~����`���۫3C�Q�{{���_X~��3!��"Z�ܴx6n]V������xl�qP|Ѷ�L&S�$Io#�x�ޠFVS��{���8�RR��JIꔃ�2@����x�����m��|�:/[��T�2C̫S��i2b@_��S��V'�:�dY֫�Ɖ�e�:ec�L"��x>����������(���DD~�აƔtx\Ρ��]�T�&(zd�^��P�-�0��0��	F�:���]�n�3��D��dug?/��l��8����¡��8�V���'�����:y].,��vi�Io Q���Ϋq۲9Cׯ�W�9���/n�mo\��7ʲ�(�}>��S&���l2���&�s�ͻ05����(Hl�V�<�ڃyq6 �*�' R����m�w�x�Ӫ˭.��{>z]����9R��NgPV̲v@CN?u������K"��F���R/�|��������Z���ҟjP�&�3Šw��t�T������|G�10�� N,�o@7���g���;��v��lpPRQ�.�'�Q9u�[����uDDS��uނáyP���N�t����7H�͎$qML�>�Ð�3;���h:,+��}q�2<���5����_q�o�+A3J�W������4��޲f�q�A?b�vE��V���p%��q�����v�k[z�9��5-��g7�� "��|N��+-����W �݉�"inN�����3p�#�?ߜ.
�8�z�>�[%�	�%���s�P�j6D5p�v6�#o"""���-w��&�m�0p'�Hk���\�c]���N��0�DD	6���r�و������`���Ȟ�DDc�ڭ�W��M��B �DD���Lڭ6d$�n'��}�v����N$�4������$å3F���+��冷��]�Ex w��S<Nm��$�&g�iL@41p�`���,K�Q�}"�a���T���;����<t[�=ڝȈ�b��6�s���P��jX7"�)�U�����-�ݝ�h�
�:z��WvboMS�c�Nr�N"��d���4�7��EgF����;e�M�^����������j�ne�� ��)��w�sg��H�����$���D��?��9Y�ND��ܡ*�h~kK�p���j�G=&��u�!{#\ǌ�^�:��M'PS��	�N�)Xcf��SDD���g�ZR�������|����C���;���F��ĝh���ܹ�BD��Ts�6�$گ�:�i�u��0��Pq�4,DKNŴ�.w
�O�$WE'G��W��E�DD��Z���S��˒������]���ԕ�h&�o'#D}��h���%Y�ND�${�(�܁��VPxI�w}~�aV�-��>~w
�"��u���h
S���%Ѡʶ����d�IVd��φ,���l�h'CDQ!��k���#vrAD4���߅��9�U�(ڭ+^��:��Spdy̟)�w�XDD4�ds�VE.��TQ�u��֊�̡�;�6����F���hD�nTd���D4���PY����$��,\3���G�u�SPd��c�Qw�^�NDD�D��^]+֔�bQ^&�R��mE4��2f�]��DD4@�FnF3p'�n���M���h�ha��w����>y'�4%�3� R/��2u�`̟Y��	wM��m?Ӡ�H����G���z��_��i��=V�W�~�DDC���k��M?�烤���v���G�h����OI�.$2l�
��5!NCdڰ�/
E��]�y�Q�yd�	�w�2(���]����atۦ �Ĥ$�&k��;	���\�S20�}}�|�-e��B1��{r�������j���@ѡx\�uv*+6D��w
�Q�>z' *܉�(Й�<w��,.G�ɀy�
|��ӾEy9ڥ����0�`���o_�v�'*mAD�Mg2���%%DD�&k.�ډ��om����n�DKNEؗ����"I�1�j���!�}�""�o��K`P|����Zـ�������X^���X�������A ""
�d���f-ѴS�F�R��Q��V��1$��(zRr`7%�u��)$2��W�K>��!"�Xc~��>|����r���������%�}iy>��ka�)����O��""MW��������(*$�A�ԫ��DD4���>��m�):|>�W������]$� "�Q����rN!6��#�l�s�ވ?�2ޭn��k~r����V�{��;] "���W���s��8܉�A� �,�嗁��f���2�SP$I������<�:��DDc�x}��O/�O݀��9H4�̽7�[�'������D���66�����?����ZADDc��fW^����EK%�N��� �'#"��t���1p�����Jc����""O�݉��E<~�uXW���3���V����7���UZ0?U�	�w�%���E0�6+z�׼�7����Č��W�!�E�l���j3��.���(�O��E�<�������z����N��E�%�}�gϾF8�SO������2^K����vфD ���>�o]�_ڴ��}>/7���f|�m5���)<��4����D36�)��KթX��j��]��ӭ] "��tz$�|/��y��3U,�;!��{��"�b�#3��2�9�.A{/搖�h��S�unV�S������b���=܉�.������؍�O���ׯÊY���e�������n��pc;�7u��ώn�C}�O���l�cvf�kϑG�}�������p�y,��h2��t�Id�;�t�̡�VDD�MGZ.�F�&��z��H3=�z�nD���="�`m�n��~�nXP��o\�5%yC�Z	fl�]�M�j���='��G��mM�ؠ��.'ź�ګ+V�9�p�⛑�_K,1p���<�~�N}��e��p'"��x��m*�H�mK+�qv>Ve�b�_��g�{�Ve�<Y�W�ׄu�U"�K��������"/VjW��Z����������z��#pw�b ��M����>m��+�SQ����d�-&�1�v�.������g������w'����6,�Rf���V�SplN�#i��G����?��(�>���������(�H����Ex�*��)(]�.{v��Q�{hC	����@DDDDt��XeKDDD������[	���7�-e�Sp�{��9�ɣn��쩈��� """"��J,�"����
�𮃏�;EIe{�rEyި�G����#""""��I��HDDD&�!����ñ��[��6w
ʎ�ִ{V��C#��?�]�'��r�#"""�J�F-]�� L��0-,B|/�og�NA�q�e����+��|��.��V��z��
w""""��q������!���=6�XX+�)��_������kV^�^5��N� �]�E���D���="�����]�c%p��`#��3p�Iy�ȹUn�o[����"""
�,���I�D�X�NDDD�K>y{X�K���>��?V�����{N����j�_R�����.�����܃ם��=�������z¹>6�g!��hRJ2S��`��sM�I�:wX��MNr�����߷��fI��=_"""�i#�<Zۭhk�������N'�b�#5Մ��$&���ȱ1X����ry����aG�ͭ�AQ$$X�KV�		�q�1Yh)#1p�)y�T�ruŖ�l^P���$<��$�Է��8�~�U��g'\ޜ�t\3���r�vLsO?�U�c�:y�D��U�q���h��Gk_?��lh��Cmg/�v���=� �M�و[�T��+���N�m�²�D�}�Z���[mڥx���e]W/�����#X?��r\�����[��� ���;ap����B��N�5����,����p�d�RM(/KGNVB��\��g�u���o�}��n�v�x�x/e���β ��}�/��1p'""�#�K��o7m��O6����$��9�P������Q�'���;6�������i�Ə_ۍ���u_v������=v'ޫk�ן~'�;	�,��B-d�i�l���<�<������{����k�����G�֩�qPk��,.��?�v!�u7�hf�;�Te��t��>l��c��-pw��Y��:���V���]�%��iW�&-pw:Cl�)s�T"""��8.*�Ǔ���=��E�xp�{�Yz���1/7}�6��U�msLv�vyâ2�������/4U߿xs/�7�c�|f�-��8��r�#�߼��^	V������Xɡ�1����n�u��;�-�j�n_�k��߽v~��^�<��N4�H܉�����l����T5���ٴ���N��H-��!�C$����M����H0k�+Jr��������uZ��ܡ*|�w�ms������ڝ��WCu[�v}˩Z�n��/n�B���`B���1b�sD��On�\�=����i����_���'k��9�u��3�:_������P��XJ�.4����&�ߋ�=A�t�٨].��u�`�hqr��?y}r�MW�ʺ��}�û��׬��Τ�#����v("����2Sq��uJa������M��a�N4�Dw�h���%DD3M%""�	��2���W>�Z���Q�=��0>�v�֣\��K�q������LFQZҘ�{�W�G���_�Zʜ_��_��v|�����wߛԀ������eڼ88Q���Ϳo^	2͓�̉�"��=""""�V��D�+�mΉ���;�h�^����n���{q~x~����bg�G���}'�^��Y�����Ӯ�C����Vj�
i��	������p7����pӒ���㯍����|��_�օ�?~T;H���7`~nnYR����p'"""�~Y	�2���_������Ǫ��߭��`�W7�Ү������q�����o��'��v~qە�fA�֚F�*1��h�t�p���R��������ϼ���=>��E`��5��?�<���?�ލ?���߼Qk+���h��ւ���hڹ�	7�DDDq��ٕ	�
w�7������}Z��h/#l�W�w��O�ԟ_��ʺ1���YQ!/��~���j���$l�]�^��sd����R&|������s��4O�4#I&~��͘����_������T�'�C���I�.��D]������"���(J��GD4��&e�}�܉����/�6��?5n�zko���{h��Wׂ��yfg�j�e%��ħޏ�|۪�/�N��8���ꚇ�����U���kqŜYx�h5"�?Ò�h5t���C����g�j$~v�&�JOƿ\�G��⑱�ߍ�ʆ�|�
-��t�i弡�oP�����[��<�K\���þ\�DDDq����O1�|�I���0PQ���w�e�m�e?�����K��!Z̬�����yt�q|��G�����e��!p�̠�c���Î�}���~fc�b5������l�6����;���
w""��g7%�5{6�Z*A�לS8h*M�Ư�HEn����M�Qw��%���]n��3�`���C���^�C�u�Q��7Wz�N|繭c������]����H��|��!�j��ǣ��ዛ��"+M�������,+����\��y��dіID��DDD3�����p�Mȫ?����t�g�!�ő�n�Vq.z��oA)���w���8y)�C��4Nj���Du[7���&���¼�q+��.�c��9�	�c�@��z%��J�����lG�v)�-�c�p��Ҁ�o���z⧘�������X����?�:
"�s�"��"��ל;^�oA�a�{h��gKWE��]`�NDDG�>N5w���,g�೗/ǯ��xL^�p��lä_C�)��<����C�s�|��o]i>~���H6��}����4U�����9i)�9]�}�
�	��%7i�,�g����y��e�݉O?�
^;~v�>�7_�*>+A�qg�N4���LҚ3E��sԭ ���ū~�ճ��iL@�0p'""�3|� ~�����7oX��e��VY�UK��IǦ�����Z;G�p!�=#�d�Š�Y�C�٨�E�����klǟww=��,�vA�V�^������0oD��GwG�-/��]���W���#�2�j�%x߼b�p�����A
�	\�d��u�ݎ��k���d_شK
���N���F=��Ƞ΋P_|nb���e����H0cqA��r���ַ�/h|��ƿ�x)>�q)6Vi�#OD��DDD3OGf	<z#��wC�N�ȇ&ϭ走�ߒ��a�NDDg���8
ӓ��ͫ�1���_�M���k�g�Ǩ犊l�"�+W���˾�f���'0��ų�i,��ͯ�9�߾{�V�����-�~q @�b:�ډ�o;����9h'�M��)J�uQ���[�����e��#��|��7�橚Q�]^Q�ǋ;zaT����o?�����ۮ�<��iQ��8h*Q��w����;%O�˪v@��A��4XP]�A�6��š���/��]�aqa6R-Ft��q��/��['΍�\�K\L�)�4�H�������Ѫ�߭�s0TA��y�h5lN7zN-��S/ۭv4�X�64U�]���8�֭�`q���W��N�V�]6;�z���hT'1�H�}V��n�u�J݇���ms��~�e�v�`mi�vpB��W{�'��DCw�"��?��~��|/��9�}^�,�`�N�X�NDD4s�%e���2�Un���3[��nJBU���iy=�DDDq�hC+���-S~�z����z�O����Ԧh�[ӤMSe�;��ېl6��jՂ��<ޡ��������7��o�n��NQ�c�;ь֟��ʹQ~�]�]vPx�'�kg�uL��;�6�S�"a2a���>�(�1p'""���dT�݈�S[apr Tݩy8[�>Y�tb�NDDDDDDD3�uQ��Q9wJ�wA	s��W��/���$���5t]�y�ۼC�e�3��I�ù���E����;Q�p�85o��uH�m��ާ]���Z[��Q�Iz�v!�w�ȁ����"���2�z3l�X3�4&h���ۼQ:���;Q�ArVK%r�C��A҉��m�/1�����O'�DDD4JiF�6h�D�L$h����h���ɘm=��K�kC⩭�K�BM�
8��3p'""�czE�¼L���py��j�BS�u���d_�j���M��O���Z&�E(��� Ei�p����۪`w�_���$��I�;�msh��s���o׮O�Q����!�bu�Š�AQ`u�p��DD�4�i"�.��˘�fK_;ʪvB��~���ۊ�G_G]�Rt�Ϛ��f�NDD�Dh��+W��/��v�m�x�H���6?��y�XW�?��E+���-B�k�Ǽ_�߹n>}�b�t�=m.7�v?}}z��QϽ}��yci��ǻUuxx�1�}�6���D|^}�￤\���I�g��Vl��� """""����T�����C��/>�F{��L��2p'""�3"l��Ǯ���Ƽ?�b���K��0��9�'���;\Z)�+HMԪ�]��X���Y����FRd	�赸��_}~'��g`yA���b�D��}��cSEn�ݳh�����[.$���N��֥s����UZ�x� *���V��������p�������x����'"""""����v����x:�uE��+�g61p'""�37^R���iU��Z�f���צ��i�iA�D��;K�E[����_5�X�,P3��������ub��d��,*���Z���$,.�nވ{}%���<�T���j�4�	�	�^f&������J���.�ۋ��_�ً�����n��?o\�UŹ�}�ܲ���>�؝���m-����zDe&{�*�3l��̖*x�/���ň4�DDDqf}Y���ܴx�V���.��f$�Q���͋����r�?>�7�h��իVi�M����=���4�:ro�{=�d�K�h�y]W���Y�O1��7p������E��� ��2�}/����Ok���-�m�����~�DDDDD}:�e��C�����R	���֜�}�DDDqf�Ŋh����7�G������TE��������`D��Aˋw�Ap�h�"�����c>�W]�ｺ��}�v`@�����C��w���4/g`=�ky��9�������������O����v��4}���nJDoJn�^��;Q����MEX-���ڵ�8��~�m�щ�e��g$�����䪓�0"p�j����=�֙���K�3w�~x�$�XA/Td�a��1G�p!�_����=Q$I�~Ii�.X��@�K���݋���`A$0p'""�3���'y}�:�ŋp��B������{�5���T�qh~mIn^2[� ���~����)� w��Ks����A	�����I������2�D/��>z��c^x�p%.Ŀb��D��Ý(*8�M7	>�:�I=͠�P�N�T��鹗��m0��;Qz�T������Mq����D��[�g���������^X[��M1�+ܳ�C����q��a�\��hזi���~Q�˒
|��K��!�<�T��A��{��p'""""�����3���Q�.���M'ќ7/��f�NDD��ۺ��?�����߀99�0(
~z�&����ן~{T_w��u1�h�_h.�q1�d	�Ɓ`�7AY�D��Y~���\�_@~��R\��T{���2l���Hze����w"""""���i5�ؐ�x=�����N܉����'�a��Z|r�%Z?w1���_�$�����p�U}ۜ�y�W]��#�0;��m�������?4h��ۙ	�-j�u���?�+��p�Y�F�^o���U����y�DDD�휈hqw$����aBo+w"""�<b��T_=~�~��%ia�����ͽC�k��]o춎�����Zp-K��� �Xc;���:Q���4<8��ma�������C_�
�5�����6�Z��W��;*���#mw�ADDDDDD$(gؗ�����h9�ލ7N��'�.Ү��*�l��o��s�G�J/�H�kD����x�%���D�{q�@vܿp�:���~��^��vAj�?>�+W.Ղ���r��8Ǜ�/���mw�[�.�"�M?���,�DDD3�s��]���M�T���[����ܟ>X��ݰ	�	[ʔ�%i��;����`�lG�viw{�gJ���BR�J&�u7�y�����-���H�]���w�������%�C��%�(.J�M�}�N	�E�֝u�E���4�K�BZ�֝5!���ρ�;Q�Y߹vV�䡶�Um�8�ҁ�͝�n�҂�5�}7/��=��φ�G�A�;�����s��3~��L#nZ<�~-h�>��i���+��������p���U��=?��'��r�Ͼ3j��Z��Ăb.�4ྟ����Rq��C����6m99�э�~;�,&V�Q �p'���Ѩ����Ѡ@�W�����;�C�p�ś��Û.�?��ER�w?�- 饣��{��-e�gU�?>�m}�Q�=��(*����˗aUQ֘��w��^5`����^��^��;�>Q}/z5t�qQ9nYZ����D����3�g2� Q�`�GDDD�-��hf[?��NDDD��x?c/�ݰ���k��u���/ڷ�x��ܲ/�Պ�'�������A�rީ�7�����Şs����Vca^���"0�t�V�~��u��J�׎�C�a� ������Onل��.�`�.<��0>�b>:� """""�XIR8b�X����^B��DDD18�`��N�Y�����]ޘa�����￴K
�ǽ��CUڔ���YiIZK���Nt�.z��ͽP�$�X�W��^9Ok1S��5����6�m��
w"�U���$""����_��m�x/���e2p'""�s�G�&�w���cԶ�Xc�'��G�z!���^�/�����z��/l���@DDD�.�"�IG���� ��;MѶ%���]�`��Ql��]N"""�u�h�q{l��w"""""""""��Q�Qw8B���5RL��	����;�L1�M�,�+��R������(qי������p)FF^��D��;��(s��1$Ԋ)�2p'"""""��X�����"���aX���p�2B|/>IF�1p'"""""""""��pT���S�.ˡ�ݡV��"�a0p'"""""""""�0b#,�b��L�+�}��pc�NDDDDDe���KDDD�#�#pq������m6���`w��@]���h�#-͌�LL��X��������AK�m����\p8<��|��$���bBvV�:ozN��^V�]|�1f�`H���DՙN44���{�]�v�5�����,f��!5ńX���g�C]��9��ͅ�;�zq�T+2��{IGf�%�;+܉������M%""��t�@���6T���s|hj�jSɬx����!���)�^:��� ��ѯM��Ip��!�+܉������Rl��Q�c��}����+Su����б�sQ�*�p'"""""""""��B	�cM������n܉��������DDDq��c�[և}��i�,=��.Q�$[<�0�>H�i�~x�F|�٭�s8ADDDDD���7""�xǿ��ǣ��E��4|x�|<u��>]"""""
]�C�є0�"�i$I��k�^��4I^5��尺4��;Q�|<�sX�NQw��2�rUI���������(8>I�&���kb�KgDOJnؗ�����j6bvv�6��8�,���Qȸ�MDD�<�5��0�z$�����Y��ֱ�hnn[M%XY���M��es����������u��W���J�(j͙����,��;� 51����ञ���7��S """"""""����
!���uf+ݣ�79�"�|���1�����X�FDD4�t�ς�@�;C�icMHÙ�5�Ir�^��;ͨSBz~��"""""""""��!{�(:�(��d��� ��H��;͠����S{�	����"""""M�^6ьԑY�]2t�,�)	Us6���#�Z�)hF�p���o���> """"""���8Q��]�$����=D�~z�ep�M��z�)h�߯���؉��������¢=�Xӥ���ae�����2�u�i{M�4%܉�������x���MPT�xN�l�TTUl�ְ]`�NS��xADDDDDDDDD�ӞU:�^��0t��~K*�E�i��@�����v���<�$��= ���������(��2K��d$��a&��:xey��^Y$e��nEI�Ǽ�79����c�NA{��m"""""�0cK""":���Cf�Hީ�t!�OVi��#{\�/G�d�s���{�����+��p�nJBwj�I�Q��DDDDDDDDDD1�ഡ�Ի�%�KL���ڔW�i�h(�N�y�ׅ�;M��D���eADm�U{ yܠ�B�G7��Y7�J��e�YkWB
l)9 ��Z���hf�;�Q~���![U��uH�nBm�Jt��O��3p��]�|>}�*m��w���G��+�N�I����@m{w���F|��uHO2����(��+'<U�(\z�*��-e���f4�ˎ٧��Ȱ=lD���]h̟�������)h	
�S��ճ��wQ�����"�b���6��ߏk�_�a��L3��_��W/����NDD4��b���b�uQлa��

7��C�3Ӂ�;Mɂ�����t-l��ҠSd%�qmQ���m�82's����hFa�.Q�|L����f$�ہ�[a���"'������P�8�����������3��6,.��ݠS0+3+}CEm�@�X�DDD3{RM�v""�G�vb��wa���"/���ϋ�YK0�8T�����l^~v���%�rn���@!��(��z�r����������P<.��~&[7h�d�V�+I�/Z��`�NS6�0Gܗ�U�٩з����aAi�6�����h���~�I`�;�L!���S[a��M���*�$9b=��S�F���W���D3�2Rn/�JEK[�6��_0t��}n""""""""���[�lg�]���h�S[��0
1p�)�W��EE�������r��*����ng�;���z]��I�2Q�����z	�NP������`Fc���.��;m�NsnJ._P6�qi�7%᮫��9h*�ÿ�D��CTDDD�N��`� �����[tw
��K�y�G���۸�MDD4��?�:�""��"�����Bb�)A?��DDD3��Q�"p���;M��]��;0����T}I��`E��L����q�5F�.����������Q|�h�(x��!""����w���v֦X� 3	&E������x/����S�a�ɘ�>�N��kj���K��3��_lO_<]���z�~+�br���t��rjS�����7h�l2C�$B6'B�)iP�i(���H��:�t
�:�dI��KP��)����p����O����W�1+c�;j���;Q,��v""""���(KGQAJH�ص��~'���4�E�!-c����)?�-e����Ue(KM@�|�݅�]���xs�� }-M���b���æM޾�Qw�,�X�z5>x�&�&!ŠC�I���1�����S�7#"""�<�'""�3���C�Rb�.�hԅ�^BM�}���S�q�c3�6*2r�ڤ)H�-��O�
�݁����dm#�4�����==��lp������О�s���Wk�.�����6��\��ݦ�����	��/�
d�^[��hR�,�0[,HINFFZ
r3Ұ���υ,��7:M���D��x�9#���D![?�nC�b���,�c{���I���D�G0�cbM�Ɉ�.��M;$E���M��ǂ]""""��
��\�l��B}/��Nі`��{7�GC��?;�������aIa����nU=����8X�:m�x1��8�/Qhx��h2�gǗ���"'�6�c���ew,��4�	�.���+�Ǔ���� �W͝������ۧk�e�S�L~�\""
��g""""������:5��2u^1O��~Q�:�@�o�^���uM@�>H<�ww^��?�3�m���c��p���̞�DD!��(Q��iǗ�""�OM�p�����"&ΈeK���3V������}(;��r£���˖"/%1���=V���(�HAv��X���e�ד�.1�ODtQ��� ��/DDD4��#o��;+�)�dj��
?�2R���ދ�9��+�<VT��62���ʡ�n^R���.*2w"��H�"%""""���B������;�8=eh���O��8�pS�)fc�c��.m�T�jf�%�YZ�W���67D����>�EN�7)Q�X�NDDqHl�JKFIF2���Ku�KN�I��2#�^�'Z����n���׊��Zq��-�R�ل9��(��@j�E�ۅ��V쫪����ȡo�a�Ǝ��t)��T
�Y���H�)h�_��u�㽗��71����w���z�6o����ŀ�-��]O;+�)L$�AQh�=J,nvQ<a�<�/���Y�XY��t�iJ˲�=8\ߊg���j�m
K�m�7�4;+ʋ1� ' �4+3k�⩝�a������=66<�8��a�NAG]�t��n._�
F�~�vq�񾿽�w �6销e8��������D���KD
Kv����f1vߝ�����$#� 2�UŹ�tߦe�l����ϻ�����rsS���Mk��S͘��3����X��c��z��:GT+�{8r��?�|�)h�k��#��?���ׯ�z�m٧��3ȿ�]�]�p��3��-e(L�Ý�(T�"%
&"���h��˗��Wd@�0;+��t�z�
������c�N���3��c�M(�ʀqĺ��p{<HM��0#5l�;XY(&փ�;EQmg/ޮ�Ŧ��1�?Tߊ���'�6�/�W���tpz��B��
w"��k����(n-/�����s3��uE5��o݄/���?�V�>�p����Ɖ�f,))x�Γ�Z��w���5���]��
�`���������N.��	a=`��r�Ӥ�/�Ć��d9���n���s���Ҡ������}�.�4-	�]�pJ�$N12�[״G�G<���[�|}m�"Td��5���>��v����|����ь"� """��sâR<p������%2"��S��$o}�|�����3A?�����8R��ۜN쩬��v��׊p	G+y�6���E[��6X�����Z ��2HM6!;+�pK�Xi)3V?z�Í�>tu���eC��pNv"V,ɏ��ca�N���\���;���VkGm.7�{�{qz큿 ��S����Z�y�5�n�w��f��[�u<P'��z//�A:���[�+P�����!-�����;�8>�� 
�< ���M�=�^�~�1Ɠ���ĻV�y]�z<�����'����ǃz��/p��h��B�͎$��஻N����F�զ�Qأ�.a��9��w��q����=�v��RS��� �2P^���tK̴��ο�ק�g}C7�;m>G���w�`��BJ��ŀ?l?�MI&��{���`�ۋ�����h��b�]\>���3��VhM�&œۗ���7m)zq{���S������uB^'�aᗷ]��ܿ�;y��{�g�[�N-T��K�����p��;NVk�wY�Z;�����P�ۃ�G�Q��=����ݪMy��2��Ⳮ�����V8���(�߷�<�5+
c�)w����#���_nه�&sߞ�D��A����hJ�7�(x���HDD�G�p��ۯ��Qt*��>��6���Sk1�O���y�Z?�}5�>V�"�jj
�O�7�GO�P���ӏ�0�����~��F�"|�DE|��w�a�����*�=!���]���;J����Q�W�ğI�!l�A�Eb�N4��IDD�,#��G>v�6�Y��U�[��i�>�aQ������q����>��E�"X?Z�p�^�a1���?�B���M]��ñ'J�kB}/b0ՐIl)C1LM���9�"1p�03*�?{�G}�}�;�M]�d�W�c���t0��!r�܅�]ʓ<$OrI�r)��rI.�r			9�!�^\(��q�&�V׶�ggT,Y���f�[>o^îfgFki5�����C�@ ���c  ����+�t���խ ȹ�Շ^v�}��ㇼ�	�e��e����;�r��ӆ]�*��:n��X0WuM-��=�u=��[w�SW��w$mޔ�Z<w�{��՛�ʆm=�j�lm�S�����;{�N�:^%A�o�?�4����#3ZQ!G�`P(���* @�Z4s�ۻ�+�aW�:_~�W�q�r��C�����_Y�U;����ߖ�գ�y}K�L���k7�X���Q^��>��
pw$m��*]}꡾Z��aŅ���Η���_0g�.9�}��}��<78[��U �T� �y������LO��_��<��m7��ECݝ���/^���P��4��{|����]��`s�Rɠ %��R�bڨ�_���}~�8���]�KB]��t�����
<�,OZ��
 /��  �jWΝ�i��n�:BE���\��hL�~ߩC��gO�1zy�Τ�w�R��v��0�Q>0�1(SGV����)���Sf��0R�OюQ�ˋ�]��/w7�8�d����E^   �(;��9��7]p���=�8������PC��.���7�U���LD�;2Da(�1��QW�sgר��Н_�k�j�ڶ����[���xhF����i�� �](pdv$�\W��1�����rٕ�dx3$�KΨ�Y�u8���ħD'tw����Ń�ϝ6�Duk]�2�m�d%&ӊǞ�J<P9����c�f��r�E�O�1��������Z�x)��0�%<�=���6  #4��+���n6�{_A���M�
/Fg^& =]{Ҍ�lײ�K�~��n���KN��q{>p�4����Nؾy������xL8�m�p�TN�|���YcGh�;[�p���7S�}f��V����k����+N��D��D.��i�����n��5Ǆ�)�Ƌ
��X�?  �B~���;%%۶p<���ro�䔙��gVd�!PS�pm�v�j6,�?���c���Ꚕl���6s��>m�
�=?�T���C��=��rwНҵs�[�p�wl�*�B'  p�{�N��hDv�U�w�(0�Dh��f���k�jN���o��xݩ��4{�p��U�L�R\���;B�XDH��c���Q�S�}wڬ1�u����v��E����9�m�7��S�L��  H�y;�;p,XAWl�zw��3&{�׺S�x߻�4}��W�����3�+w��,��;kꘌ�-Eôa�9���E�mBz�3K{G��]R'wڰ��^��;9������=���c�v��z5�ء�]�Բk����)�ȊF�oc1KK,+k�-���cU^S��G��I"  �"�+�_8&,g����]p�S�h�W�ۭ�eE�TY6���������"}������;�Ϟ�͛�yѼm��)����R&
�jӌ�5e�"-Bj�5C�G�J��!pǐtos8����H9�;{�S��p��W
��-�����~'���R�����w**V��46j���[�F�׬V���Ao+TY��U������*TQ�|u�[��ͧ���ڗx�����3��@ߏm� �3�#�Q)B�p,X����V�~h��.'����˶��տT�
Cz�ӗ���|P��L|v��IS0M��]ϸ����+��T龰f��m+C+4�B%n����/*nRcϨ��5���|/wd��pT/o��ɶ��������S��w�2m�9խY-ۣ���:�u��˵���4l�4�<u�F/\�`���8�ծ�Vm;HX  R�AS�cιؽm�O��rzJ
�w5U�TH.2|kg����15���t���/T�nvk\}B���~]��j��{-�T�;�~�}Ʌ�Ή�i#*�Ξ:e�H�Pf���^RAk��%C;��}#�*]ܑ�'�ڠ�����-��Q���u��U[{T[�|R���W�'�	���;���.�;�\M��2VW+4Eb  H��v6�;�v���t%�m+.����ѕI-�fw�.��#:���yС{�F	�gM���z����q5G�����so��Ɇ�3F����h��35e���{!�h��y�/�����$<S���N��,��/k�r��}D�=�7E��_um%>�n}�	m{�)�^x��\}��F�T.k����| @F��U�웁���񚺟���a ��Y��rN�y]K��>�����<�G>}�&W�����;�q�#gM��>y�ۮ���b8'twں��E'����DجL�q�ٚ��e5��j(�������ަ[�&��[�9Z����n{��={��Sq��w.yQ{^{MS��F�.�4g+A��p  ��#ܣ�H7�8lL2����ɍ���8G�^���c�6�}7���J����бy���)�s�<q�����U�g�*{��3T��e�4�
�qNV�Kݞ�N�^[]#���X��d��0��e�Z��Kxr-pw�Ǭ��m{�ie�x$���S�^Z�9�p��jj�K�+���p  �@K ���EC��F0( ����*��>S�]w�n��)=��^�����Ǖ^xu��p��}v��w\��z&���k<:��צ�gɌG��|��P����{��s�"��V2��;�D_<�Μ2����6�j�{�������杊6p穓F����N���n}(�{Q�؜�J��͛��O�Km�3��f�֭Z����O|J��;O���%��/   ��,�P�n�
�� ���(S��C�E���O�����z�	�/�����/Ռ�W���n�Z}�//�y>z�a�cTY����3����9�o3�1 #J���Mש���Ť�r͛8J�=�$l��5���U�4��L7,�����/�yw�^ظ=��Ϲ�ȗ#�/w<��޾��n��l`��Zs�oԼs�f|�:�B$�ѿ  ����= ��#p/(��0{xq��	tT��xϳ����������t?R�޽���_xK_hi������:��=���"7Է(�C�c@�P�{�~�a�!}d�,w:�>�Lq+�;���}�7��6��ge��yDͻvk�g?'A��Ys���   ���  igw?�U0���U�+J5�:F����<�mr����������������2N�~��u� �v��45��P{�H5w��'N�����&��}ڈ
w�՟�6l�]+֦�鹗2e�ā������O<�l������_����[)�J�; 	�!pdN(��	p�X�w�
w�U]2��+N���kϕm��V�_q�#Z4c\�ǜ���O��$��%l�TY\@��� pG��+u��;�qK_��Yݱ�m�g��j�~�%�Pٻ��ֺ�x�i)�	dy�����������?��y��/
�(E,� @*u/!�s�n�Gk����84���V龳�Y���N��-�XJ�vGQ ��D�"pG�f�<�g뿞Y�?��v��o�ا����^�҇{���`����_�v1`fo�K���{�>�\��޻z�'?ּ����,|c�Ĩp  )d��8����fw;L�+N���t�[��}cӐ��U��(���;��0���p�v�s��t�7�;����5��9f���^yE�O����uz�~�?�)��[�   R���1����=drAE�7'�����:��;���̓چ�a��� 1(҃W�V:4Xꄊ2��Y���#+�����m�?����S,[�4mߦտ�uNd�y�U���C�|���&�x��N  @&8��ݶGf (��?�i�e����L�/�)���:!�)S�;��a�����G��@��}~�+V�o�2L%��R�j�-�J܏�J̰��hD�s?S,ܦhӶ�m�� H%A��:Cwg|�G��2�u��wy�;
�ĠH^iHZ��қ�_y��F�i�p���r�b�~g���.;C��݁Uw76k�zm�w ��1�w+ћ���{��6�s�*f�аiӕ-�q*� @
u�poݿϓM�E%*>m�
���1g[2cQe_,�?�;��m�!�m�ZV>�H�n�qO0q�
py=6���ۯ�P����[�5�u����_�s������R�B���uܝ�Q_��uzb��}�Ο>AE�����ҋfN�������<���m���{�v+���axկ�3~�ì��!p  ��U�=@����<[�����170��T8c���R�ݷۺ^V����xL $3c�}����?���H��vw����"��ܑ�҂��9;��N�����x�+bY�s�Pt��)����������+� �T*<�
�
�����v�Uv,���H�p�~ؽ�Nmm�:��C2�d�V�,��o�x�a ��|
�8ɝN�n��w'��Qv��P�n���1W���cl��ߑӶ��9�Z ^){�)���u�O�Ֆ��~���+�HI��(�"=x�!i�CD&���N�m������9?���ޚx���ny�a�;�<��LG�  R)0i� �YZ�N�|A���Lo[�t����1lw|��eZ0i�f�����{�.��;�����o�Tb�\���U���
N���pT�}�О��tp��#+��{����~^�.n3h*     DSTx�����7}����ilѕ�<�Gn�L5U�>��0א�H�_���N��!�w���{�U>۵t�&_�~���LF� Cdd�%g   �5�}(�����79z��iG}�.��!�C��p����`�#�ԇ3{���7�Tӎ��k��������?)��    �Hk��L��/8a�����?z��\U��s���B���s0�w��6Pjv���#
Uxߗ�+T�    �I������၇����7�O_�I��D�;҄����^���_^x�Z��#���\���ի��^�^Z�I�]�Le��    �?�0v�@��UC
�;m?��Y�ޔ��;ܑ�U�;>r�'�Z�i�2�Η_�me��4�������    ��ކ�!o��g{�a{�gj�đzi��>p�T����^�8��e�}��'V��yQ�t!pG����]�L8�i�v��}��q�D��*     5�4�i��~q���ۮ�Pkv���;o������B��������:�rp��az�#=ܑs�~�5M�]&okS��MBO�^=cw     �ɞ��A���W�k���c�a���Mt���L��-��}o��O�9�en~hP�����mҁ�9�0���׭]+;z�}�M�ж2��    ��m
��
�}'l�ja��H����3toK<��׼�k�����/P{�ڦVE�d�&��9%���2�K�R�n�Z���M�ܾ��a��fM    �'�޲�^�GV&���,Y��=�\�~����	��:�_��o\�����rN�H��`��t!pG�)/�y�c|x���w��⑰��mS�ģ���y; �a  @vY��`ҁ�����Wz��+�������n�8��?�X��q=�v������������_�M�k4n�"���w32p'o    䛍{&���/�ї|�߰���_��͞���2����=�l��<W���N5�1����ٕ��5���n�{@@��#�L��̠����:��a�o-{�(�    �͆�����~��;>v�.��;lw$���ilѵ�>�g��`�8��3��V��@���O������ղg�п�ݙ��5    �g��L.��څ��(�7]��;a���_�o�~$��7���oyĽ�����.Ra �hs�n*ܑ>��IQ�R�؈ک����O�r�t#n    䛷w�Wk4�T���s�4�X"�i�a�%��2��|��=ne���>�[4}��@���i)�t2ܑ�.F�+�������}$��&e"*ܑ�2k	    sD��ܾW�M���<m�B~�����l��T[�~W������/�ﶫ)�'_d�l�nE�q�B����2+(�"���e&BI    @�Y�5���qݼ�C���x�M}��e�|}�pƸ���7n�N��I�V�lY��?bm     2ǫ���g�91%�6�I�����]�	�������o pGz�#'|�2�a)g#~m 046��   �ҳ��-T�}4=�L�N��[����҉�i�7M/)���/_�w�+(�g�D&�;     5��z~�v-� �^J��w���:�4#pǀ}>]s�t�9e����il��ww�u[��ݫ���@w�q��������om쵌׹f�̬
wQ�п@i�2Qf��     H���ژ��=�hqG�B�����	H7wHa����aMQ�c��g��p,�6l�]+���՛�e>���I�U�XϹ�4T�˰�䂊
���i  �bȖ�D�%[�l>�  2��olз.9]#J�_D�E��֎}Z�s��t#pǀ|��9���N�N��Y�ܩ%u�߻�k�ZhiK�s�ZVƵ)�!�/S>�   	~;��xD+*⳨_qw���:t�bfb��t�Fǭ���S�p&�;  �8���}y���x���=����Yt��)lw�����kO���r�����Z��ǖ*Z�qe���*�O��
���L�� ��AS��BVDe���~�sB{�OL�W�uc�ϕV,*b�G"1j��|AE̠�� x�w/����9IeA϶i���Wa�ꝵz�͍�w$�	�O{��O����O-Wms����{��鶎9�sF�S|L�M�iy�[���6LS%�ǫa�f����㔉�� @�l�>�5nZ��A�mB�/��b�p�{ˊ�9I��h���
/�V��  ^q:|�����Ug��{]1g����E
��>�ڷ�٢��H���`5�˻.������Ow=����_^��ְn�nq�uZ�1}��ţ�n��W�3p�0e��I�	��b�6u�2�I�;  �Cے�^��2M�3��,�R`�l ��߿�Z9e�N�M;ؾ��<~�n������mخ'�np��#iS���oy�^����z}�ʳU]R�~���և�l�n���ڕG)Q9{��?��S�	�(���  �0��_P۫Ol%@f�н5
��3���`�����l��m���";���&Ŷ������_��r�  �Bܲ��??�'>{�
�G�^��N��8�ܑ��� �Q
�z�i'SlI�ܶG��Qm;Шt��(�W�9�m-c[�pH�����p  �E֭T������0fY���JE�2K�;n�����XF��}�4T���� ��ƃ��:�����1w���F����  ����3w=�?\�>�P���W?Y��(lw������A�1d�#i!ߡ���,�+��RK�}�('����g�}ޣqKonߧˏ��-���{�S]����04�ڙ�KKU6y��7m�>�e*�� ���(r�m�Uz�MnО�0۩�w&�e�4������{߷K־��^��� �W|k�~��
}����wk;a���@~ӛ��gϾ��W�#�X#pGҺ�z��j-���mK�(nۺr�T�2���U��'N��k��_{[����*o�9�k��M��+��P��*e�Q�-$p�&TY��)�T>�"  ��0����e��U�v'�<Y  ��w[��ϧ>��!m��sk�����Y����W��}Y@& pG���5��\�v�¤�^\��c͑���9 /\3͛A<RaԂz�Ow�H�Ɵw��f'SQ�    �!�-}㡗T�ܪ���Am��ic�酳=	۝���V�ۏ���2�;�V�˥� �t(�Gf�TUiĉ'i���{�7ֱ眣LƠ��Y�L   0?}v�6�?���\/)�@�Y��s��Ԫ/��=��=���I۟ؑ��}���q0=���2�e=~�"���CA�pe2M    �oNO�W6�ҏ����[���kٶnm����R�6�
�4��L"�8c8S���
w��'�t�D5n٢|6a�be:�v     ��T��p���7q�>w�I����)+^k�����7��Ͽ�{�iK��;r��O/	���Or����?���U�qǩj���tT���H   /,߲��k��뚓���5wl�B��e4��[�d�N=�~�xs��"2�;rJ�4�)Ӎ�7OæN����o�ARg\�1e�v     ����^���rw
�LMQ�)�e�2�"1SuI�*�B���Bj�D��,[�mj���M�Zר-�b�^��U붐�	�;�VUZ���Ebq�5��%�zl��jj�h���=�񙆊CA�$v�v�]R��=�-�\�f}�Z��oȶ,�1g�������P�#  �WѸ����w$�}'L�M���޿��7��_�z��)�4��T����=���5���Sf��W��C���/)}��,�n�T6i�Ɲ��=���E��L�>�!      ����2�jX��O�<Z��ׯ�|M��]ZX����3��Ȍ�^��իռ{�r�ah�?|Z�aÔ-lJ�     0 �HZ��qB����X�ĉ�U�냧���~���P:�b������4�3�Ѳ�~GV,�\6������S�M� C�n   @�!p� :j=�LA����>uT�ʋ�+�?x����
w���0����̾Q.�M��"��oU�*�\�i�����      y�;�ֽ��i�2qx�6��)��v�wV���s�����j�E�i�Vm{�i嚢��tʗ�,3P��� �-   ���I;<z<e��}L���p�<=��m���]����go@:��T��Q{���\��м������ӷ�;+{_N    �V���*��*�0e�����?�U�`'�w�g]_j��ے���åU��ɮV���@���^�{�Ա�{�[:������Pןy����J��}�E-KY�45��?�7~�S�{}��]��������l�    R �|Pf4���	@.!pǠ�1}���ʒ�^�}��S�lӎ�?�h��$;mWN�◴�W�ԮW^Q�*9R'�����F/    ����e�����#i�a�N��M�����c�z��J�h<�+�;>�����T<f�6�_���Y���/~I��re;z�    �fȖ/�}�����\�t pǐ�0qt��MQ�t�����04��kT4z����[��ڔƞ}�f�SY9@j_,w�(N&!mx�  �������I%�@Rܑ�lx+p:�D����.0��*�<Y��+ܸA�*XV�ٟ��F�?U     ��p���E�;�w$mݎ}���+z���
��c[m�ҡ)UeaP��x�h-�ֿk�%Z��;��W&��4���',-U���P    �?�W��#d 9�Hڪm��)�5Fb9��Cc�:K�'����ޫ�O?u��,;�ڧ~���s�rm7     ^����F#�!pǀ�V�]�����q�@q�f}��tɥ����ڞ�����|�T�\y�F�|�r�->L     ��fk�;��@2�1 �A�����/�S�j�Ĕ�
G���D5W\���=�mO=��=��� PR�Q���1g��V��N���#  �ňdg�;����c@>0��M���aڼ�2Qc��EE�t�%�Դ}�j�x]{W�Ё��r�u�ܹy�~2�����L�}j���U    ���֖2T��ɿCr�ܩ��Esj��gWz������W.�d[+�۩|T2n�;M��r��Lû�y�N5mۦ�;Բw��maţY�H�z��B�ʇ���ZţF�l�d��LQib[N��|v��1����fينb����UM��LӔ�4���ϐ��-��U� q{�ʍ�e�z    �/QV�܁d�#i!�O'N��_<g���{�0T
x�-�ϧ|(.V՜9�ԟx8,3p�a]��*�,-��� �K �'���  �ɈG���p�C����=�m��8a�H�(+�ކ�ؙ�����8�y���y    �Όgg+\��H
�;�6����i��Y'j���=�qv��}�"kj���ھ��{��6*������C���s	�|ľ  ����p��w$mxIQ��?s����m��<�T3M�ĝwx�!���    ��cZqe%���#pGҊ�C�n��	����+��މ�_    x#[[���H�;�����=�����- �
�U�`��  �Y[��g; �HHZ�׳�w���>��Y��Ñ^��������ieg?4d���B    �#K�k�b
 )�H��w��=n�:���)1d*��BW^$ �W!M8&  �-[{��|��A�����4�o+Ƚ�eg��2T]8����!�    88<r�;�ֽ"�%��-[,θ�C�q^O     eknaS�$��I3{�;��mٜ.�gl�' �`e��$  @Je�g$� 9�Hگ�]���vh��*���n����.�[��P���|4    8g�9� W�#i�[�����l�'�Mxd� �z  z�S\K�.w�������inI�     ��K��F��AUV�ڦVŬޗ@9�ls�Tk|E��hЪ����Ԧ_,�����`s�����~��:-dJC�v�y    ����a�'4��E�����&|��^��q���^��Vw�{h�&}����;��m�f��Ϟ<ǋkF�S��]u��� 0H�  �
w ��c@���T}�����X�g�>�(=p�U*
�d�9StӢ������9�|� /�k�     /Y&���ܑ���%�����N�Z���1��������N�;�$ݺt��44+�
��q�ڢ �   ���pr�;����*�oS���]�63���E�(*���}T^X�a%�nÂ���'_K��,���o4�c    �K�An�2w$mn������|j�\�7}|�ex����WKL����bwwd���     o�>r ��#ie���юv2S����/]�c�w��W�@�����+�ᕫtù��q#��<���4G� e   z���m�Hځ����Ѹ���ԯ?rQ������Kj�m�9#�ܯ[��m��/�i(n���
wx%�    �����6w$m��}���r��-K?���:e���<��V=�n����	%M.hL�0��p,=��	�ᕈE� CC�;  ��,q���G�^�Y߽�,�J}TY�>:V����1��_�~�Y~{�>\S�/�2۝��})�nw�i)oD��     o��F�M1�w$mہF���}��9}>~[�[�t}��uљUho9����iy�!�!�1�     o��� �.w��\�i�:c������7���Ǽ�Fׅ�&��W��o^z+-ϑ�2�
� 04�8	  p�����e���HTW�����?K�gOV�gj�������������=YQ+����A_��j�����/�Zʼ�v�44��{��qll�|���J�
��q#�k��j�}�}�
w    �ײ�����c�b���}u�;�Ϟ[��{�sj
G�N�,�p�������wɊ+�����9y��Ϝ�k/^�y3�*S�Z� ��b2���]}�t��VIol�+     �*���e�H��w�?&�7�M����|'��v�m+���9�������Su��4e��WT���J�e�*-+QIQ�[o��[�L�$�V(dGn[t���dLiA�mt�����e�o��2w    �'܁�F���s��
��Amk,�x]A�"1ى��xL�榎�QM����I�HX�p���� <��ikm�o��w��@�y�J{�0�w�z�e�u��í:@�}w�t�N��wO�$~fEU*,)9�2�=g�����u�et{N�߯ʑ�����2�>���?Pa��U
����g�zZc�K Zs  �"pr�;Ң���8��5Ž��{g� �*tRri��4��Ж�r�g}��h�-���o��sN�����ݣ���Ӹa�=�M�    ���;c6�	@."p�����'��yGiބQ�3f��+QA���e���O��7�@H���a]{˃��'.Ӥ���cˋ    �l��A�Ѱ �wل�2]z\�.�S��F��w�'O/'lG�[��Nt��Z���i���3�
w ��   ���q'pr�;eڈ
���i���?���˯ܶG���k�����w/�r'�ij|E)W�    <S;m��XĽo�����9��N�{'���(c��@��j: ��#iN��2ӭ�uZ�$�%Սw>�h��mb��w�� 0��D�-Ŷnh������������&��T"a�m͉��cj���(�����m���R-�VFQ�  ���b����CWs;m�/;~�Ψ������紹�ca`0ܑ4'h��KN�������e=��oK�q�A   Y�0eV�P�s�+���#/uU#�������|�R2

�݆��bQ���HV\v����$0�D]|��@P  �	c���g�q����mvƏ���w$����K�n{�!=��˚0z�~p���?�n���t�   �lg�U���O)��-�>}���>�s*л�w��`�*<�r��/'�  ן:�G��>�R�L����* C���5�E�}̲mىi�i]��Q��]O�� 2���˴�)ٶe���$��i��-۟\լ姺�)0m���f(�Ƌj[����c���[��s�/�� ` ����|̜H��;������%g����B]�輮yš�.�;U�y�  ���j�  C��k�_�м߿[vsC{e�w�/�í�rv<&E#Ð*<�2��|�&�W9R  Ɣ������	0p�H�ۻ�t粵���ɪ,*��؈�J}`�^���ʳ�q���q�   ��c�-9  YfTY����}rwڈ
���j
��1��ܑ�=��统��4t��1�tΔ�T��������߽O�~~�[     d�1�%G{��(D��;,n�Z�i�;}�/h�J]<k�[�~���N�OE���i�/���z     ���r�w�wٺ�u���gWhBe����i�h���#Ǽ	���Sg�_]#       �A6�;<�����ə
~-�<FgM�3���7�w�}�]�ml       �w�L[4�g�ou'�S�^�%       7�~"m�A6h      @�"pGR����2C�=�;���\��%��6�#jh�@K�����6m?���       r�;��T�l�q:al������{l�~��r      @�!pGҾ|�sz���Q�gh='hn�6}�W����      �\D���-۲[7���~{�b�L��e�bq�6�hsm�6�;�U;��u[��@�        ��c@������k/Pq(�5OC����g����	       ��;��76��t�G/���G��F��O^�xl�����nh       �w��}u����O���\v�����>q�.�=Y�x�uwp�H<.       ��4g0�-m�B��`@s�V����Jw       y���R
��W��V�w���z}������       ���6sT�n��M������Ϯ�O�Y�p�62       ��;��#t���Ұ�P׼�e������g������ض������5��m{       ���I;n�p=p��UV�1�o���is���]����zR       ��ܑ��ߧ�|��^a�@�       �\E����3\/nڮ׶�Ra�����~�u|}�0}W}�        W�#)+��q'       @��       � �;         p       ��        x��        �       �w        <@�       ��       � �;         p       ��        x��        �       �w        <@�       ��       � �;         p       ��        x��        �       �w        <@�    iP�o�B���}_,�����zF<&ò��&�-3�#\>Ru�N  @'w    H��*ݵA��?   ���    ��RG�H�"  �G� @J8���J�O�/�?r�ο3��5����w��?&Ӷ$�6���j�B���lw  �\��G�  ��)ڿ]��<{�el�_���=߶e��}��X��c���P���Sٌ�ۗsv��X�헜�]�ϖo�XÈ�@~1�  r�;  �IU��ʅ�5��PZ��<���a���ew ���_,����m�F�u X�����B����)  z"p  C�k��y��w}����Iʽ��|�%��g(p�=�  r�;  ���ԙS���w��i���״���'��~�qB�;T��
� �a� ����(uC��C��9'�K�7=�f��ʴIh�|DK  ��G�  mJuE��/�5IcGT=YF{�n���G'�   r�;  �Q�E����ڴ�^k$n��3h�ӫ��mTN��M��L{�v�	����s��   �!p  �v�ko�S_��)�@P�hX�,���@�$�@>��  @�#p  )�w����RH���K�9��9  8�;  H'p5�	N�v��� ��;  @��	� @����v�̮f���'��   9��  ��S���U�nЃ �O�l�A�N @O�   e��"���T����'�   r�;  H��{�[�F��)*�s�S  pw  �2����!j��,  @�#p  )������&l��   �� ���M�⁐|�6A�zɐ�y��n   ���  ���ǝ���$A�;��h)  ��� @J�C�RS��`tD�$�@~�-!��;  �#p  )�T� g �����R�-�^��;  H�X�P�@��5ZK�b6 ��MS?��\}�����آ�_}[�z�h��"�v�   �,HPG�N��3�x ���/��s�*+֗/���U냿�� �A�  R����݀<Š� ���W���9���3�� t"p  )��v�A�;����"N� �ĩn/��z�o
G �� @j����ũn%t�� ��&W��ړg��ؚ]� �8  )E���Pg}+�&��VR9�_k�2lKF��e��m���bXq�X�yf�kÊ���X�}܈Gۿ�w~�<U�0��~�_�~�.^x�B�CWq�޹O Љ�  ��i
�(n��,�U�k�i��c�N|��ў�ʭ���ŉ�lZ�%�C���UX3[��i�Q3V˷� t"p  )E5wo�L  �l^��òSX��	�vm׏�Z�k� �;w  �R�Q��	�mQ�
 ���y�:��p8� ��  ��e	�:O>P� @f3��WU��brR@?� @JQ�~H�O�� r��e�����#�* �!p  �e�w�Hfl  2Vd�r�6I���# p�w  �41��  2Kt�J�b��#1l˝l�33 z"p  �E�n�M���  #�ш��7J��S�n����� @J�ýS���A�;  �(�w���I1�� �p�   �8`mg�H r�q9Ǫ���� 	� �B�  R�
�F�O���� ��3n@V����d
�`�:@� @jq�ڡ{K!KL>L_]�@���|r���  wٱX�=ެqt���F�  R��@�ŉ��S
���p�&U��__:�F���A=�a�  9��Eo�8:*���  ��a�qR��]��?�+lw�MS߾����� �U���t�A2���  ����C�rG�Y�����7cde��~� �r�[$�AS��  ���'�u6?�,qҸ������5 �i�I#y�% �@�  ���٤�0��������aݼ�M��e  p���;  H-ʁ�u+l7��d��ߧ_�����_�u{��ݝ
Ǹl@O��9˶x��ѱ �w  �4h��M;�l���E_�� 䙮�(� ��!p  H�Ca;��  d8�c��H��@�  ��p�v۽C �� Y�?Z$��	��� @jq��? ���sg�1� ��   l�=��8 ��g�$p~@_�  ��= 3�޳�جx��k{ͷ���I�7�m[�)ۗK�@PMՓ �U���u��qd  ��lu�p�ƃ���*۵A�.ZXF� ���8�Hm� ��  ���v��s0����J��
  ��� �F�  �N^�yH��y;�Mڙ� �'#sNg�7��-�@a	��� ��‵��J&{{�S���pw���6 �-e���e��   ���`t�|��c3N�t�eX1پ�  @������ @�ضbj��J�����3��2]��2qwB9��j���;;�j�N ��  ��]�[�A���V��Q��W�  ���xH� �� �ԩۭX<.8���j����f]L^� :��.�]@rx� ��  ��}�V�hDhg[�;�fY͈��`����h)�{��b@8��7w  �"���F�V\��/#�Ou��t����PvrM �8�^  �;  H	;�&Y�7b��y��y{GwK���CӶ�s���% ������#)�XD �� @jĢ]w���aO���V^��}�8uB �]ox6�|H���@o�   %��L����G��
���6n��}���b�� Q��{�r�H�  }��  ��q�mJ��ƀ�[��X6�<h)Ӆ
w �e$�H�m�z��;  H	�[�_���s�j7p7�'1:�& �9o�� �v� ��}G{   +��u1v��hY�-;W�PV��;<�
w �]�=�-��Hm� �f� �����cq���勆叶)ٶ���j��������`��=�; ��  }!p  ��3]jmj�Vw�)�,�/P �x���0H,�b�ţ
��2����:�<bu��X�{{Ӷd�c*˲w&���w�m����wZ�3�L�8v��ٓ@�!
�M�`�--���Zh)t�=h���&찲�N��L�I'��mͻ���-k��%���I��I�N���=�{X�"�l춍lV+	6Y�f�Y�d5�f� sk3e����@�Cw �x���X^ �w   P	��[LNc�)�V�I�;�R��҈KM'J�".=K��$�c��h1���@Bk���]�QX��1���.�l$����)$�U v�b�204q�;('z>R�� ��:   p   �p��r)Ng Qo b�t��'Kדb&X����I�[(�����NS ❈����: %�  @5\٘��1-�`i� ��;@�:��ay �   �'�N�B^
 �P"�� (@�    �����]C��������{��u P��]e���e�(^#�{�q�^R{��gJ>�J��IӦ��u�|�s�T   �>��5��wX| b�v  ��]e� L�8�w�C�1�_nQ�_���Emk���)��%    ���  	 �;  DD�2^"F�qN����[kZ�^1�m�Z�NX-f�I��b2K��zn[�J+D�.���   ����C5 ���*"p ������DQ�P��՟���ѿ~|��y�C�M'   �D�� ��l�Y��� ������8�ӈq��P{�l2�    w���׽�.
�  �A�2Q�:D�j����)RA����l6��8텺<   H"2 ��A����=��5  (A�2VRƵc���4�ˋ͌�ܹs����<�j����F�J    �{�  qA;�� p��]e<��}I�Vw���\X6�    �� ��   �w�)���� ��PwR�H����     ��� ��W�C��; �"�*c��kH-�a�wÙ����j7��"�D��O��ECJߦ�hE����$R��M��y�&l�d���V#o6�#���6��1�m��$���gE�dxK^���N�qε�  �&���  pe㎈�<  �C�2�s��8l�N�P�io.& A����$�Ә	  C���Xz �]��:���
���| T#"pW_�����`�َ���4���� � �`�   ���,QJ� ��4M�V�� B��h���+�]���� ;�z!PXv �vס�� ��*�y^��[,jnn��5���A�;��|��6��㥿�5%%�0A�H突㸈�4��koo/�Z�y��ٶIC���m�j�mҥ�`0ؤ�4��٥^��3����CX��Ɇ���S���ٽs氍    j8>  B�2Q�q��DuuuOt:]CQQ�D E������������=�%�  Y(���2���G�T��"  %nT�q�&J�X,�< ��z���*��	t>�:�@  Y�!P"�<����5�� @�����p� B�t�" n�z��.��t礋�@��q\ @D�M  ��6 (@�>%i糞�8� 
�Zm2�����D��hR  "�O��;5Q  �v=*Z��p� (@�2���Die�ٚQ^@��Y�u��|��I @D�ع� aɉCX�-|�  (��*S�45^Ik�"���~�9���  DR��� Q_S  w����K�C�&�ɪ�� �I�L��[C��K��!�  ��C/�p�� l�SX�-���X���*�%�RR�j� x����ZmЉ�F�iE� A<O }�� V$��;  ��������b� xd0��Zmj���y��   bD�; ��'I�?"w�V ��������l:H�gz��S���v>Z���d2     �%1��!XXN �w�q\�4��X,� �t:�tt�����h� ��h�A�ٸ��   \!pW_��Z��~�<NE� =�9���m}���=N�������|)�E_J���P�	�}�&�33*�a��Xr�$Mo��)��ǘ�r��A�O����������z�Ҵl�X,��`��[6�R+�K��#���&  Dj�C f�  �.� ^`� 
��/a��X'�uuu_HW��u-+�#Z�z�t�:�d�)ǱЖ�,ev?T�=8Bky�;&������Z��Zo�Xڤ�Sl�4dHߕ,�;�/M��=xRO  1"��!����:    �՗P�`&��B����D�g��l6��N�*��  �,�3 ,5 1��a;��a   �*Ei�,�vʤ����N(�"�Պ�R ��u (���>�7bo�N >a� 
����yNL�0�q ��֐�^O��
 @4�b�K�(��   H�՗P��Y'�<:Pd�Z��  �() vX�4m��p0 �!pW�(���Y Y,�>`[d���  �P��;D��7 @��k 
��/���D��x��K	����| @K��;�2�
����]�p�6�S@w�%��$� @�~�l��`w��M�{ ?�0�2 �����sX׃o� %�U�6.�N;�V	�g,p���t�Χw�.�V/  �%e Xj����/���/X ��*�y�k+[% � �  1M���b
�c]~��  pW_��Jk <��<\�%�= ��Dۤ�u}!��)|��{[�CI�J� ��*K����ߋ� /BԱ�}��#[x  a�/BD������*�C@w p��]}	��) oX�����9ԓ �0��! ��� �k  P�pT}�vX���Y;��  � Ċ�2rw�^�f %G՗P<A�2����ɱ�E4e�T��Y�OA�s�F�hIT�	*����x��Z�������z�:�{n�G�R�M��j �/A�b��-�]a�#�V/_�m��y=��L8iS��Z(ڈ�kC��y�&�PZ�K�8�l�|�]���*���? (�^2�Z�Ͷ�q�����)�E�(��!_>��Z���f
�5��2O�S聧�޿����J�F�Wr��TiH�2���{灂�Q��)�d%A/ڋ
A?��U��38=Fp�E�^Z�wzy��^+ͫk>lǸ�h#KG;i����M �@��mDvp:2JWL6�L+YLF�;�ue�5� Qo�]B�؃x��J�m��#���;5�o8��ށ�F>�A�z@�O��~��L�W�z�� P��]e,DM�#��ߛg�X�"����Y�Q��vH��MZӥ�D�D[  �c<:Mrñք��}NG�m!y�:����ϐ�h%%-��ȐB  �@��5��:�u�Ld�h'sk�Z�l6�Ǥ\v	�$u�gj���N�o�b2��{;Z}?X���%w��?� �t��A�e�v� @	w��<ϡ*�Y� ����f������h4�㬕�4�i���m�%
]��h2�u��N�E��|�7��!�\:?�
�V$�Cdm�#��Eyb���W�~�T���3r(������z��鴃GP�����O�Ğ��|�,' � ��ʤ2��!-�EV���綴yD�՞�y>_�>�@m�o���Hx�	Z�G�����bCԁ�k��!��=A��t��gOʗb[�!�4���-#O��B����K���d��EBs��N�����n�8i�4��C�\�T����P��W��(�����]�y��F������M�R�0U���p�� ��p�#�8��g� D9���J:*i�K(Y  �4��w�!p�� B),�V�A��d��{腨�}�¡�{T�D��4^��A+��K:(�  	��
P9�);6���; �C�>�ktV�u�4�V�u:�tu"AH���T�RU�݀(¡�L����i'Y;lA�`����  �������C���k���ȡ��*AƙL&�����,�C֑r��pܥU�(���ECi+���M ��w��K��]4��D��4���J&+NZ�
݁;w���� � �; �$�x��H�f�N�+�F H����΃� ��&�q��4`$A�(*c�����Ki鸡���G���K���?�SM� ����.�p� ju �
��ʤi�Aܰ�lSA��j��4�Li�.��;lŖ�����(�NS#O�x�`��Z�C�>����80�~~���� �ŧeʗ��6] �B�2���x#-�)�e��j=���-�X�bW��!-)�sD`Q%e� ��]-w;�� ��o���#��3@4���?XCA��2 �������(��&�ɢ��Xk������q]�������p'B�E�EZ�Cx`����Rin��}FΒ��~�DZq(�>:��? (A� �б��6��u�ʚ��x��P���7x�p�&h�y�U���v��C��+�{���̱n��nF�v���ђn�p���lZ (A�>�B�c���L�s�a�ts�G�h�.�¡�;��'���{ĉ�9VJ����,�����5��L��4��s- �A?r
�����M�� �!p��E1�h4����5<��!P��ݱ�L/d�ظ�Tΐ̦��1�"�C���Cw|�`��E�ݰ����R��>����*��m� �AW>���:"sxbMN#  w�a���l6���t�5���@E}�u�SzG��;��Wۚ�s�:�<�-5g8A�a�q"!pWJ��BwA�NU�������C E8���t�����5	�; (�@�Y,���(��j�Τq��=ץ����GbaF[CᘶyMU}Fa�ɼ�Qf��A� ��4-�U�#��8�[ �;�_��h� �Z�3EQܢ��X�`I!��{�P�	���M�*��ړ��	C$y����p�C� �8�z��bH%  h� ��lS���:�n�t�eB�&�bJ��FC^i>Bb9�pW���ݎG� ���GP{���	D�46��}��'(����)���l~hY�H�5$:���sP��m�3��V�$g �����)$4��6I�ج���%�9�k��̞<�{M��}���HC�&,�=��  ��2��D   }��K}�;��g��.�8n�V��I(Q��!p�8�!p+��#5�U��I/�f!      %�Շ�S �k���8n�F��G0�=�p�-��^�E��w<���]E()c�A�      pW�N�Y,��<ϯ�8n&A@DQ4:ޖ�K�E�E��A�pB q�Մ�gE�     �����8���q&�i��`8 }7F���>q*%�+p'�a�
>Q ��j8��gǣ�;     x�� ��`6�3C�t=�; grN)�F��y$d���&���zD��'�      e�U&�,p!�b��b٪��J7��m�\����?vz���I�#��=��:�R�.�gŦI��<zizE	��i4��h��.�>�[�����n�w�%Z��cL���$�.�ԑ7V@a��=�D,����     �w��<ϡ��;��6ET�(��9%�ǹ,p|����ݖ�Վ�u���]��>���D2�P�]=�o;��     ��*Cw %�N!��������V�##�;����     ��  ��5@����{X��j䡤�zD��gg5�     ��  1D�4�G�z�p+���2����^�L    ���H�ӈ�\��C�iɔ�l��1�F3��6�mi�c��h}�jj���o�*�8.�?~ ��`�	N���uL��'�y���$b�q�Ճ�[&�2��     fxAM/-�C�i�*�����:M���Zw�}Yu��m�h��  ��v���mbADI�ppR�j��J)�d%q�@�̘U ��     ����t��
iFC�g5��d]6�T�}���ƎC���*�mn�HC�>4��X�k�sg%_�qE �*��H�o�����r�n����Î�YR3ɒ�IVC�\��6]�����k��l��c�,����J��6k��9�D����-FҘ:Ik�$��C�Ե7����4�}}��o ��A     ��q����i��r��T�*�G���G?^<���UE\�=���� �WP��(�����y��y2��'݀xgNΠ��Pr�Y�=��m���FK�9�d��#SF?2������F!�$�&ӕ��XL��h&CG�Z���(M�u�=̩Y�P:�:�$     ���z6�*+�s�4<�0i8}e�pZ����uTs����; @x�Ɋ�h_os�3p'�H�j\C���*�S�����G(�d%��s�=o0�g�G�Mg [f��
��q$���������}t�
    ����OO�;��!M�J~���׌+��#ӟW���NF���%v��b� %{�`��;&�Zs�t�bY�AW0�J��@eX�C��b[��C<�*��%     �9���^B���tZ����t��r���r��p@� [k�����!Jj�0��v��^M�c�u�g�D(3��p     ��Z��p�E��œ��+��9��w�B?�p=�s�n՟�; @l���O�ރ'*g;_<R�߿R;�Z�IKz�      ���u�ܭ���)�����9r��{k%Yl�jυ�]}H_ �Q����u߿�s�x�(��e����&� ���8>      �:��%ӫw]I�K
(V�2u$e����Lm&3��; @l�[�N2�p�;B      -X���=˨"?�b͂�z�kW�u�~�:U�L����� �8�j� ��cI�]�a�7      �]z��޸���{�RL��u%����d��]��/� �H�`3Y{��<�����{���; ı{L��ǖ�^��g���m�����p�4y%*�9��;����T�� <X�BsÎ�v���6�5��鲑����):�<E��^ڿ	n��m�7M��ާv�E՚ᡲ�����6x�F'�F�r�4~@źyC�_�����ʧ!�/��  b��tY;$���rQd��Ǵ����u��[ܦa-�Z��ԏ%V�,/[��/5�"���O];�  1�������BZ�>r�4 �F?�p�����W͢Ye�/��8�v֜����y"pW+!��# �Ï���1|81���A �3�`��ǈ��f\�|��}ʭw<t�|��u��_/�J�s��Ek�hf����?p ��������a� @��}�l|}c�8�7�^5�v�:GW�w  �8IDAT��	��"��  �Ǳ6$�!p�4N�������QO�����B���DC�S�������!3ɪ��r����8�LHh�1����@����Og�џ��O�H+���a!����dA'���R ��=\�05Z��'FM�x�� ��谪<����������Np��(A�*I�M���2����L\E 	�h��U��ێ:}�j÷�y0���
����[;<��ۥ�(͠�xU�/�~�h*��A�+:���� `�S��N��k]��� �����'��z[��o>M�#�vC27-��dx������ҳ��5A�9i���g���?��
2R#�2�PcO�y:��J-&3e''Ѡ�L�?��)V��@Jʴ�ʹ�l=�CY�2�8Z��/4��׌$奥�آ|���P0Ymt���~�[f��r���.p1��b��Z<c�d.UJ���y�m��A��; @�b}D�1A!�8^@w�.���#p�IO����,d0w�Q�B�h��A����4��/@$��(]��r��������Pnr�dePiN�ɦ%#�ihn��ϳ��4�a�V���qj5�|*���׌JϛF2�^����������MI��߽���>���9�c�H��e���eZu���|X��5��בA��߾{�x�����oU��^���2l����D���wtA�WZBˤ�"�A2,]��X�n���~Gz_o{�}�:����RE�liȥ�����޽SYE_{�#��z����n��Y�P�yg�����v��B׍N/�x���;��NE���t���]���y�H����?��hً�٥l��C�?�^F�p^z�Z���ܳ_�]%�t�`�`�SZ֯U��rf�H�7��/WSMs3�n
�2�i�i���)4e`!��{���}�n����\�����۟T������t����o�,/�J�t�s�n�:;P�>�����o�� 6�u��.�N��}_~�h*}���͇@U� ��/	 j�;��{X�(gyZ�@��P���9U��"9�^I��B����jI�f&�o�C��W���&��?_��-@tĂ����1��s���mm�l�I�o��'ϣ�gLt����'I�s��5����[2Z�3��e ?N�l�4:ݾ�r;� �=-�v՞�߫{�J_�:�]8�rR�}�#�;m���ەU��,�fÚc'�����=k��Ǜ�e�����O���_�B�>�=p}�?����G�"6i��u9|i�~���=�i|/;�s���VW�����=���?���%4:-�p�ay��b�p����왽��鞷?��է�N���4�����;�B�|{�ߤt��_�Gi��i9�ъ5���K�c���� 6�1}4�rfc�Y6~(=��6�_��<� ��p�bZWGZ�C4<�=���fH&������Y#�l��b������44ӊ;�ɭ�\��l�o�'U���/k1����L�~4��}����w���sJ�h��Y4�d�C��T�P`*��q'������w+���t�p�	"����vy�o���eꅝ{|�޼����=cMP�v������~g_����A�5�khay`gI�������^���5�\�n/�狴��);��/��^|�Z�}+��Z��-̣P�o�`i�p@�m�3_w�4�\�v�M�M���c�5���ނI�H�٧�Ι@���y��@� ���<���N!���к:��@�y8���;�K� ��N�)Yd�(Z����ƀ{��� "�S���O��U�j�W�6�/�p���+7�)lw���V��AE4oH�}+������tJ��j%�KG�J��;����%����{�
k�}��ʻo�:�k��X�t��-��6����^��o?u���=Oc
��z���J��7��g��Mv�h�ѓ^�yw�������o~H�s:XWO���1�r�2���76ӵ/�P��i�8m���������x%m��-n��6�������E���R~�nKǕ�Cﮡ� �A�2�j, ��?%eDV�
M������e} �8nNTHO]7�m�C���Dk��������5F]��uU5��7W@��o�D�vT�Qy�ު�R,c���v��fN�̤ރbG�豕���QRLW/'�FC�T���ܦa��ϿXG��|�>nP�rmwG����?����z*�۲T���t��D��{�V+����_��N��ށ!k�;����J�Ւ�䯻�N�|��+Ϟ�=�ut�B�ǰsձ�����VR�q~���g�V�~����Z��K;�ғ�-���<ZM<J�/soS83���Ň�|\�ȸzg�a��UG���|�\f�;H�xX9]>��rS��LK��}�<}�����õ�h��'����=��Ҕ�B2H�3�o�>-w��cƠb
�?]���/�ȝ�����3ͭ��f�N[{�3v���[Է���kj��׎v^7((��Ō;���D��,�zl��� �; @�Eߛ)((^<ZWG���k!z��ϒo&/�Gl�������H�����NsE�ɂ��4���lx��|����-r���y���I�v�P��l�A����k�~���胳��C+Vѓk6�M��l�4��˩���ۤ�+6l ��F�|���{���?�2��qEy���;(�&,�;'���n2��{�'+V*��ys�!�{l�u���a��G�������K�{l��ϳ=�ᗴ��ԩ.�b��c>,L��ts+m?}�&+��QێS���!��tvi	-���q�ΘL7��-��GG��{}�~����CGh��5�~y�et���;s��m=y���9+���r��a��'���y��i;��;w��y��*�jD�S�-��譅;v`�����:8�N|cղqC� $���g�`s%\X�v�p�<�p�h#��	PR�:za���!6y�N:v�Ȃ�������~U�]���l�/�P�$��+����_2�V>.w��ڈ>>t��1�+�f5��_W�����c��)�N�^{�9�~����t#�[�,��Os.)�ԯ�9ȳi<���%%������S���cIW���>���cm~n���Q��}��>��J��U���������m����c��}ܮbgc}RuܯiYY�H��T?�t��8v������5pg��<�6��*����'(����~���Չ�ъ�}w�޲����h���SF�lFY��MH3���j T����G�h��wl$㹷H7j
�'�",�X��F�gf�A�p����3������q���TI���jH�-�!��<thP��9��b���\�b(:��?M��2���xp�T������p�to����q�E����һ��ſ���=pw��0'9٭�W�I�j�{
��1��Qo�Q�D�������%�x�zp�4�ͪ���	��ޮ<T���쳵t���A^�u*���V��#'�:
e�-�v�R��C׼�&���������%�)ܔZ�33P?R����54f-����;��߽R��]��y?����C�(ݡ��b=�4n8�tu,��#*�	�L�,Y���%�����+���Z �r��Ow��a�����f6�h2�y�Z���v���g7����6��Y)I�#�)iH����K�4����M�a��uK�Ք��C��iK*U߻+�]��3���s��W+��wזڻk{K=��J�����@�������V�/�'�K\ ��ng�Z���[<�|��iT_���u~�o���g�,��[��(#�޼�z��ye�iʟ�C�g{ϒx������R�s=韚B����X��~z�L�v_�$p�7������_��j�������_�@��7Ұ�9.���۪���E%��������*�7�;:�dS3��*���I�)Ӥ���w��,Xo����7�\�Q.�����=&��&̧D7cHw �x�������Oo���Ç�Eg(�h���z�w�8O�Y`]��.�bE�1���*��D�w< ���CKvO�r����O{(�4��sP�-=�$+�N\hq_�p;E��~)΁(��/��P�KX]��I+��+�!����)R��ʿ�z��C�SF��4^6$G��5߼���Tߞ�z}�����h���#c���Տ^_����������1#�����͟I�����~�����4�CKm%ϟA���s�q�Y���~�8*HOS|���
��������|�������~9N��Y_	?�;���Dc�bkk�Ipvr����OKqܙ��N{�ǥDT�y��ŋ��^D��x�Ӹ�m�Iߚ:^>�����ݤ�|��B$����yp���z z�t}�_w�uFѡ�5���  t�V���X�i�ɱ����ri��Z���P���?�s�ǰ�Q]w�⛵*�i��Z����wQ��K�ʁ��������{ǲ J�<�L��1pc�;+����khk���;�\>����b���?-�]�ɰ��ќR� �=F)p�T[٘���=�i�C=r�)�/>_O�Xz�bP�����St��� raz�d;��N�������_��T_��N�䧱Vun㛍�߃�m��d(����R.��w�y�ze�~�y�������ǫ��ۖIˑ�s�ؕ�v����+�����̱5* @�W(� �<��V@����u}TJ��陊Ӥ���3i��<�5���i��3����� �)�� ������=O�ٺ�ZL&�s�PU�^~"����jz�>�V��x����guc�AY��to�Ǿl���	��~x��_�k������|�==��,���ӯ�\O�khÉj�R.k��
9����1��ݟ���;�gi59����g\�:b�߯�-K�.�M�>���o�E�Ϙ�x`�ӮŻ�o�e���b~��Z:�ҦxF�s�v?��� Z����q�
�5��p`��C?+Iʏe�+�sX'N��������d�d���[�~)-GW<�������P.)�e~��ܻ��dȥYL}��]}��%  ��qk�疈���uP����yW�J������%S�����_���@-l'Zc��Y��d��"Ǔ?��gӑ�(��?w�y���+u.�cda��c�pD�����`��@�S��v����]T�}?�`XwG��u�����ZH	k��ّj�y0��	�=yu��-���;�❯*��;H���#����췏5��6ol�]g�h|�u�Y�{IE)-($Ϳ�>�x���;�u���+�w���lk;t�/g-�������#V{����r�:,4�Mu�_�N9^����l�'V��?kGwLK�\%�E�NS/6���ЗG�τ�·_P����G���dt)�LE�mA@�R �Sf�k�N"VAa��=:X��^�n�ҕ��o�KO�o��6����jP۩��M����}��l]��Dy�
އ��Ѷj�Nx�4��k�߮�L�`Zi�3g�����v[��Mo�R���������B�1kaY	}�d�q9IʥcNy��n����~V��1���x� r�SN�X��Xk��G��t��2JkɻxX�ܪ#+�s�߮�w��14��wX�۷o�=�6������a�|�P����R|�����{��94�ȋN���X�G��N����N��^�_7l�_^:W����K�������SgƁ�T��W��N-����詯�j����ۦp�G,���M��KN��s�t�or�6ο�q!75��KNJ���*C�e 1{�˪����{��m�<�>�Rny��S�|�.k��T��/�v*d�Z~|��z\9=�Ӓ�;p��-�����i�/(��a-�{��l�q�U��![8�=c��y��V�O\3�>�w\�Sȁ��=ʵ��ݭFҿ�\�*�ka����ն�ѩf�V�Ƶ#��_wnAz�����}�۬#�����})�hQ*��J���ե�`jA���Ov����W�<���k�����è���V=��XV���f;�����ܙ>���YN��w^?wX,���J���<�j})�N֒~C�)�i֝8屬L��A9��eю549��દ�Yq|��k��\~��#'�mL�Y�)���%�.XH�FU�[��ݕ��g����I"	���/vז u����8}F�ͮ�D����cN�"N��shh�-_K�]:׾Su�|��� �Z���
�6�o^W�=�NG&�s����);�@w�K��l��<���lY}��)t�sR$��W�"�$��Eθ��S�_Է��S|�u*�ˢLuZ����>y@>-*DW�(s�{��f+�_u�s'ì����Ν��������;�^~{�����h�=g��"�O�L�a�	­F���_ٵ��c�9�rR�nn����(���dxc����a%eXi�R?�A8�M��ҹ�ၣ-��;�8�5t�X}��c��+=�����u���M��I��[\��O��5Ј|�М�w�޽|OfR�S����뮳�@��U�<����6{��@-jt���W�f���>�qh������{t�+�{�C� v!8�ű���-P�'Ol̄�M�S�"͜�M�xv�^���OO�)�
��+6��) ��H��VJ���(5IO��.�u��Y<z�b��Խ�3�l�t�"x�������]���殁��Q��˼4��̼�����/!��0����/�F��ȭU�dg�U�dLAy:לr���>�k�u�=��&�L�v����]�̕z�r���'���T��n��2�P���R�j�D���n@f�\nbl~zh�j�i��q�7m�[9%�^��۫g%a�m����*�ά)�_���Ȗ�Ǐ�Wv�#o\�R����VVF)p�i�r�2���-pgީ<H#�g�����a�Th�?mp�S��Q��XZ��W?�d���6�V��;����m�aҺ����v��6��{�c�'iC��E�f+�w�!p�Pr\���J9y{x�)$j�����c�aN�c��GNѥ}Sk[� �rl�%�ЙbZ�{М���(�u������MO�S�4mM�rG��0Jz�=�3�ûE�˗���[�����vg2�<ׅP�� �х3��1͓�n�׏*���&�˦���+/v�˕h�Y�Q��~��R�q��;��Q���I�yrؿ`H	�����4���O���R8��1�dmW��ùQ]{;=�n��4�/4�?6�fN�x������(X���]n�b�,zc���S��qy�ە���5�k�2K�.���*��]ZBo�v?K๭����Ӥ��ޘ��n��u�󹢻�~ �0~$�a�{�+�����~B[��4+��a�!@zDZ��"��\�i�^>[d���,}~ܻx����ꋇ�% D�>��n%�X�`-�-�	"Ü�_wGg���:����p��y�
���.Q�N���Hu�O�e�YE�������,�O�Ȃ�@^�c���{�� D�`K�|e���[�6����˭ܿ:n���ڞ���^�`�������t��!p�X��9��!=�������^��;�?f���'��k�$���Ӂs�I�{�Z���4�c�=�u��B�Q.?�j���t��1��y�n��������(�����fӝ���ӛw�����������T���C�h�~�4lY\��}k�x��Z�o�9C_y�=�^��\�T~��={�O��n<��D��r=�3}i5<m�����XE�Ϻo۳�cl>��:���v�♓Oo�I'�Z��,���x*'#��{=���,d�^{�Y�!W��^zG�ζG�]���������Yg�_�2���q��i��=���̔�m6��w�9�[ ��>�o��SRF�XϪؘ	���ɔ�x�퍤�h!��-�è/-�Ԥ�ޓ�8�wU��PjeDq~��)I.z6�Y��9�ΡzAF��w���޲=;� ���I���wfM���Ե�;�g����1y��}�:��}��3h�B�yfbQ�|��l��y{��ǵ��~��M�&����������,��F����������r��D�ʗ(�.��E�=�{����6lw�_6����S&������3��;L�zL44��Z�@��C��<N��,lv�VV�5p�xe�56˃?]4��n���=3'�_ֺ�q���k����̽��:"f�Tn�<��ݲ[�q�<J��ZT1�*�+7	U=�7���'N�?�V+��p����	$pg~<o:=����r��=�UKۤ��wGv�������ق�S��Ê B��y�^鹉�2QƘ�'�x�E�y�F�`���K��s�����>[��ک��1�[}i��S�y�Hڮ�f�͇�2/����|?�N��J��]nw�������pN��5���$h���M��v-�:]o��O!��4d���k�ͰNS{x:�<\�-][�����~�T�8ԡ�jB�	^_�`���:Z�D =��2��MW���^�ZFA	�]���K�,7K�~�:�=t�wit~י%%YT.=���
ӕ�`ۅ�(��<���<d-��x6}���ݦ����tߴ	T���w{{�X��B�� �e��<>�C�w��ھ�@P�*��������k��/o�=�8���_���rq� v��t����:�Յ��B���c��Ѧ�S���r���-D?��]O~%�{��j:ڠ���||��4(?>T�55!�p6��[�6���r��Q�~�����f�VZD���l�s���W�U� �\Z�����NS#M��-^�m� b���R�h%�C����z����=;U��y��H��ޝwג2E-�X�v�rͱŰc�w]�w�.��R���>\#k���v�:���kސ��ίЍ������D��K鶉�=N3(3Cq<�[��V�J�{�������[M�en<�pw/r�	��m��N7� ������]F�J)�f5�WTu?c� ꗪ�2�������V:&��):�gy�Kxh�4����n��z��ߪt�Y$���	[fY�¥��L��}G�-�!����T��>���t������_7NMO_���\��U��J_}�]��O_�KM�P�CP�>�[ͽ��޲���F����=�9�����\"pWw ���l�u��-P�9c��{ �լI�$k�S����I;�";SI�r�huNaBqV�S9�ܴd�ec�6cdw�Ù9Eݯ���`;!��-�kf�{Z��w�B���/��|+=u�|�e�Hy`������'h����Թ��;B�q������'Wo�o�C���ӱБ�l���Yr�oe)�=�dz,���_[��MW������A@��Xl]��+��g^s��;*遙Sht~?J�VS���Z�{��>��b��٩#�~�8]=������s.��~���45M-���Y��s��t���/:�����YII�o���NӅ��TO�9�O��_������l��է�c��l�������~=';K`�n�w*��n��'�(�ug������!�h�t��T_i�ȶpgX��ߟ=�~�n���p|P	"��=��ɘ�'�R ��[� J�u��ʳ�116e  ��&��3�J�,YF��zH�^��D�m�A܏/�!JX˿���5ǜ|�Ёt��o��[�f��j{~|��:�����k�K�0�o��Ye�t턮 ����������V8AU��U'#��C�\:t0���)˥#�T}��`!����c���Ɠ�i�:�m�ꤛ�c
��-|Y,YN�?��m�c�vfɈ2:����묣���מZ8�~����7��ҵ��R}�e�+����n����,k	���o+���X�H��/UA����r+��;G��*���l��)��q#��a1[=������߬>�`�ʠ��tz��ͯR&�OM�K���	X�O�����R�#�ˇ��}�X�{���p���6�8E'/4�}��fPv&�,�X���'-3\ؙ�L���{���L�i4�_�S��Pz��k�R����\%-Cm?�̶��Į��F�R<�����i�Ѓu�{���t^�{�Qa�ɺ�����X{Կ�\!pWw %�����,�!�� @��4jt�4<I�e��,y���0�'y�\;Q�����7_����]�Lr���S�֩#��d��U�{��-�["|�������t��Z��)(�·�����nH�:���I_�>�o�?�7�6�YI��o�![�y;@����q=���Z�ܔd�>�w���P(�ʤ���|Xɟ��P8���ۈ�CS)�u(��� ѯ��D������۫�m/n8����*c5�E��
 ��{��	J�  Dݓ�S(:�<Dr�2Tϭ���;k�7�m������M�kƖSa�{+�T���H�����[{�4}XyT���;@��=	 ��V:�Ё���g��C�2ADԦ�P��'���x���gb��}  �u���^�T�y���,m�J�4�wR�Z���8��^��~��:�00��*�I%4q`>���ڑ}�����ͣm�g�gޗ��  � Ăwv��g��D���~,w�!���q)#�GA�  ��z�V��sCs� Z����O���ny\NJM\@3�����4���}zV�v��B�<w   �7���Rms����ո|�����]e�� ��c�D�j���  ��4vi�����t��SFГ��Q�6.�Έ�^ �hU��s �Xc�W���-�L���=G�:������+3�	�'zQ����O��Z��Tç�   ��/-�f)�YeŴ`� �3    ��kwѽs�S�.q"d�l�_nf\�[��� BƱ�;��i�];�~�/�o�s	   ܰ�}Ɛ"�U6�fKð���3���"YW   @M��:�V�wNM�����hmC0����; ��(�������s$Z8n�J� k�&}
 Āۧ��y��m&Y���wג���C� 3�Jr2���H���~��,�5t ��O��M�$��i�z���8/�L%A�>��Fb�n��y�!t��Q4���4����Z����G��=Gh��3d��   �?|��n�4�R�:�wl��[��w���p �/��n1��x�5�|eJ���} @tSܟ�[�|Z�f��[�)�ͤǖͣ��J��:�Z{����z�������A�����]s�Ӱ�\���>�hp�̱4q`�����g�8_�9��?����ٖv�����)��*�GO]7��*�:�0L�w��'j嚦    ��TS+���m��˦S�{f��{�|��AI�	��2r. ���K��f������� ք�E�ٖ�r2��{�ɭ�%�utɨ!�p�B+=�n7��y��z��c���c�'L��FZ���"�u�ۥs�=G�g���y�"�~�0�����.���>�w���⑥��m�Q�V����Mm���#�|��Z}!;   $����I7NNC�gS�b�s_�9�BI��� �(��Ԟۂ $�|�� b�ʪ2Z���d�f$���Y�t��}��.�z�J�y�Ɋ��ֵFG�~�̱na����t��U��ESI��ȭ�{�m6���_UZ'rR���K���u�nD~r�4������p�|Z%}���Ѩ�"?���u�[���u~��<�:u���x���C�y9�/��R:2w��j7���-��Y;�k	  b���+����_Kz��궱���VRs�)$�B�>l�@Hp�����Z�����v� "p�����jy�E����Yc�E�]T��@O~�����#K��6-I�t��?{{5�<y�"mɸr���W�T��wLv���yj�v\f��o���w�C[��"�WWͲס_�4}q��>��N44 �6f@�>k<�1�t~/ێ����YN  �v���#��7��'O��-���C� ��t��)�w��� .�+@��j�*�u��i�?��I_�Gn�i��*�e��_ic��m��d��E��xT)���E�����r��hpŨ!��Z��=I���];�iܱ�f�������I_�9�~�t�<��1e�ٙ�j�װ���:��^��G߹t�|��_�  6�Kږ�2����J�bg�9���C:O��C� v�������q�wT��83����|�����4��}v�>z�mt��HѢ8;�iU�ږ�ߥ#&����O�YE/o��h1 ;�~��w��ES�47�~��M���39lg��>�Ǘ̖�I%rK���"�u���C�S�H��<�Oa;�j@� �f�=�~&7*Y8��b����?y�*cᚈ� � �%����cf�; ĉ�����K�Ғ1enk�UGN��ﭧg)��e�د7�w���z�i\7��w^YA�	�i������Z�=F��}s'8M���}��Do�fv�A��j��_��F-Q�y�oiI���l��ڥ�7����i�n[���;�j2I��t�=:��  ���;^�����R�00�bU}[']�w��=���i; ��Ea��=8�; �6�y�.�J���֢���=�����I�Vy齁�ڪ��쎍3:����i���65Z�8���מ���~�S'�����lrz,�p5ݡ�� �)-� _�����/: H@m&3-}�]z��+hfY1�v���y���oRe��U&H�w�G�S�W��fc-�y�V��]�ƥ�>F��,��9��cmA<��Z����b2�Zx�_-vay��Pt�}\wG�l���^z?XR��ƧHӺ��'��x[�H;@X@�b��kw^�V����y�m�ܦ}r)�h���m	��J��@OV�:���i�C��h��L=M+-���u�p�g�x�\R�4��?�J��:��MR�t�1���d%�5Z�N�?-���e˭��[ Q��۞9��4D�N��@  �x��m�k����q�"Z:.vj��m>�������~!pWY0��� [-K�(����\��V�)��M�~�F�Yk4Ӥ˩!|N�?�� bSY�Lz�Wр�޺�,\g!�QV�ݛ$�Z�SJ��z��>g��X�vV�a|w`��j��Pms�om�ڦ6:��!]�J�;hO�9�������=c�\҇�p�]>�~v��i؎�L��������>^�Lр�o~}	�(ȡ'>�B�X�����A���Tz�Y򎤦�/�7wVѷ_��:-VHdSJ�� $0V
��/��Cu�����ڷ��՞����g?���Մ�]}�<����� �&�(�^���p���ȼp�b����v�N�\0�,,�Z�0�f5u���MFi�.���MƐw�����SG���� G�����>R*�������壆ȟы�_�TJ�����+�*��s��__Uu2����'�̡I%]�>z�L�a�0��+ik�Yy�-�g��ճ���0�M����d������o��Ƀ�����sg  ?֘��O�������7_*7V�F�m?(o煣�w�!pP&�FV�5a���3^B��`�h4�'���@�yh�Y�:O/-����p�]��Gr'~����P�D�*�;o|IC�g˥U2���,l�ڋ+hg�9�ǰ`��_�}��Wl�h0up!}u��q�
��'�_G�o�'ܹ��~G�+ҷf��?��A ��*}��A7fRi�|�� ����i��^��_9�n�2����6;c��ﬢ���s"p��0��k�����լ�' ��B�;���`��+�o>@����,�aЅns;��o��}�~�l.-W!��+�Nү>�D�N�S|Li�Ly��u�z��>�5u�9k��xV���飝Ʊ�����Ϡ������/�3�m�{�x����]d�^��z��Ľ���#�U����D�0[i��:zm�> �����ae�^����Y:�����|����^Q�UT @t0�6�n��c'���k�;����81v��%�q���6Ŧ0�w�#��N]���}s�����wo�N��gЕ�����3�y�^�j��w������ơބw�A�V���	��ټ�n����ױ�]}q� �-tO��eO�A1�# <��!A�%<�Â 6,������̵r�p�|(�\.���@>�j�c���
��Z�6���D�OVï�lb�|ZZ�(,������>�i
���p���x 3��zv���'\]c"?w�:X�<{|�J	|p���1���i	���At�n��{v�k��v��AD� ��y}L�̈́_�����8'@C�W��d��Հw�!�� $X�֍�UlG�D�N'�K��M�8Y��S�TO.���1h-��AN�Uu8SR��Zbg�%���kU5�:>�y�DzL��%���Ǵ��YX;�vȈ�t���E�),�v����H܉N����~v�жV�?AD�폿=R�ҍ�Ra��^pk�l�Grr���>�����?Մw�A1��� �����j���y�������}1b"���|,ݍ�.s�l�~�v���76�u�lh���y���9A�;�R��Y�`�� 8��6P\Q_l?�����"� :'�N]`�WK`J^6���FwO����v'�V�M̽���ǂK,�� �]a�$D��f�m�X,ás�8�9�W����Rә�7A>JNb�0X���& ��A�k�R�װ�<��������G�����nI���򼰼
�3q��_A����n�!"DHA�UB۹VY��Ե0$_�-��u�V���^�A^r��� 7)r�Ĳq��Q!������"�0F��kePP,$����݉ZqW�	���M� ��f��X,���ī��h�A�Grt8�8e$L}}��O� }ϣ5τ��#L.�I�^��W{Aq�ӭ��KWA��]�O3F�o��|Y(���񔍗Vn��{g��}'��X�u<��oP�ټ7{l<u6�8�,��� �D*�#���ֱD�ƧH�����f[ =g*���=��>�2�a�0F�ê�@�ǌ~9 i4��y��"h�.���7H�R��DǱ��,K�a ��RPf�,�	��AbB��G�X��M��5��_��+�r�L$�Z��_��M�������NhJ؞9�'�:���j+��k[��!�?��?{\m���U.�U�����=��@wE�~�Ε4�Ε�X��
�Z�..���*xJh+����x��=v�=��!�����AF�EI#1�o��8uŔ�߂�S�d�-�3atNJ�EA��)��{O��N������S�Ze-�U��;�wÖS��WI��Ov���E���� ����b�N]�Y���/O��-`�q��K7i�M	 �Mڢ��+)��m	2�˼'Ϋ>.�L��<�i��ex�?a6�S���@��4���9H+A�7@���o��x�V����g��&k��#�ߛ=&}~�Z��On�}p� �86,�Ep�����q���_�"�ć��C{��lUm�OmǙ�l�AS����Nz|�T��O5�ٯ6���H��� #��ٕ��N�N^)��G���#��55��B��B5�^U�\����,ߕ�[|$||�D�M�i�X\`��ە�g�\��?����CGrS� ��qC$�E��V�#��r���je�?�u��oڒ�&^�\it�� ����a,�ǊJ�b��h�.?���8^�!�����/�n�m��.^�����(��F������fv]��Ie�WR��ࢩ��18���P�t��'�}��s�Y���i!��w��8��������b�&Y���!�m6��`<P��4�-�A�Pc�	�	�1CӁ ��@�	2`��>���;���5�;�8iX�>{]Flx�N����p�r1�I^Z"��:D�ذȿR�|/�`��٩�����u§��1�E��6��k��e�{(&|�� �Z����b�����\

=�5 J�k�����P>�?q��]�="��|�f�w����������
ɑm�m�-���|:L��r����HϤ8�������^�	�����L�������,��`@n/ (����]�x)�!A���;] ��w�-�}��E�t(Ŀt��u���k���-x`j����}�Zr/�A�7e�E����.cA��f�06Dn��qp�%����Ӹ�bw��q�0����NaHp'Bvl6�Q�łw��M-:<�����"3�t�� �����>$ק�`��M�E����� ��	.�W2q ���jFlt��fq�-��?<nx�sU�g�ڥ��\��-��EN�!E������
��p%��R��:J�_l�_�~2�7<;v0sK�ZM�#�'L�zfݱs��p>�9r��� ���0":�6]����KlA����=F��P"b{��&�k�M�O���Hl�2�s���-��"Cһ�� �c�p�|JU�Ǽ0i�Gk{G���?���SF}	j�?5�C���[*�-��?]���N�0VD2B�0.��B�z���C�[��˭�7��!�x�ㆰ�r��0v��@��a���Z,�n��p ��f�U�'��F���&L����E��R�E&�ʀ.A�k��?��ݢEQ�^Ϭ��� 1""���[����b6�E���fq߲쎿98�E������<�2�`J^6�}S���w.�����b�������P>|�퐦���M�ė8O��e��]�z����x��"8\X
��p��
��V�M�
��3`B��]tI3�wW��]-��!����pg[�d�9���5�;��c2c#a�����+�8"Z-�Օ�P��Z)���%�����S�sGq�g�8���"�,�g�������u�w����OP��*#����i$�-��w��}@w�r����5aL���2��N�lX���B*< �)d�8��3	� ���Y���Pӎ	AAq���RP��+r�T٪I��ǋJX��aA����M�B�=xO�(���@ϭ�/���}����2�Y�����7uOci��PQk����&�w'/)�E�<[Z	3>�5��&���0xw�H�1�a��Y)�
����v���^���b��s��ά����kK��Dw0���j�����.ʂ�����v�M�0���:3<��Z��H��u�X�{8RSp�Ӆ��&����Y~�Bt�3mhlر����gB��-��/������Y79_�:������k��	�
�>܁ ���l�j��G�]x�p'���Z�!�����I���	�C\Z.n��^b��iK?'5q'KW��B������=�]���;����d��"�ms��R";�&N��l�jy+�aW���S��YJ�
���0е�bנ�!��Ć�<�ǖ#͊�"gJ*�������������7���i�ܳ�]}��>r~��*�F��$�@���c>���7���W�E�ԕ��	�����Sl��oo���g�� �;�[tW$�g���fq���`��	t�6��2�qh=����8��(J_,�dJ/�V4�5�M�\DÔD�~���E��n��Rn�~��FVv��8/
�#�}��HpW�	��v����b1	��[�N'�z�n��1A~�M� a�FPq�<���֞�zD$<�Upw�`��w��Em�#}��`dv
���F���P`(����:3T��1��\�;5��G��5W^[Ǭ6��ԧ�_ ��9�%7�w���D���`fd�����4��}���!��W�+��D�gbd�=Y�J1�[�&�h�޵�������Zu��SpW������.69��j/熸�����x߅+,��q/<1z <;n0[����9S-J���T�؆B3����=pK�,����(*�E{�;�G��������_xn�P��� c[�%&�#����n/qQႩ��m�
�����w�4x��_C�p���q.�a��#����x��{�����|?��݊D���Q�o�v�O����f�m�Z����@���X;Y���z�d��QK���Z��X��d)(6�-�HBx�,����1��n)L��x�a���C��k�f�&�`��R�Ps��%���d���|�77�V���R�[�^��v�m�.������>`�SA�$W����{�W��9�w���mO�qY(�r��~��R�<�~tmw}������3Xq�!�ú�����-������i(��anaN������C��}jn���B׸&�g$²#癘��B�qL_x|d/�kj欮��wG����9�.���_ϖ��<w�W"(ZcL��'����&� מ��Wթ�[�ĕf..����sX��l-��N�5�{[�l^s�w��.]�����Ĭ�������������Ò�D.����9����}w���W*]�Ԯc�	�A��Ͷ�b��j@V�m����:g���w�Y&�8A���-�Z��0gD{�P[�����]�����~P�s@�D���롸��TT���q:xz�0(�����Zf%���vr9��t0mp.�'D�ղ*X�� Xl�/<�o6������Ȋݝ�e���`>,�
�j[v�%p!�_�پ��c\��Hpw{���ܼ�=���q�ŧs�1om��3�U�}WaE%K;/\�m�	���Gw�
y]@�`^W�;	?���v�?zfσ�v���h�����Vתj���c#rᧃ��������+p��ΛĠ��}TVL�M��`W1t�ū�6��wܷ�:�.h�3�d���T�פ;��`��+���4��R�����X_?2��"����p�~8u��G�#�לZ
�Z�޺k�ך���\>��Rf׹B�
h�>�/���y�����؞���qCX [\D��w��x��;!�t5��?��1����G%eJ�	�A���~�b��<?�� ��;Y���Y,�_��b;���i6�� j}����Of
�D����D<�0�����&�/��'�_�?	�� ���f�<�nK�q@�����?sS�����9�_)����.���c�uG��S�>)�v��SLd�y�Pu���g_.���9تc\.�w��������p��>�%�կ�t1⣝��7wqK ���dn�G�\�S�J	6{/��7?��Ά�]]C-�h��:�;|{0�V���N��]��� �Ji�:�o��u�Iy��yk|�����x~5n�� #s#��ihm�f�T��/���Ő���J�S��=��g6?K���V��}��m;��˞���w�|iL~�+X��4�T��*�����]�7�8���绎�|��ۖ.4�u���]?�68�D#�v�,����y<Vk�{p+��b����B%�Tk��o��0��<���
��c���V�E�/
�Y@ty-܁'w� ��d{�9��پN��t5���,&HM����@!�o��"G.U_�ƸZ"�u�}�K��N���b�'P�Yv�,Z�x1������!�����^9���
JLp�������`i��U@��\�	޺m��릚�~�ry%��V
��vnH�'��f�b��ݮ�?o��Vϗ���\��?>G��e]�
��l3ۑO���o�i1�c����&�i��-
��5#����Լ,���ŕ?2Ky���������ٓ���Z�LqE<��;x㾛�A���m���;��sF�C�m�w���â����4Ǯ�B�5�8j�Jh��1Jh�V�z�R��1P��^�]on�W*Zc���u~���Ůc�ǩ#!/9��1Zs)��1g���x���X?�A,�P�	�h��~�l6c��!B�Bs�v^�Y>A���U9_,� _-���`|p�$��\�]����J�s�e�Ait��@N]s��ŉ�ы�.�,~x�����s� V:{/����x�����("�z�H�jX	��I	,5ES����������e��~������!�^�]~K�l�<
?]�j�w񠋙�������*_�:�|���OK7�~6�=��˦����8������g��>��D����=Z���b+|��h����'�BߴD8WҲ��l=u~�d=�q�MLt�j��jeL}{	�w�D�/��Ar6E�p����%,x*��h���P�F,/{\�o���Rf�lB�l8y����ַ�t�H�+QĢ1�}s�E��볢�?���o��,$��N��f�o�Xpy�r�S1Y���� ����A�ٞ����_�~?yL�׭E�������߭آ�0j'ǎ��Zu��v���kp�?@tX0�VB�E�m�ώ��QA��������m�f�ѓ�'���>=]���Ҕ)�����{����N!�=��ɫ%�>�|���ݑ���+�����=�i�ݝuB�Z���ܓ��͹��R^W�
돞B~.�U��7����,!u��] �?�x�gB�}��(\0ik����.� O���M��k����w�͸��/6����٩P�ʀ���w���?�Z�GK����zw��^���i�&,�[�9t1�0֙3�<y� HќK����y|j��l��Pܕ�7z���"�!�ժ�y���� d�У�)y�������`�o?;
.���b��|�]�D��2�!7)����ُ����/���'Ak[�W�;��2��ʪkAm�zzXf2��i�?q��_d�r��%�]����ݳ]��n�5f����.��G��~���:7�	�X�4�6�����lp�g�x�,��z#�I���ʖ]��p"�Y<BP�\�?�%$#6R"� 5*�:�^���G��Aa���+�T��������m:~nkX�껔�n`ө������J蟦��ʟ�<���Qh�﫱AP��{��[�݃sap�.�/<�`�MAx�	�s��N�l��B
c�@������wWV��?�g֑�ȥ�J6��D-�'��t6^qyޜۘ�I�����1���o���Vo�)�r Xx�]`oNLj�=\$��%��s��A��u.A�Z����ep�����}�2Y�{�3��Y�U,���~�\�!�i��n�B{ts��/������/���]Hp'��A��f+R9��!B��E���E�v��>� �i�*��q0�����&�]u�JM�İ�F��%�'n�W�vxກ�޶=�Ke�����ؑ��܂���-�MRk	<���֧w����X�����߸ׯ\2ADk �]aP\��<����|^�$�P!��(�wƵG�P��T"$�k�&JH��ct�����A�$F�B���6o閛�1p�������w:A��"�w9�	�F�	���0����iᡡ�ή����&A���9#���'���R��?����������`^�&��Z��('>�R������TS������خM��rcNL�׍���r�q�U���-}�`j^7x��5�s���:��aR�L��	�_.� �JLHL�����k��b�E|���@�=�����{�*�^&�΂)y���U[� ��R܉c�Z�m6ۍު�OU���<o���B��*���1��霣]�5N�\�����<�'|fџ���5�/�K{��=�&¹脤���x�p��V�;,/����g�($����`"��PL��O�v�=h*���AD@���n�02;Fd%C��h���ej�<?a(��l3\.k{�:����p�{��C�Q��A�]�KD�����b�Vղ?g}�P�F��v�was���AJy]�c6���[�-�blP���� ��ڡH��ߧ��Y~�^G�/��ú��|w��y���^l�kP��KM����w�gA�w�-�5G���cg���	�#�^ ���	�s�BH�c�j͑3�k�D��Լl��+���⎓2CZGsG�1!Q�Wo_�e|�&L���,��|�{y��q=����z�A@�}�}'��h�\0�-���N(Ix}rr�+>��E�ٴ�D���;�����
@D�'(H�&D8)B�0�m��kw�w��H�5&�3~�dc�?{]F�09�
�3��G���gH.�q�H�mQ��q�2�<t��s���a�0qŲ���ϕV�܅�@<=f0;��j=��jj�>֩[��O����H�/.c�z?��sB�KD(�N���@#\*�j��/�mO�7tKe�y�в���ǘ��K�J�w	6�Ix�3>��q����y��S0w��k:I���u V;\�5�̜�ڻ;,?���@�k��ť����A,i\D�x�axpd_�a���,�(�o8y��,@h���v�iL4Lg�����_g����;��ˁ�]��}\k�5r��Up��$!/s3�̤F.��h�o*o�\i_�e҅�L���Ut2�+�:�)��t7�x�4��	�	� ��� � �ݠ�Z����U��Ē�'���hâ*92���77mt3<+���}`M��;�5z-֥��qۄ�헚 ��!#6�y��sEl��b��=8~7y8{���{�������v9E�4��ca�P�DpB>*'^\���A����؄爬8��}�XpO��U�͂Ԩ_���־���M���+�x;�����$���=���6:��M�9g*sy.Sj��*����e|w� ��1y��S.��u�J����|��\{.5���쮠e~�r+�͂�E�����a	�ʖ�a��|��pR�����E���AM��RJ5,����,�'�ʀ���G.m�.+5�Ϭ�1�H�i�X\�.�VZ�-傘4,Rc^&�f�4rh	r�U�Z.ud�*;/�������w� /��@f�2<�d�N�߃b�Pa4�_7�ٿ;��n��G���?_�	A�E\(xf�`x���[�9���wa��[<-�A$��Ĭ'�=Ђ�LZ
�|�B�����^z����0k@w���l4�뷏a����:��[��C��U�t���$��k�d���.%36�~d:����P\�m�J��~�`ަ��-g���#'`Z��.Ǖָ�ƭ�a���"���/b������5�<�Cs�M	�W*�྅�]\)M���.8���xa�0xpd^#K\��c������Ѱ�\q��ӎBPdG�m���l���l��.iǇ3�7.���t�d��%�ڤ��;� :s@�jo�f�݊͠%�>����rA���pU����� T֙A+�y����Ǽ-ul�փ���~��傻��Ka-����K_}��ܕG#S=� �]�hr��	��[����7�����MTѲ����h&P�SAFǐ{��^�Ɔ�Ltn}�� <(�=�I
[jn�Gq���?���]J�����<B��(������{�����{���vq�$Ɏ���Oot<.����_`���/����A8Â;�p�N�����YX��)��������,.k�!��0 ��T�|�'���g�дd�k�V�5n�I���Z����������#p���g9.*E�����mw�����'��U��li��*��w��ZŲ�Y���M�������������2��@���E�Y���Y���b��W�j�O8��#�R�`���m���n�76����\/�'Y^�dAR�b�ۙ������w�M��-���ma��"���m��X.�s҄2i_^��of;զ��18f��|9���n�Ӧys_��H�;�a�v	�h�k�iD"��0Yq�����`��\&����U��K|�"4N6P E�>�-X��@�R-�_�5�?�rLy��n��.��	N�Ω8	���v�`E<O��ܜ�>2ã58��ی�,Ք�	�-!r�+�ٓ\�i)�Y���� N�>c���^��������/�9��H�����x�Ǽ��������,�0r砞LP���P��&�|�qq���w?�?��!Fc#ww���E��N	m�;S޽s
�}���7����]Y��9�,.�#W����C��Lic��W��w��p��[X��w`Z"}�&0�QA.��&�݃��s��-�랼��c�*� <$t��~�W
�җ5�v-4  ��|f�ǔ��Cxx���e�����v����e��h�������� ��-����oX\-K����&�	
Y^"#]��q���WiBlG�����.RYY	�/_����FyAp���i�\��\�t��%&��u�߱���.+6�cz������ ���0d�N�w!�k�H�� ?dჷ:Et���*����F.
���G8��, $�ג؎��Z}�U����0'�9��d��#���C��fZw=d��0������b�t�uIU-���RX��Y�����z�Y"�m=��1��WM�]�����u�!%����e�Y~lSO-����^&ԣ�>�1Z���g�����X�`�_Qg�gV��߭�#��+�\�\Y����p���ӁE�C�W���}�dxp�r��w�vD�� ��>�&�w<{�0��o/�U�
��!�?�2���^�,@����{_Ht�����`���p��,�uI����e1]�<�x�O�88}�4���[p���ѣ���+���Q�ŀ�Z�Ks��,X �1sf0��;�ٳg;�G�]+b;�7sQ���k�?>X�VV��v���?u����i\Y+4g!�z�jx���l6��̚5��~��x���7?�/�f�x��7�b�����3g9s���D��aZ��W�.��&	�
��h�p'��a�����J^��<��!��@pw����x��"hp����\��$h	�^raWYQ����u����(|��(D*�b��W��'�#]-�v*��`���o������-]��/��������t{2wtC Qؗt��mꢩ�UE�-�;|>��Ô����Q���PX�P.�f3�>��|�CR�`r�n.�������s�U33S ��x�<=�T[,���5�.�<�E�Vx��z£��^�q�O`����0�p�-~Hw��bk�~p��U&�#�����%�NKq���p?-��ඥ��LlG�?�N�b»���Sh���+V8El�?��S�<y2DG�����⁵~׏�fc�Ǎ))�zvV�_��E���aҤIХ�c���?쇪:��}���0>^�h�r�-����^#�]Vj8�f������Hp'��� � ���Ñ�;A�Ǻ�g���}]^�@�(���R�����VmՔK9�F��fK�ol?s��1_���&A��ߛ�3W,v^{�*w7�cA E�;�[����vM`]�d�a��\?[�r08��E���l
�M��ґ{�{l��@<�*��:�M��w���矁=/C���\%��A��蛔I��(w���%s�+U`ʱ{\���=�@nB<��7,��;Srs`hZ
D2�y�c�8�`���p�c!-J;�3r��]9v�� ����\����ʙ���w����#//������󐓓F��N�E{����5�ߡ���'�8E���d��K�Bs�hю��1XF��D$=F[}]s!(Hc��deeA||������+L�2���HFF��5,���`�镹�;�w���t:�fӖ�Ah��n�y�r� ��t���>�o7�����;~}/|��8l;s�	�(f�����<3�����ڙ�K-|����k�{<E�����3�*EP\A7 j"�߾�Lcw�^Z][�/2�$Z*w�Er�x�~���h,~x�?~�V�.tD��<�Ҷ�����w����=���X����ڱm��喞�Xj	�,�Ā�.�剟�������;�i\�trDVr��Z��2��H�a�7�� �������JH�i���գ���O����K�u���.E�}�����0�fZ��]=w�}7�5�Y���A�\����n��a��@�+Æ�Ç��2�e1D�Y�;)��>|8=z��	���\��q�X�Ւ�l�����,�C�AXXX��L��d����!L:N7���[�3D���F�	�A���b�G?_����K���}S��.���g{��n�=�<��Q���ES|������쀿�p�x(d�m)n�����g�0a�Ĩӹ����;�D8o\@�x�<|w��f݂�2v=��/��w�p��矯�i,jE7��6[��SAMZ��돧]	�Ņ9�_qA貆�
^�	=��3��9���s�\�<�}��`��\�
���k���|
�����^lw�� �ѣ؎�F�ÒGg�����{� �jPe6Ø��Լl��'r\���{�<v����w���W@mPȼ���Y>0?��b]�G�vL��]UK�r���e��6�U50�Y^P@w/t#��q'$��7	�z���H�Ƽ�ױn�n333Y������;��OWk����P�&��L��E��ڵ+K���ڻ�'�@�(�0�P2����9�w�Ðw�hB[1��N�zp���C,�OM`����vk֚'��N^)��R�k��~<�ȃ�1L0U�@�+��n��cz�n,!X&�O��9��j~QqQ'���	(�{�;/�w<+�I��/�}���jb��X@ڐ C#W9"(xr'�\HY���'r��Y�[�|���	옴bq��/,��n������hr^��&BK�������p����e��/�����Gvϛ�'�	�x�o)/("~1g*T������1�U(�WN��\���b^p���{'��׾P��>���sE,��>�_��;�:l)/�3�a�3w���w�G��j4����[Ypt���~)�-~>H��w�D���%M���x,���o�of�:�{;��~)-���7=}���~6�4����rYg׍/y����JHp'�w�h(���v�	� ���WXzi�6���+Z�y
X��&�\�>�y�D:񩵴mR�a#L�=x�&w�X�(8a��\Μ(*��:��}s� Λ*X�ަ��Ի9:s���M�;�cH�c�CwKH�p�(�4��?�>.�T8�&w�f$��B�)�.�������C��Ȏ�;��
���w������̀��2��.���`\��n7��%h�$�P�^���.���B^&	y�L^�M��{�
��J�Yߊ)92���:Fd�4�K����Q�ӏW����׾���;���
���u,���^��:�&Xq0��{65�]�^Y������`�3�����;�j0���	�"m/͕KFl$�u�����6�!Z���q%�o�ܕG;-Q9Hp'�V`��� ��R+%��A+�I��0�w����~�}`�w�0��bm��;v�ȇ ��&����n]�r�"�&w(�i���Wli��p�c��B��ɷ�e���6���o`�b���h{9������).b;֓�'�úcg`��?������ES%|��K��E���Ddp�.ps�,Xu�4h̋���]FQ|w_��G�1fZ�}�g�~�0/�s���=��g���ӻ��s���^\Y_�:�RT0��IcyA+ki�u\dג�.傩�Y�ą���EI\�!hM�;�k4𰴽H�-��=,���`H��C�c�uܵyϴ��	���N���� �=�P�#��#Z)�c�n�&Jc�-�p��'9��\i9���qSV�-�?K7�3c���j�F�u�@��f	V�=*�11�	\���ܶ����t�I����c'h�"����vtà����xi��s[(��Å���E����{�%�Y���|�O���v|��!��ܥ�=�cBKw�/��o������Ⱦ�ܥ`^D���Gf'Ä�L!/i�#1��=PsV��^�O�	]ϡ+4���/�Y�#�nµV�.$����x&X�8	��Zn铭Y�]JS傮q1AWtD�쵙abٿ�iW ��
�q�߻l�Z�PUU��n�w��J�V:L����=z;�3���R�^�G&r��e�r˫��p��%�2�3����v�MH����_�N�cR���0�}PPP��z�/���N!rU2QB�7�R��.����
�#�U���� �A����Sl3��B��k�w�c�i�}�~���#L��/R�����Ne�/-�๢�.��( �B�ĝ;5��Q�xO�]#����0&���Ja��j�:i8�� �	����E������w�3D�i��l�Ƞ�D�5��w�b�Xh�9v���I��z�ݾ�Hp':��j0�LÁ ����3�x{�l6�Ơ� ����V��H��`Dq�Z���,"K�j�]{�<	� Z\Š���\�D; � ��d�kp�m��c,�:��H�~�up��g;���ˠ`�é,��d�փ0�/��"]%�d�A_sk��:��w����zr�D^D+�fp���RaXF������[���T���nɿ;��j�JAAAD�fe��z��y�u�B�w��pG� 	�����0�"�>;��}l�	�zLZ��8t��{6�� �u� � � � o�,(�����'d��D�����j���Hp'����������C`F��d����(����R~�	�޴>�u�;㳐 � � � ��?)+��{I� $���  B-]�K�
�_���e���Av\�2s4<?�:xy��h�!
�BAAA�����UV:^zIVсw���t:�	��ʋ�z�� �O��E{k����_��[�֟8AAAA���eӫO>��w��0v���8�{�*:��uQ	��E;t��caDV
h���hX��t�z�)xz��`��� _���[
�xKi0Xj�f� �Av�0��8��6��兿VN_c��N��WqA��\`w���AA�L�<o����J}?	�D��w)c�:f�A��]�{«�n�`��n��u����p���b ��"Av�H�:f��yk��,���M~��1��>X���C0X#+��������_��u=� � � �� ��'�^y�_J����W�R(�d�p�q�����ԘA�e��~���������'� mPWy1�܁Sz�g5���f�� ������`�؏�lV��Y]��x�m��͋���8Z��-���s� ��vc@���&|� zC0�	�o�>Xx���`���G6[g�T�6{��n�ۭ�j�h�qz#( ���R���35�]o�y�ޯ��_���AF�	 Tð��%�l=��=�ڻ�Cu�`�e�#/�Ӷ6��v�A�����б���/��z;�c����U�'䁟X[	1�� A���������.(|;��/�^}��J�	�ʣh@CQ$����p�cB���{�Ô>������$H�o�Ah������兣�3#�zՊ��BO^�����D�	�����Q�����֯;����?|�����G�&��\]
���E�o"�ɾ*�ۀ�*�7�o�	�,����,k�؈�$��B۪�<G5z��"�@���P�^�Э0<3|	�.���!4��~���z�f�-	=y����!����j�i��A���;� 6�a�i�܏���$�+�0�j48(//��(P��n�7z����#�߆��&sz}�6X��FEEAXXX�c����A!��[�T���V%��'{2�#W�v���p'�s���\j�(�j�d��+�	���/�L�9�]
���6[���ҝ ���n%�� � ��`�� _����L��"�/}��O���$��@ee%���x�7E!�)Z+�[�V�6���7!��q��W#��4���k�۪ �>�3n�
��_n�.�*a��| Beld�NAȌlA���B�;A>�oم����*}��%��a�	� � ��Y㆕���rd��U���	p���Xa	�:�էF�A�mȥA��;����0�{b�?N�;�&�O;A����Z�0P_����t��ǜ������{�F����f��D�g�0�ޯ�h���}7�M�X 5���!�n��AA4��\����|��j^����]��)��<�&���I��p�&�_1h�`�xc��	g��q6Zm�
�� �g`��S({�7��XcP��ݭ=6t�Vk7�q:]��~L`0�:C�@y,y�Y��/��Gb�q�H�Ւ�@�:p���A���ս�h5A�Ϣ}��R�kL){�	U�܉6є�^���ju�7A��,��1|xͯE�ȃ/v��犀 ��R�-;�n� ͋#�N�K�q�F��B��*O�p���r�F��'�	_Ǽx����TZ�ݨ�.���5O���Fێ#v��5[�8�}�2i���p���ho�WHpo��|������?Z�[-��|g�"�Ї5Д�V��)M��D<��Pyy�xB�s�-���x~r�kOnU�DHpW���FmF^�\Z�]zxw�6�w�����>c4���B�Ӧ��:�6�;�����@IP\�N�p�|}!Ɖ���fq�u�v[�A�ۃ8�Dq+::�zy���a�*��]�E���(���RVV���5o�y����-/X�L����Spp��G��}�y����`��m��K���������"��PW�>�9�)�o5E@@ �KK��OC:�}���_���
������W�z�S��f4ٽR��R[[��U,b���$r祮�N�K%4x��§���t�z���_��K��\xg� rֱ�qK�=?44���e�����2o�1O8Ό���u\�P.�K�A:�OF��|�X������'��}�i�S�A���UE��o�h�ɚ��xZ���5�I_�ؑ�'�aQ݁ ���-#!/9:�`J^,;�Ax���.ep<�b�٬�/[�q��rN�O�H�d>���Ĉ���v']8i,))VT�q��JI�K���y���by��������XoKK�<((HV�qX.׼*�;�)�wb^�b�x3/���IHH(뿔^ls����h�l�mh��r�			�/x�1����F�(���f&��x�݈�9�:����V����x�7/AB^j�ܔ�U,�����-'XoQ(Fo �	�O�ǕJ��{��q��[��Z��_>墳�HpW���Xž���VJ`�O�$�!�� 4Jߔxx��~Йxz�`�	B8{�QP�8)�ӚJ
NR������;�7���¡���Ehh�"�"
�ee&���E���h��P<�[��E",���2�((��n,s���x�pQL��� �.�vR(^;9��}	��u�c4��
��b���E��c�BKdo��ϓ�aGAỴ�����bn��ж~��d�Z����5�ZڃXǼ5��]`����u�amʋ�;��6`��ܤ���jFlGHp�3�pWS�=�s����2�O�_�m�D����{�?q����ަ��D{��BF�d��	��"��'D�[)p�U]]��*C)��
�J�e��hY�4�x���R�u����}9]�x�Z!J]�(���`{����J{Q2/���
o�
q�K�*�V-�o��&��hʭ��(Y��o-��=-���!/%�}�Ҡ���b."�w)�q'��m�!T+_�pl��R��t^p�i[w��@S>ePl_���]�1HpWa��Q��ݡ�o�<�˶͵� �F3 Kj��B;	�U��ف��u�+���t���|�C7�V[^�u:�96e0�Yn�	���Cz��N^FmjpB���:�8����'P<VZpǼ(9�C�LP�W���,������٬�;Bpׁ�8�%L��X.�&����+	��ro�wG,��rewR`���_I��ъ��q���y�2:[� qAEJ�,\�Ep%��1%v�S��X�Q.�,�������"��BqW����;��uLI�e��]5�;J��ؿ�5/�vk��:���y��B������5�� | �o���Iq���'����{[W	������N����(�XR�P����%�R�$<�|�+Wl��"�7A���)e�,.�x�\P���TT�BK}o�(�����;�����J�v�8��N)(��X����ȋw�VѵÊ�Lt������))�L��8�+Dz���,1/�@��)�M��8�Xˋ�uL�u�)�����J�1o�ELv�O*�����	� ��A�]���؅`�&�Ʉ���A^�z��[�q"��5����-Z�ykR��N)9�5�7'x�ﾺZ~����a��Q.�̅�`~�%�8v�*��ۛu��I��b����sX�ʿ��v�ɜ��t];�v��(
or���^���J���8�����y���c�V[ؕ�6����r������yJ�r��q���Ѽ��[����>�|�S;AÐ�N����:3�z��Nޤ=�B�K��WU5LZ��~��+�8��Z�&&&z}R��򡲲ڹ��~~�x�S�'�K�$U�"ܥ�b��B~<�/����'^���t���ZSK'�Ҽ �k��䱩���5��a(���;^��ʎO�џ6�_)�M��"�T���˥=��D``�b�����Qf�E�];h	n0���]rw�{��͙o�1-�뀟l�~Fc���o1Ľ�g�(5�#�C�L����_���t��mP�|����3,,��A5���׮����뛿�q�ߚ�a�j�p��]N��&�>������H��ր�RVV&ۂ{LL�jy��2a�3��5m��	�A~L^r�t'#2�{:���Ŧ|�9� ��Y���#��8�>{��,g�F���s���K\���ӻ�E�rIMMo#͋�u,--���ǲ�b�.v�;ssØ����pw�y���r�%11��b��^��ڡ r��gFFW��{mׁ;(���V0/FcH��g]4Bg��n��:�l�ңGN�������ҝ�C�`���ט *99�^_d����v�,ߕ�� IIɠ���PTT$�wy{!W
�k\<��"�H�w�f�^/�?�| �;5��l�#�3Y����Ddp N�?t|�KD��]3]�|�Z-Zآ�!P��Z��28��	�������ǝ��:���\^a�ہ,��[�*�,ko�n�l3��_N0/j�ו�r����:�@�k�������HD����hm�+��BZE������'����O��	�A~
Zv�G���OK�M�'�� �D{��}��P��UC���ȋc;�N���j��#/���i������]� (���f�̀��Z����w\��x?�K���ZZ��U�������p �����/��ڋlr�����x�Z8��W��>���AD#�"Ø����Ax	��.et���Ɍc�o�}��v����b����o%�q�D���F=�]�r�"�f �ƿ/��qG���kH��P^�oW��ɍΏ����O�2�-�u<L2��-��ޕ �p!>L=?sZ�w��"|�|\`�-�Q[�a-RQ�5-���+N�Q5��Qԕ��]��4,��}�{���u	�Z�h���:����o\���!�^� �SK^}j� $�wf��N�	����:�?�
Ax���5��������".��~T.�`�� �ȓD�X�j�E�_,_��*�w�җ�{��I-�PƑ�vvm���aoS�R�x�ue����^��<�=P��S��G!�� ������ޡ�� �
� �D�g6�Z��I�Ů�gF	�B���_y�[ S_ԕ�*�Wm�@�:����)�]����NS�_-����w��Տ��/��p'�V��?>	�A~HBXD�Ќ��A�����V�ک�)a����y�wZQ��Y-QD�rQ7ؠ�אΏ\d�) j	�'�]	x�����/y�x��{�0$�A�!4Fk�mɦB������dF����K�r���ǟw��Ұ�cy}�QOG�����B��y�J�m�я!$�+�w���$�>
G3��W�*��l7�l@�v'�r�����w�}���x_�:&�=��͇z[i(y~�D=ѝu�C�:F4�?�	�W������Q�L8����/Pu�\� C@5�0$�A�!�3��85f+��v*M-}�/N�l6��ą9�Hm��~k�y �U8��X.�,�kAt�!�rh�D��/z�#/�!R��0��lN8�}��$w� B[�-)����B^r<tvL5u@����d�H�)�����n���5���f��kI�.��-��nW}G�\uL����F�E�5$�9v�h�|:�?���'�K^�·�1=�)/�Kע� �,�	� m�o~��'���τ���b���*8��1��/�����)/r ���ZYi�E!���ڐ��gxZ�p���v�?���k}��
�GmUN����QG�_��/��i��;3����R� ܨ�5��{�:2��[pWs��ȋO����ܰ�Dٱ����hT��s�u���KyB��.5�l�C i9��UP���8���-�ƒ�Dj��T'�p.�/��;�w� ?��w��+�@�w�8}�����b(����F�v�����1/8�Z���!r-P�␚�y�l�Vy��5Q[��C9qG�����V�-�2���)���Ý�r)���$��ٷ�_s���MP8�0�h7��\� �CG(�����`���6�)��-���܋:j��K���!5Mt�#�஦�.���-��O3Os)�/"���O�q�ǥ��"5�Ga]'�yG�;��а� ��:��TTAbD(tV��,p�b1���q���QV�c5'�����������b4��W`�4�f{1����r�}x?r)ӡ:��ϼ�^O���) b]US�����=!�d��q�̥�W��C�{']�i��� gJ�;���c�%�Ҡ� �H�G�"�"�%R�Q�e-�'�r	���UoV�� )EM���\�j/<��Z��d�ΰs4U	�v�p�"��a�t��y����N�.6 ŝ ��×�Ẍ$�,=p�+��q��.���	��?h��=�����,u�0�)���kU5p���U۱��&������ڠV8�:�q��*|W5U�@����J��/-:"�!"8 "�`��"8[R��؜�hH�r,�j1�]��r�^����IhhY`�	�p�7E
˪`י�.��9��6c�*.��G�ûێ�!�M1�G*X%y?~�.�7�c1*8��Hg��c��f�m���U����!'!�!&$��k�����^�6�<ߦ��ct�4�Ϯ���^�
�)`�����D">>bbb�������L6���@-��#""�=�!�D�in���U3/(R����񯴬|�)�5Q\<

��� v�x�b�X���Xf��0�����-������@!/�s�F���׌���=\t�Iĩp�~՚kA-�������'O��55��k`0�;�ϳK�.�^�s�s�>�r@��b�0����V�K`` ��ݻC߁�y	�^0�5�w��b[q/�;R�{^��u�9傟��PM���<�1l���:\��E-�kj�%;;�e�M���`���c���}JM����l�'���$22��>YD����-��vYb=�J�f��X\\,�;�Q�G�G����?��8��\��a�3������N�4��L�G��/�9���W:���`�x������CϿ|ŕM��H��P���I-�F�0�'��G��绎Õ�j���L��n��w� ��5��
,�w��+j�؉����	.���d�G�����0w� ���{�]�?6��7�	�(ࣨ����##z�C70����7������[ࣝ�=`�?O�f�
�{^ �]/.��ښZ�����F�5�����V�+�����m�zB�������_�=���\�,U�v��D�� a�b�ŷ����'P���`c�K�2��u�$���NUk欬,�	�3@���`]/L�/���������ib�,B{�&Gj����޷o?�X(�G������g�"'��2�Y�`	��cy���#����=&.���~�y	����`d僋|�Ei��w��6̋��W�:���1Q��}_��^J��T	և�ҠA��c�$������b�/�/[L�z�AVV7Yb0�%%%��_m�?.�b��v�h3�El/:7�u��g��m���m���K;V�����$�lX.Xxo1�i�/��/�Iq�����cQGh'B{�6�ֺ�}LX��^������4꓅d�5�/v��~�ncu��lQ��]4���h+���~�>Ҽ���v���_!/v+�,�����_ay�'�P@Z.�9�m���iǶoU%/�.���	\n�,߇y���R����('3SV+{�M��h;^��%���a�1���VQT��G�Bi��{	�!00-���(ߜ����,�����d���i���
�u��]�(��'���y���#𻥛\����� O=��8(�I��܁�����&��AF��ޱ���Ͱ`o�:��jSW��_�󙐗��9����n�g��Ovo�y��c��=[<�wRl��sZ�n��;�����wfO������\����#80�Y�{��i�d��I��#2,*kj����A���A��&ݭE/����U	�YY��'yAB]FQ$���U�;���9!'�m�����(R*L�-��B�KpPP����@�9A�<X�U��
y)�j����@Tx��߉m&>&�KM^w!�B��(��v��[D����R[[&�ɫ傻7�����D!�\�c����MZۏI��@M�5�u`*�t�a����ܱ\>���."wm��'����RRV���K�po�:�bnk��:�u�T��fu��닇8~		v�5�"�ul�L�O�Џy�\���*����Qż���?�󯬮��*�-��y�EG�*P�wE���q�5S���:���(1.J��T׶m���:<���o�>��(�����U�z���ܫL3��.�`j��Sȍ)7$B1�Mȓ�}_r	_��mB �u����)68�����{�m�K�,��zߝ;�V�2�;+ό����GX;���w����y!�!�᎜����4 %,n3ԫ���}n���uΨ��;.���7Ӥ�W��T�mnT��@��'��>��f�����D�4����pP��Qr��jZZm�y/�s:>g���UA_�?��)h�݅3��9��Up��R��һg�
���iɢ������/���N�8H�����̳��q  =9Y�"�B%���Xa���1����$��0#�MbB?q�Wi���-�^)I	~4=�m�y��LW/�ꨥ���]�&%�ꄂ܉Ya��d��lw�e�����2�9��A�X=�l!��=gi�y۷�-\6��C�ͤ����l�}�&%vЌ����`�5�~o��w�KMN���3/�������n����_l&�������X�fA[��K�*�e��㨿��������3^.F�
g���N"���kz�Q���S�	��U>VV�X����lQ&��5[�Md��&�"!��G�Aw�H��ҏ��}׌����o=vƒ��e�0��]7r%��P}Kh�'�j��#�4,3�F�?�R�|�\_��k/��6|t~o�9NK?�Eߚ4F��<��썃�N�&u}	�_�Z�T�VgĦ�Em���(����	w�5�ϝ���ʇJ+u.��������v׫�
$kM��ʱ�L��m'�����py�x�׾9�Fg���8���y���W�%+\;b��v���5���Q���)��;�s��L������c����6Ս-�[Ew^u]5�y��ܕ	�͞�H2_�d��Q_�x������E]��j[��k���D�yh�Ό�x��J3�HIJ�f��q��t�n3��	gP�lw� E��t���P'��^.t���2��L||��ma�9�e(������&%��V3I]�~um=55�̪���2�
�t�rI4}�p�0"rF�i�dn�z|I0���c¨���sے�n�f+y?����+���03p[��%.���S7#Ut������8:r݉c%/�j�(�g�d�Xiv[X������;�C�;�1�$�E� ,�σ'�\�}�ݖ�g�O�PZ��;���	m���s5��-ۜ����K����<^7m�%����0}i�^Z��-�s�8.��u�Ͻ�'�;����;ݦ1�{��y<�����_?�1������w
&:@Ψ�zp�8��;?��];���K�x{{�qz��<J����l��Ab��b�����<�g���:���>�w��ghz
�7h�D��/�=ۧs�����[�̊��H��"V�]��(���v�)�j�H� ���_�VT���53=U�m�F�;�k��O��2�5��	������[M�������d󃺌��,nK�9Aw(�_?k��ݮ��u�9���ϭ��3:���������`](��� �dR@������]e1�Z.���Q��K�=�,��bƝF��G��X���}7���b� ��x��NU����0����bf�;W�[��Δ@5��hr'��c�걲��Ɣ��'Y��Aw�ï�#Ԋ8�"#�S����;@��g�I��x	M1���no�QK��k�r=ӬhheU8���	�C�7x]�v8�hy���2�,��nC�4��1�a��?a���.�MR�lMC�4���6�5ܵ2��Tr�7xz������T�Ү�m�=i���?�c�O���S������k�۵a5ʨ�4��5Ho��\WmۯY����_Z�w~߾f<�${�B����� �`;S�P�|agU��Ed便Q��Aw�����:)�f���@��0��D�j�����Q�uL�u����*:v���� ����ѹ�t��	bA����D48�#�c5�s�`��"]�`�K:�T[/�B��/��!��y��w��z�D�d�*����!�M����v>[�Pߗ�m7����Ī`�����0F߁ ��Y|�d�>�^[��ǌ��ɩ֞'w����d$�ֱ��;�1Iq��@���E���x�[�k�I�����o�l�D������St���/&�޾>]��q��^`4�P�A#P�ܭ�y���50!�B�ݭ4c�%"��ݔ�л�
����e���^�Acq�=��2���Xzh�xZ��^]�~�`�i�!{��w]��L��M���܀������%�z�����>Ӿ:uV��*�����	������X�N��UO{�_��n�7����rmUI����:/Zd�/�����b�ؓ�n�<�w18��<�!wd��M0�-�Mş�K���>#S�@/�^&����.��:��P��$��W߿ΐ���䄄���xW:?���ܷ^��rQ�r	�]1h�+���]$�ebp�`.�ҽ\x��z�����F��?3g�;��1����pq}~�v�F��UF�kKr��k���q��;ױ�6��D���5��ȹh�[R�������O2~�W��[�����//1ت��O�:���ptm��Xdل�Xw{x�9����ƴ�K{��۾kY��Ovv��to+���--��!�>�)��� ���Kd��9��a�����[��._(^&b`Q2�ӽ-��F�����ü���i�RxR<ֳ���1�擄zeN��0��{_�HB��O8]]G?[���c6E�7w�l��8��j��A�w>y�����g�Z��&�����#��R_�����y7��ܫ5��{K|k�kѺ�����i����ց����Zu�c�d�j�e�O�.֎V�Ҩ��.��ͣ?l+�t�ۥ��<��no��_b� ŗ������{ �I�70�gzO�#�Ϋ�:����L"��Z����k�r�;�߭�H�����z�~���p ��<��"ͽ	F\��̣-������
ܺs=�j�����������*�'����V煴'H�с-j��Ui_szl+D>���Gū-�v0+�/���"~���Ȼ�Y��}9X�~��
����g�&�����p���,S�u�w&yN�
��?v�ƪ�����w�6��������˥��Gk��Ύ ז��3��8�<P���1�����}��C+Â���/�Y��V�����.�}��9����;��bp�_�����oǂ�q��������
��"���NU�Y�E����PQ]�1M������������+�&2���Z�.nz��4�I�sw �F�A�bp6}oJE�����ڭ����у)��6ߊ�&:[{>xXx�N�*jhTvg��[�po��p��Q�it��ܦ�׾����a�3�]�W��L��Q�&>F��A��{�#�%�����{�r�W��w�v?N������?m?t~S}�uځa�;�'�_kqD���e~>c0�q�q+�1�F��Q|�ʸ�c�e^��mq�W[\����{-�|�/�7����H	�Z��g�@똥{f�"���E��\߯G��[��H���#��d�3�)�9#���鱽X��iE�Á�;�3I��� ���������f� �$����ꏨ�ٺ����s��qkw�����\�Iܮ3(u��A4e� �|P%�j�z̵�7:�k~�2��42ս�Z�p���E�*)��޳C�ި�V�ŶSe��p1�{�<̣3&Қ='���V�~[��rk��n�����[����guVy��z��j{�-)�l�   �:�b(��7�H 蝢:��p���N���� f�����>���4~@E���~�e�d:o���\��!�)�tY���2�g!����)C���%��Ր���y#�@,O��W�%���^Y�Z�m���]R��ڝ��r���I�G�΀�,���peп�����;=�Z�=բ1�Vg���r���&�,��Á���;  @ ��q�\G  �Ȃ8b[��G��p��{��R� }���������Ewy���k�:@+6��=���Sz�;gЭ���﷯KY���m\��{0~��}�_�o�R���j��$�4ʦ��);��m������hE-���(}��1���b��뼏�gj���A�5�s���I�����l��h�������Uh|�!=��lé  +,Q� �L�)�sI
s��aQ������k��~���y����t�x�=��f���F��v�	9t�gߡ����9~������t͟KӬ�v��>Q��u�����^6�2'���4s�o]�c垃��6��/I�@Gy��Kjt}>���zK�(9�)�m�Mw_6��־�Y���[�FxL���15��ϴ�g�/7���]��y��镭{{4�V������Ow�</�M�Y�=  @��  a��Nа���p��$rj� �Yt���5���o�)r�v��������qĹq|��t��lg�2�iTV*�>eeC3�t��4.']R��-�ػ�vJ�Xz��Y>Y���mTPZ�1�x����IN�|�h��7���w
�����^�� -�}���x�7+��p�Ǵ1]�ߺ�2=3G�n7;�΅�9�~_I�G��`��,���2�i7�JR��Nw{ϔ�M�{L�9r0��NG�USH$�  `��JqG�; �7s�ɒ��;�;�M��� 2zǫ��s�Ϥ�S�(\���(=���!5��D�?�G{�\]w�^玄��H�~�� �������iw���d\%e���&��Gf^J�5��:�Ӂ�%r�s���9)�4c�@�_R�1P�w��"��w�8�����ee�����x�`�1u��:d��Aq8=�2<3�NU�Ҷ����y��'󮡗��g�n��w���u���`�+�1���m?<[I�!|�o�<BO�0�c�q?��{�Э/�	i;sH2�   t� � �EV�~�T��{_���v ��7�\��(*��~�����<�!��|������5j�ϴ��V�{�zjS�K����;f��R��3�^���GIM����w�i��wRr\��kNɣ�ş����y��;�NGi��y���\�^�|~���bT�c�����w�ߋ�����*|���u�U^e`j-[0����w�#��x��F�~�}�����3{��Ѣ�y�.�j���A��l������{y��ݖݴ�Y�Ӹ����累�S��L&�d��y�|��_����T�N]�\��?�y9}r�4}ZX��oy���m�C���Z��s����YAY,���g�iW�9:Zn'��p���2|]���O��c�������5klk��w����w�^޼�{Zs|jVmr��u� �X��8�b/�J!�^���ho"c�L_�)tkHʺ�!�z��&���,:�zV���@�1>���&��#��)�z'�$�b��k���$2�S����{_&I(( ������}�9�eL.���f���t%�r��A�9����>�^�D����C��23.S��8�qK�o�lw%5�˂pM��WD[x3E�%�Q����0�g���/�8���Mt��V���������5�g�� ���*u�:��zO���I��dH��8����U�ݻ��k�G�)�h�Fi-o�T���4m���K=0y�߿����/�d����<j�?���hڒպ��_ݺ�n�NS����s�����N�s�EG��g�ui܀�:�s�wϢ����o}�9-.9��i� �R�NZX��ѓM�����#�5Z����� �ZJ1E ��6� \��Wޡ�Mɣ��8��{GB��xf�VQ��b� �{��-z�S�G�i��~y��n��{��}�D�vƙ�Srshӱ3ߧ�γ�'������sE�^�K�w�Uc蕭���Z��Uӳ�>���K���'�n�g�O�U��,���P�=᭺�YtR�R艓5M->��$�s��_o�I�{��sZ��������i��_�	2�Ο��/��:��j�xI�(	�K��7y�ڶ_�<�M�\��M����
�E��`;kn�o��:Zr�,���1A��'���1��  `-E�=�  >$�E ��6�Y �������Bzr�U���ydi[�kQ�|���h�����ɤ̮N�O
��n��2����矵r==�Jz`�$�~Ԡ����L�����Uu���Dw�p�z��}!���N�bu>�'KE�MGN�����vӧG��7M�9c�h�������ͻ���]s>�M��N���	Įp�k�Ӕ��&�f��^7��zv�4��<�Y⭡�����!���|�&�n�8�g���i�/�"����m��K�f^A?�y�OI�������؞y����on����?1�*�2l i���8]Fϼ��v�8@,     @ �S�����>M�^� ����6�?��K�w�}׌��g\�9Ц�V�:ڜ��Tz�~jXf-ߴ�>8xҧ��?����饭{�+F���d��OV���_�AQ6�l�$ʨpƴ�}%t��5tݨ�tk�HQ"e\N�(g��H�P��}��;�r��f����]d��w�ܳ�J���kG^B��)�3�R���j�q���`�ז�M����K!d�W6��W��w�yV+hn�������������W7��>8��'�o��l��f�B�2R�Q���Q,�]��A�i������b��tt��ЃKм��NZ�y]5$��g��T�����v��Dz}VX$~�&�չDɠu�<�@���T��v     0�Sn=E �>L"*�=a, 譸�3�~�u�=��4VԎ��{�g����}��?UJJ/�A��R��DY]�ؼ�g:w(���h��_�Y���X�]���Z]Vk����ߗ���`j��ď\��U��F��0^7��.$��1��.|� ���(�/�9J      h�a1M�0')�� zq��'�OFB?�~�`�3f�9Xd���V�'G��S�g��R��    Ɛ���   B�e9]d��a�ǎ��Ͽ0� ����9�ו��%F.�E���h@JHN��S�Ŋ�\2��������4��1��U]P)    �I�QS  ,��#!p��*_|�l�S+��N$ ��%Fx`��2�)     �  Dt�"�}���C���;         \�� ��Aq8ߐd�/ee         �z�6g�v���q�˞8��Ԋu꯷         ��$�~\�tQ�ԨE��)9�SV�[	Y�         `Ez׾���=J�w��%��>��5"i!         ��`TTӿE�����t:�r����      aO�]�  �{KQ����ROw�=Y������c�         �$�p�����"�Э���H]�b.)�w         �Xv�����G(B!�n$�&����׏���      �3�� ����$�u�}bE0��ӳ[�O-��F��D�p         �0�伡n���(�!�>�_X\���K7�$e��0�       )  p���2ќ�%�P��;h�_�Ha��˦v�l�'      ��� ��J۝���e��`;C���|񉳉���C��&          }�Y�S��#G�A�jX�X=�bFj��<��!C       �g7q�uD�ü�+���M��:o����U'Id�w���*)r��YC�dZ�-��fEVZ̚�gW�`"��F�"�6�hg~��?*�>wn�c����x���(
�R�d     xkT�H��P=IR��N}Ã(�2�\T
)K��&�g�$E�%�HTCNٔ �Mq�;l�l76��Ô��洵8��ٔyK1�ɔ���؜��o޺ &p��K[����_��c �r�z��O�Hm�lR�$i&/K�6�²ڝΨ'�yOoq(	N�d�"E�*J"X�/�Lʼ�8+Ť ���A��i�,Ӳ��TC�IY:�bJ�SR�3���cZPHR���כ2o��I1%�!)�6�s7�1oY�V��iJ&Z�B��q���j;�8�� ���~�   K!�!i\��9���R�\�I�T�}v�$��HJ�������q2�D˲�@�M"G���H�Im2�ߠC�,9b$���dE��-���~����$EI��W���l�:*b%)6@s<�+K6uc�!�d��Ԗ\��o�������?�ϳ�S�u��֨�"��R�(�ڡ(-�N:U֪�*l���j��NE	�R8I��	6I�C��w^\мIR��4%��n��N�9��(RZ;b�L	6%����Y��)�M       `���d��MV    IEND�B`�PK
     `+�[�AWv�'  �'  /   images/97fe1122-b934-4e82-b9ff-450ac31bc7af.png�PNG

   IHDR   d   G   ����   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  'IDATx��}�\g���^���:���V��%c9��f`{�a�s`=g��93òs��viI;,qI�����%[�[�[ju���9�7��W��:Jm���:�~�7������4�G������M�XUU��:4��U�z&1�隦�����Q���I���eK�p���ͦ���5�5EA�R���k�	�|��o��]�����~���Տ=��i�`9���&�3�ejE����}D���G��p��\�yV<��k����o6�2��^, Z�N���͊��T-��#��ό��F�&��I�V�۶���ݵ&B�?=�~��)=����+�F</����77��u��yI;�%���ȉS�pjDz�9D�]Q�}h:�^�֦��_i4��OVT����M*�Û�:��T_�ޟ���C�P��1X3Y�Aw�l {^���͚�+�[C�uEX{��.]-���j�*�jEM_� g(WG�JE&��#���.�??|H���5Ժp �z�=p���ڻ�Fo�y/<�&b�JSS�PLD'd�p�l�D�--x��9��FF�r�
M��
�ZZZQ�q'&��}8�n"B	���f3H&�hnn���en���G<>�r1Ϫn���a��y��F�e,�C2iF.�C|rR�2�����N'� 4�B>/�V�C��	.�K�Ô�5�r2n{kz���_0Y>F�XB�&k��x�o�t�_�{���LH"^�����&u�{߇��p���!���g��U!�jMǪ&�2��-&��\�EB���<>�قX<��	�ha�t/�� ��b��L�*����Z�;Q+�184���#��j�J�rCã�s���8�;,4�����1x�l��MC#h��d&�H
�7���kr/L!�B�	9�h
E���D'&��ց�^����^���'�S�i%��!�ji��t��/���Hw�a1�����.3��e��C!3pf��j��s?�)�o�k�Wg[}j M���N���M�������.�O{��[�*��cmںM��R�7c/}�o�I�]w�!}���X�Z>�����x�ͷ�Q��o穓���D�u3���w��'�*�s+׬�B}dMf~\e�c!�޷�fy����[D�p��P{o
�84,v��'��h�.�k�*�H|[p#�G���k��5EhMa�ҟKE�̒P[.��ua��M�dab=� -=ҿ�RIDKezG�>��X��?��C�wG7M���|��E�wߦ��X`��q�V�����hJ����6�3����z]��{��Kg�_}��y]د��&�+�"�֓���ᰚ�����T���)d�[:�p"�Êf�S�ϊ^/[8�}:|N�ѻ�*�a������(��D�^�TA��%b���y�V����hJ�"�F<_B�P��j����"�2���(+�b_<B�I^,�c���U�|�VU#�퍈9,��+�$굓��JW�bQ����\�����3+dMJ��1�_߉YRϞ���6��݅ÿ9��ہ��و�>�G�s�+Ф��A��5��W<O�V�r�JL�H��hcCK~}�.��n߄_��q�ukQ���=r�&�nz�@'��r�lw�����b�$�t�aGg3���Qx���n��N�c�쏴���'ӏ�ߏ�k;p��+����H�I<E��=��a?�9؝v�a�&A&S\n�-�!��2L����[-&¾вw/�|�=z�6����A���FE1k�=r^��������Vu�l�mf�
d�鰒x�TI�)ܝ~�O�V�FO+dM��*�
���%�;s^�dt�tϑ�a9M��\F�w�w� 4�F�89<AT��(d��{��� ��F��1�bI��!�O�3���Ne�`�����Qy��}�D����`	Q��>E��=˖��+ۼa��b���gq��V�mY��hp]�qΎ�Ѿk�p�N@�k<')l�լc�ٻ��%qU&��˄\�n�!���]l"��B��=G@��ʦ�&xm&�u�*1��z��mD�^�_�Ӂ�޿U8�a�����e�����"�YL2';�^�8��Ob-G ��Pd�rYj4l�x��s�<�n�6�`n$�A���1�{���-	!�e���0�9�{)]}9Qi>�b���3�L4� jb�U�e�w�U�*e����_=�L�,��qb�(Y,^+�<]��3�ݱn�,��G��3�&�aR�L4L�<V!p"Gq����c�J\G�P�R`�l|�����8q���������8���pL�3eIH¸��T0��f�'FR��1"uQ�&��c��3�L!����%ƃd7��lZ��'���n�(�V�ɜ�O���~?�������"}`pY�P���6H
���I%H,ؘ�9��#<J�:],��Q=�vV�×�B�YT��lY��9Gt@� @&2�
Rt����H�a���X��N���l*��� *��P<GH��+gp�\M_���D����N�W�U6ҭ����������.�Y�.AH�V�����oF���V7�8E��E&��K1i�H�^���J!j�����0P&�P���3����f�̍t�\���,�>�#�ٌf�È���iQ�p��6�(�}���d���!Dq�<�ѧ"!ǤNQ��,��fo�%�����y��!��G���ԥ�{��/4�����5�}�Oa{��6s����EM�����Ѳ28Q�ua��Ѧ/�RG'�k��Z��5��K,�9��M-�>�K��QIٯz�G�V���ͩ�8K�G�*����>F�Y̰�O�DW���01�C��OE��	����ǘM��Qu�:̡P�~]R�D"0�3yr11����##8% \=u��1$�w��^X)rI��cN[K��v�����⢧>z�N����b�D��}���#ŝ �÷��??u?���h�p\D�l��|	T�\N��&b�-���N�+� ���u���D+�����7�
@��|O��؛NyW,�b�U4����!�Ә!�c�7|
�ɡ9#�J��rd���>��={_|�p����{�(Nۧ9����֐C��?��x�xN@��]��^��A�cQ�+C>2(�!�P!�!M�p��v���y���Ȫ��H*�Ⱥ!�������8���"K3��5KcQ�!�{�����x���h���G^�+d(l$S�k�?����6�����;N;y�q�D�kAAħ��x۹*��H@��H��0�ʂu��<��tG�c��1�d��4!3�����P6��Tw���bV V�"V�u�V|�g����}[GXD�g�v>��+��{wn�k��i���.#���D�,� ~WWI���A'�����R��	�|��?fJ�������F��OW�Q���18F����n� 
Ԥ.�k&��{�i|�/���?��HV����c�0���܃���e�\�>E⥄�Hg�����?;���,R�%M.�̛����֐8{�hqM��C��g-}z��%+�׼q#��7=�o9�*׮xl��1Ό'p����5F��qAS�ۿ�K�^�"~_ϗ�2�r ��?߻EB����N'7U���q�����~]�v;y������Ⱥ��_w�K�����+s���5�f�pfk*ݫ)ߺ�[">4�.I��$��%:"��e�y��DA#�'� P��Y�(�a�3��w�ڀO�y�8���Y##i����x��(9�W�!��?�\����M#�X�V��gmJj�m_Cr�C׺%2?U�r��T��Zd�l��s�%dd	�0�3��xʖJ"nJU���{��HU����leUmN���R_~���v�Y���K���p6�n�X?�7z~���׽��x��9��c� ?�r^�e�G$j�K�P��[`�t���$u6�	"٬'�
�|l>�����a'-�rb"W�w�D���d��ݳ�Du�P&F�B�*��n܂�dB���836IĠ���������,	����fEy5u�\m.濲����oߋw��GPLV<��cx�C	����[�B�g�P	��87ï�����7V����}�n��X;�[���C#r��v�'A�u�a�HN�oN�OE{�����3��0c"�������D��_ہ?��/�לC�zf�|�`����'Ǔ(W��eD���aj���by�O������3�|�T/�����Ș�
߲�U�!��ק�	B��k%��\�XK#˅ƹaU�2��Yъ��\n�����<���4��F��M&�b�RV=��|��ĉ��%�\e�M�u��#
�8��%���:XAN�?��bSsH����;�W���\��0���&E<6�Tyw1�1��_�6���UM~���Z��;��O�$>���N7)E�o�J��л��h"ϻ��m���L�In�f�/��lf3ƲY������QBF�\���ްG�cN��ȓNI8e�s���(>���𡛷#Cz�3���^3Ǳ�KISq�k��/�ǌ���p2m���nx�@���D�4�����q|��$>V+�C�
^��g�H�a�TI��+�X��Ȧ�/�������U5�&��ryO$S������1��������}W���x��riN�S5 ���h6�l� �Pkd�X�+6��[͜�+�մ+��׺����w���r��t����l�J��� �y=bO���ux��lz���W�Aj}�������&�A=�W��	܍TJ�M�W#_,#b7�b��AR�f���O���X����v��,����̍���.����0?�O��<<���ۗ)�̸��x|p+}�R��D��� ���y���18^x��P�Úm�3�cɑ!_�p�۠8=D�ڦ�Ρ�Z�#��x�''A�	"���+Dg�T*�05	S�.m@��l_=>��yӶ=>����ڗ������+#żPPN�d�
�#~�)۹��ۘ�4����Q�j&�d} �*�)\{���\:���Oa���d��B�
��ƞ/��л�ʎ�e/*S2��g��0���c�jՋ�2o<-��,��V�	X��2������<��h�/W��j��JF�^*`I�л�������R��<���!�{�(�k��]�la ���̷�z�}�>�EI��~�0S�x��ev$�Z"dp���n$p:MW�'��fy{��P���[<7C7]�^���Վ�͏W���(U��z�Sr/�b�<�`�<��*�'�N>3B��)k#ߠ�s�z��l�Z��HLo$��f���|�`�� �]�,J��3=(��M�*R�ڴ�q�<�-���2�ym�f�,,�nk1��\;�oEϙ��6l�+�� �\ Q�~脓�'�	�ˍ���زj�+�w��p���A�Vy�i��eR=����k�&��)I�0?�,|`�<��!�.�t��}}*��q:I��/]g	�����gr@��nF@��iB��[|��p��0�"��Z�H�ZQ�@��,�i�P�]�dS�ڼa����aE�<铣1������E�nQ9���b��9&D(�,T�s�3��l�	������Uzn��H�.��Y��ײ���dq����]�gДź�A�d�#8u���KkIE����!��ɤ29�mf|�ݸ��%[�����#,:g<����$��{W��/�Ð����J�3BdC�j-�k���x�7��۹�۷YR����+͕H4'a�M6��gxq���4�������|^d��!|Z��+b�����yZ��r+�o�Il�X�w��R�o��S�NUU��~Z' j����$�)>�������hB6������?yN��.��b?/���)���+Y"�'��&�x��E�	m���W6:�C��2�����s����	���3E�ϧ�O%7�a������u������Sק�#m�T	�JY��M�O_c1Ϣ�3��7�Ğ�frzݢW��W��(�{�5�1���8��a���ȧ$ZT�d�Cn���;���e���K�kπ��F�Tuz��z�׺
3�����=�pR�z�N9
ᲨS��\bc�n^�02�$��9���bW�����{*i�1��)��^sRֵ6�� �?��{I�R��72d�<v�}�$W���^q��6�RW�C;UR܃���ŏ޾���Νh���x^�x��m��j(��I\,;J�Kv6]dŸ}�R�wx5#�59GrL����ᧇ�Q&+t<��}�Ŵ=u�H�
����;ФTH
�(�Z��o>��[�*��[�Fb�|��m�w�ݏ���8K-C���k�H�]ы�?��;1��Sݲ�l�s�l)�	�y�����B��U�\>��U��d����;�~��LW-�����V���ǥ/��+��-17_�6�I�%��K�8��D\�d><�;��d�^��k,6Ik���̥$Lf�;��%�9Z��h�@+�%�l���S��%� �!�,�T\R�a(v��1�l׼
e2m9A�hA�׿�nYl1�iU��@lyr2;uO��e3�>���2
f�SL�������[5a9N�հ��:��l6�ݙ,���b+)hC.؁�dǯ�XJ[�:+���#�/,8�3w��
Ӳ�=z9�+�YZ�dߓ�K��,{���){^����'Y_�93?B��K����W�1Gi5#������kژR`*蓟�6Q����mX�x׵@iQ�!����@o�T��W���T�P���#Y?rU��{��:���LO�3�~ǯۏt[w=s~���eE�Q���U��p��.R¦Ji*
��*sz��7��m̫�n��5��R`ͧ�V�s�VD_����\����u�]�=_٥Rg øn�!##�u��]D�Z])F^�,O-d��'��'�CtB�
���|
w��3�YC7N�KEPn^����;7��� ��ֈ�Ҍ�>7��9'��;/�V�鮭4Y> s��9��m�&��M�3�K7������!& ���J���Gsz����x^jʢ�TE*@(HFV֚ި"��֕�
[&�P��Er�,d=�vs��5��_�_ɽe2x�@s!�+<g�D���YSVw�YY�2y��vh�D�g����,�a�wKN�䦛1�fuÃ��h^4#��K��*��W���kծ@�OR,�t:Dp���c5�jm��iZv��l4N��H��F��J>�B��������"��:2'�?m�y�N���]-W�Kd��u��/�4el2��|zZo#��ԓ�/�x�N�I��<{�]s�G`.�ꈁ�g���R��-JTp2�ŊLSjN�F�,�@y^ʰΓ�+��)�(+��V*��V.����f��f2IXs�9�J앢��U��s����{�|��N�Cz2�o�pS�,D[�p�q�s!@���ݸ��[�"z&��7j�)d���$}!�U�g�wk6ǒ��Ջ�q��Y&ܥ��s�"s�B#�&�R���p���M*�RVO�}�Ej��F��0�6ü�gV���7�i@5����e�éI���8�0
��! .*�00.%p��F&�ܻ�8_�t�ɍ7#JK��r�����r.9HDb��ѥ�q���b��ܹm���\Ɏ����(�Zm��z�%i�sZ�+�h.��e�U_O_<Sa�e-�-k$%SJ��{�l7��DJ*�m�j�ٱ�T�2���"j*o����u�5���N�ry��\&_���7�5�p��u(T�S�f�s���tFb~|v������(lԧ�jE4�t�*�a!�f��o�3��~x�>���͉�k��3&L���_#����c��P�Z��v�c4�Y� T��4�.;���	�9�:.��%Y�S9Y4ƙ-�����Z�f������XmS�	��cؽ���$�Z%M>3�i�X�����ˉݝa�/HI���ܷ}����K�W�^c/���1d�x�5S��v���ӯ̋���R\~]-^V�sGt�>��w�VΑ��͗f=��Z��)bi0�����%�_�Z��_�ӻ&Ԅ�!?~{��C'��F�2����2��� �j��O��a�������Õ{�'�(�,.���h)���z�ń$N]��Z>�ӣ)�vZ���Ta�]���K����Ӆ�,.�5�+��F*�V�i����^���D�{�źA-��4^�V�ɱ��i���u9�Z[�,����\S�Sr�z��IJ�irp�Az�g$��ÓS��a|x����q>�����\A��="�:��?��V�JԠ�<�Q�?Nf��{�z��/�J��_ݴM�<|��焈��C���əd���]�U�)�ͭ�f6*����=��H��!"��NQ_�QOי����!�@oٲ���}�:�o�ح��TY_\��m�����/eߕ��.�)��x����W�HQ��D\L�S�.��-x�� �$�zFcx��v�j�Z\�9؃�ˎwl_�GN�㓿~�|�p�$�Wց�5{k�9n�)^��.?N(�.��jE1+�rqJ��W�\��X�!�qт'��̴�I1��X�a �϶��ƚ���<�{���l���.eEЫ�26�$���M�06���Ef����4,�^	��9[�<n��ph�ϴ���q9�e7)��F�����>�Q>�@��%�lV&����m�wY�z<��?���6y�'��Ғ�l��ہ�Z�x�h�T	��i�JA������G1Q�K=�{U��(���S����摈��xb��N�A9�An2����.���Q��J�p�nΧq�l^If��&�aP��������)�*%����z*y��U<�S�����D��g��7�'Ŀ��wH��9~%)3n���>@���!|*�b�����Rɪz+m]�u�oX�͢dg�9
��ɴ4U��3o��q���b+o��?�SgT�����;�U��U�l���|�R	��F���g��:]d
�%��u{�(����X���S�+�|�ӼN8��B��uY~%(@:$�J��aױ�Z"�nf�Γ����I��rh��:���$4���n��#�j���G�4\dFo�y��{���瓹�g�h���|'�v8?����>�+���l��w���8��}���B]:I3��'n4��wt�$��Q�Ei<kB��?�Q�Z�Wf�G�R�3gΨ����$cQaϞ=�3L��9��I�802xUI���#����عs4Z�ѣ��Xy�ahh###س{��L?�s��7���KL�="3qH)�¹�'�k�n�`��S��!a��c��#.�G��~��Ql޼I������[��>zz�s�ކ@dG�0$ݕ:�plժUH6���i�W�'��������v������H�rE�,g��d�3պ�F]�\U��_8��;Z�q�ļc����?���҂�p�8�Mblﮝr�V)�{�Cx� ��G �{l��رCt
Ssgg'�ڌ�a�o�N.z�Ĵ5s� Q��a����s�Vy������m-�p�uw�]������{��O��@%D�%�}JU΂������~��I���|�����q��]{�����r\�mo�MB(1��H�'��G�]�h&ഋ#���R����6~�ͣ�Ik��U�ں�����T�E~�JWl���׏�FQ5ۙ�1v�EK�l�ѶM_TLf?��Y�0�$����[�_b[2��z_����zm^����Z�S�@c������C@z�����`�l>Dc�*��֧m�ζC"V�����2��h������D!G3y��A2>�� %��ۺ�_��$LO��K7�Z�'����B��j~�D�c-#��"�ʹ�	/��;v�s��O�����m^!�:��b�+�&i�_�%x�� �48��4    IEND�B`�PK
     `+�[x^��_� _� /   images/d5d3b89f-59ab-4c38-95f7-2948dd30f8f5.png�PNG

   IHDR  �  �   �Zd   	pHYs  ��  ��"篻   tEXtSoftware www.inkscape.org��<    IDATx���wxTU�?����LH�$X%B4���4E�"(*(�O���,�����HY��
X@A��6��,Xhb �d`���"�������8��I$7Sޯ��qιg�O�p9�{�0�LDDDDDDD>�h4��; P�; """""""b�NDDDDDD����&�DDDDDDDn�	:�`�NDDDDDD����&�DDDDDDDn�	:�`�NDDDDDD����&�DDDDDDDn�	:�`�NDDDDDD����&�DDDDDDDn�	:�`�NDDDDDD����&�DDDDDDDn�	:�`�NDDDDDD����&�DDDDDDDn�	:�`�NDDDDDD����&�DDDDDDDn�	:�`�NDDDDDD����&�DDDDDDDn�	:�`�NDDDDDD����&�DDDDDDDn����� 44M�4A�z�P�Nԭ[!!!P��� "?? ������t��s����ٳ��ή������ȭ��� 44�7FHHBBBP�n] �����w5���Ɂ�jEqq1�\�b�_�x�Νùs�P\\\�?y&�n$   ��~;Z�j���DDD�y��hذa�~����:u
�Fjj*RSSq��&�DDDD�S�ի�֭[���-[�D�f�P�f�J����8v옽�m���j���C�A�L&Y�A���� �o�w�ubbbp�w�h4VK,����ѣHLLDbb"v�څ˗/WK,DDDDDU!44;vD\\bbbмy�j�%77����HHH��}�PTTTm��2��hLHHp���L�u��ݻ�K�.�������<�����رc�n݊�����uQmڴA׮]ѥK�v�m��K������_�}�vlݺ�.]��|tӸqc<����ի����;�r��Il޼7nđ#G�;"""""�bccѫW/��ٳҗ��AUU$$$`ӦM�����Q�!y5&�>@Q�{�x���q�=�@Q�f����<��0���7��
)))X�v-6mڄ���*�>DDDDD��}����ǭ��Ze�'33ө.   U��


�e��]�{�L�*t/V�V-0 O>�$7n|S_+--���8u�Μ9�3g���]��{�V�fMԩS���C���ѴiS����iӦhٲ%��� ���������W_aժU8{��""""���C��w��7�|�j��ĉ8z�(Μ9�ӧO�ܹsHKK���m�%iQu�Ա��~�-� ,,aaa��ߎ:u��p| ���c�ʕX�~=


n�kџ��{�F��o���뇠���~ff&���`6�����C�!==�
"�S͚5ѲeKDEE!66���7�P�j��~���C�UA�DDDDD%�o�#F�@ǎoh���ɓHJJBRR��ߏ�G�����
"�S�ƍѪU+DGG#66&��~\���|�2>��s�Z�
YYYU�oa��E�ׯ��#G�'���i-���l6c���ؾ};<��U�5k�.]���{�A�v��g�R�~��ￏ�G�Va�DDDD������Ϣ}�������,�ڵ;v����ۑ��VEV��`@ll,�t�Ν;�U�V���!33+V���U����S��z7&�^ 00#F���a�P�F�
�Ƕ���͛��?�ʕ+y[.�C �8.�<.��$��d�Z/�Q��\)�B�!BTUm �h�������H �+�3v���z�B�.]*�����u����w�u�y����/x饗p��V�=YYYضm���{�ڵ���y�%)����B�pAU�K��dJ)���
!� ԔR֗Rֿ��n!�l!��@�r�߇���W�^�ի��
�����X�x1�����~��{0!z��	& 44�B�p�֯_�իW��V;_J� ��!�HB$�~��GW�^]�����ZG	!���n�����ĀY����˗cٲe\#CDDDD7�V�Zx����SOUx����f��_���u� Ҥ����`�Z-8W	a�жm[����� ���� ��s���͛�_�~�ׯ�֭[��s��q����_~���}tռysL�6w�uW�����X�r%�o�UU��H!��wR�M���X,U��Ņ�8�FQ�^ z����6**
O=�z��	??����'ObڴiHHH�ܠ����ȫ=���x��WQ�^�r�����o���U�p��	W��?	!6+��}RR��J�:����p�ު��BDh�3��ѣ��֭[W�koڴ	s���Y����>�G�.w����شi�/_��j5� � X-��"%%�T�|�ڴiӰ����' ��d�I�&<x0X�4)%֮]����#;;�j�&""""�иqcL�<]�v-�mzz:V�\�/����&�� �B|QPP�����n����d�0P1���v��x�:u*��edd >>�~�m%G�}��{���P̞=qqqe��R��ƢE�\%� ��`0,MLLL��X�J�6mB����	!F hY�zݺu1l�0<���ϟ�믿��~����%""""֣GL�2��#�rrr���K�.u5 ��c ����\�͟�Ett�] ��$4���������w�]��ڹs'&O���/V~�^�	���ׯ^y�r�Mۻw/�Ν����Z�B̷Z�_V����"�111=�V�x!DO %����[��/�w��e�>��*���cѢEݨ������\pp0^{�5��۷�v��������"33��b-�f��ת�U/1115UU`���N�:a�ĉ�����:/^��ɓ�s�Ϊ
գ1Aws5j��o�Q���ܹs�7o6oެuy�����?WE��-66�NUU_��Pj�{LL^}�U�y�e~���$���K�靈���ǵl�������l��/� >>Ǐ/})_񑪪o��қ!�PL&S_ ��u�f00p�@<�쳨]��AMRJ,]��-r�?��b��ƚ4i���痙\��Sϛ7��A!�6�����b�Qձ������ ��j�n6W�����/�\��+W�`ҤI��W��IDDDD7��ěo����@�m._��y��aݺu�/����o��}��<.�!��dz�t ю��ׯ�	&�;���o�a�ĉ�|�rF�Y����v��a���e�w9q�&O���\�^J�*�x=99�����]['3@��)�����o�}��.�[\\�Y�fa�ڵU%�!ƍ���~��v7n�[o����UU_�X,�,H7%����C��s ��x�����o�����|��ӧ��s������P=t7ԫW/̜9��M�֭[�Y�f!77ױ:GJ95  �]w��V'���W!�;p�Q!0h� �?�̳+W�Z���xN�!"""�rF�ӧOG�>}\������ٳ�F���:�b�l�� =@DDD��)R��p�zݺu1}��2w����Ą	�g�=BukL���ȑ#���ϻ��,;;�'O�֭[K_��`0<�i��W��m��)**�.�|�b������o��f͚�|�M���믣��-�~Q%�U�.\X�)I��ɘ4iΞ-1k������iǎ˯�8=ITTT��(K �����&L� ��a�������
�-1Aw#cǎ��ѣ]^?v�Ə_z�G����?���<Ytttw ���ꂃ�1s�L���.���/�`	(((�� ����H7�k��|���(�m֬Y�ٳg��ٯ��S�%�ʃ�Pݺu�t�� ��a���;�����ѤI��I)��[o��>�)R���!��+�`РA.�lٲ�'O.=����r`JJJr������)����:EQ���b�ȑ.g-�ٳ�?�<����
������P��d��G�c�̙���/��������W9j^1��>��VנA,X� 111��Rb�ܹX�j�NQ�&�n`	>|���.�C�1�#2�:>o=
�{ ��y�L�:�唛��D�=�I:���[�.�-[�29�����/��;J��%�a6�������i$�\	����h4bƌ�ݻ���͛7�|�!�wJЕ�x�^x�er��*fΜ�9s�8&�yRʑ�����ߘ��䏤�� �}��3f���5����~�eODDDD�v�����]&��ϟ�SO=U:9߯(J[&�7�l6_hݺu!ě T (,,�k��Vf>a����O�0I�ύ��9�ƍӼf�Z1y�dlذ�^'��(�|�W�5�jmڴ	-..^���.**
������6oތI�&qww""""S�F|���0�L��O�:�g�y��fp[�F��111J)W�e�5j�{�9����bҤIؼy�^!V;��W�>}����׼VTT��'�H����k����۷�laa�} 6��,F��K�.i��gϞ?~�NQePs��q��;v���J$�Rʥ���������M��> ༭>B||<�t�U�f�*s�}�:>���i�ӧO�ܔLUU����زe�c�>���511�^1���f�n��a)�
[]jj*�y����k�gذax��'u������n�ĉѭ[7�k'O��ȑ#q����9)))�l۶�X� }��b��`0t`?�j�ʕ�;w�f��� ��_�B����
���=44���F��5[r�i�}@B�F�������z��KV�^m���!�\j�;r�H�k�_y�t��A�������<��<x�浳g��g�AZZ�c�����Wu	�G%&&WU���2�V�j�*������CBB��{�!88X��� ,X� !!!��gϞ]z����� ��T�իW[-�( Klu���Ǹq�PXX��^Q̝;���DDDDT�L&^}U;�NOOǨQ�p��9{���L��a�XN�n �����}�ǫ�h�3f�py42U>�O��x�DFFj^��O���Ǳꈢ(}-��.U:)�LII��lu			�2e�暘��̛7z�IDDDDP�^=̟?_s�jAA^x��<yұzfJJ�l�$$%%�QU��?lu���ضm�f�x #F��+<���	z߾}��#�h^۲e,X�Xu������l����2RJ�~��Ä�mu7nĢE�4�GEE��_�->""""*��f�B�ƍ��I)��o 11ѱ�����7t��,�UU���.�}�W��~���=�bcc��gym���^{M�����1e��c�2TU}���'t�Jضm[����_��{luK�,qy�àA�p����mРA�ܹ�浏?��ĞO 6�nݚ��T#����Q  ��������ʕ+NmfϞ���:��]Q����l�7�q#�|UU�X,f]�$'			����� ��>i�6m�;��V�iӦ�nݺz�IDDDD��v�m.g8�޽.t��+����ի��G.��� F � p��yL�4�q Ӯ�P�<^��2����S��������r<�9w���;���# �T&L������4p�	�CQ̘1Cs������	�%�����l��5Hr)99�� ��V���_�x�bͶ}��E׮]�
�'y]��1c�h^�ꫯ��?8V}����.�Q�Y,�$ /��G�����5������w�N�QiC�ATT�S��S�NEzz���*����x\���|F�q�]��ҥK��o�i��2e
��W!�KЧM���� ���'ObΜ9�UG���F�]����% >��?��s���O�m_{�5ԬYS�Ј���蚰�0�;V�ڧ�~��۷��B��)))�Q�JHH(B�\�4�7�@VV�Sۆbܸqz��3�*A�ի:t��T/����ӑ��k�*B�5555S� 麨����2��;|��7����+kҤ	F��""""�M�4	���N�'N����k/!v�j��-=c��c6��	!���z��g�b޼y�m�;�C��|��$�?^{#�/��{��q�z�l6��%0�a�%[J�7 V �x�b������p=�#"""�i�۷G�nݜ꥔�1c��B� �pS8�g6����u��W_a���N�E�+��!�����IЇ���P��.��w�q��)%%E��mr;�e������/�������ߟg��Ė�iY�fM���If���XrKF�� G��[fΜ��as\\�w�wx^�+����1B�ڂ�T+ 0ZJ)���n���� �Wo�f͂��� �{���;<""""�ӷo_DDD8�gff���s�ڝ���D���%$$䪪��Mu?y�$V�X����^��`�3<��	����5wLNN�ƍ�e!�����z�F7/!!!���ѣG�v�ZͶ�>��^a�$???���׼�x�b�]���#��·j�[�X,� ����,Y����;���?�gh^���z����'�Լ���c����gu��KNN�`���h�"Ǚv;v�]wݥghDDDD>��CӦM��?�իW;V-LII��n�Q�RUu"�, ����5ۍ=~~~z���<>A2d��Α?���f��,�|�رc�z�F�K��" �r�
V�\��nԨQz�EDDD�3E��O?�ym���(..����:K����Y,�� ����ׯ�����.,,���ȣ���@<���N�RJ,ZTb�])))_�U	��|HJi_ôr�Jddd8��ر#Z�n�klDDDD��G�s�?z�(6o��s!�t��rY�ب��p�z6�|��n�С�ѽ�xt�ޯ_?���8�oݺ���\�qQձZ�3�@vv��+��gXDDDD>a�С���/��ڗ���Y�懺EUf�Νy f�ʛ7oƑ#G�ڵl��:u�34��	��Ҽ��'�82����%(�r8`���z�j���:��ݻ76l�ghDDDD^-::&�ɩ�ԩS��Kt��y-�#/�����I��(����5�q��rxl�~��w#<<ܩ>))	III���(���GSe�B ����W_}������<�ޡy�h֯X��q��|VV�R͆�RSS��Ͷ7n܈?��é]ǎѬY3]c�F�����_���O?u,Z�f�f͆䱒���!�c+�Z�������s-Q%FϞ=��333���:V-���^i)�K P\\����?N�x��G����xd��x���ҥKغu�c�|�p�y�wl/N�>�ݻw;5h֬ڵk�kPDDDDިO�>�''mذyy����B�=�Bf�9�L���k���{�1(�G��n�#��������N��|�M�����?�50ҍ�l�'��a+�]�V�]�>}t������[=��C���K����f��b"}]{���ŋ��O?9�iԨڶm�wh^�c�Ҥ����?ORB����MU�e��?��#�\���������qy�F�!&&Ʃ�b��89IQ�=�bf�� �n�����^�z��W��A��Oe��ߏ�'O�˪�~�g\�?)�j Y PTT�~���M�:uСC�C#"""�={�Ԝ��a��������E�e���Ν;5�z�����kP������O��ys���,)))ɺE��b�dK)����{�vݻw�-&""""os���;թ�Zzpd%�~�~����qm��j����������.�C���w��ũNJY:Aw�V����(kl���݋�/:��ԩ��1y���`���:՛�f\�Pb���F�u�-!�o��j��s��z��u<*A���C����>��g���B�/􌋪Onn�f ��'����S�[n���v�ޡy��;j����?:S���:5"�$�Xm{������l�6L�o�G%�qqqv�߱þ�7���f����qQ�IMM-Bl���o�^��5󂈈����*�*���F�`�-���o�\=��_uj����W��Ֆ��FM7��)�}nͮ]�4�d�:"""��Շ��?p��{YU�MN��k%$$���Vv,�B��}�<*A�:ޡ�� ����(
o>FQ�� $ dgg�8��&66B�C#"s���    IDAT""�X!!!w����_�\zÆ��P���s.�t �{P�<&AW���N��EEE�������y����3 �Y��}��ڄ���E�:FEDDD�����48����?o۶�y�"y5!�O�קN�BZZ�S���8]c����h�Bs�y������Y�EnC�����g��d2������Ҭ7�͎E���V�Z�d�ʥ> ��o�z��<&A����5�SRR�;5��SUu�����YU�V�)''G��������[�z��}n��c�����n��'��ذ}�.���Q�~�HKKÕ+W�ڸ��3��Sjj*TU�������(!D����Ç5�p���yL���	^��ϝݐO���?��VNMMuj�Q��I�&N���XG���M��>�Y����}#<&A��A�ȑ#�;Hgff�5(r			E ��)�n4@͚5������#���knW����Ԁ|���hZZ��ӝ�4o�\ט��G$�B�'x'O����R;v�X��q�{�R>}��f���P��!"""�T��L�N�r,rṗ���`��K}6 ��}#<"AoРjԨ�T_jz�qC"7�(�1��3g�h��M�����|M�6լw�8�و|µ��N�V�;,,Lϐ��G$��r�f��s���A�8)�	�kW	:oDDDD���K)K$�R��:�D���V�;((!!!z���<"A�W��f���Xt�SA>EQ���.\�l��DDDDD��3edd����^B�tjD>Ea c��rxt�^�(�4]�!wf�+dff�j�:5�<"""��խ[ש��&`B�?��O�R�s0�c�����G$�~��7	!�E��!�T\\|��ZJ���L�6�A�O��T*+0��9�DnIa�gddh��z�C�yD��YY���z�C��`0\r,k�P�V-��!"""�TZ}�R��{�����V�`��zyD����Y��`0�����������B�6F�Q�x����<�V�۱����)������\�r��ct)%����e!��'�|��R(��������ADDDT>�>S���� ��6�t�]�MЋ��q5��M��rn�A�����c B{�[kp� ���]Qn���bYn#���E�8DDDDDT������wEr9��G$�ZOc���JW��@���h��'{DDDD�'ǥ�6��o)%��)e�}o���w��	��t�ι�8|*�v�����4T`/&�������^��@@���E	�+rO�:u
`�C���O�����ʧ�gr�{�-r[B{�j�	���=;;[��v����R��z�C�)''��g $$ĩMVV�n�y*���c� ��)e��:u�h�a���xD����{�LQ�$|��j�������DDDDD��3���6{�|�����[��f�+W���7����/��&��jC��!�d0�O�����6d�NDDDTZ}��	Xff&��>�"#��_�H�]�R6,qOh�K0�TUmn{]�a�'xDDDD���3թS��F`�S�텫�7���	��s�4����쯅�5��B���v�l8r�Y""""�?�?ީNQ4i�ı�Bǐ�=���B��]PP�˗/������;I:� ��� �T��̙3:ECDDD�\��BCC��^�{�u�������ٰ9s���z���<"AWUU�)^�f%f�DDDD85"�!�����iӦ�mΞ=�[<DDDD����Ӛ���o)�z�C���ŋ �k����{_?�H��ԩSNu-[�t,�ըQ��n�[B( "m�R� W׿dff��Gr����c�t	�ܒ"��:$$Ds�ɓ'u��xL�����TW�N4n�ر*Z��ȭ���� �V���۝�>|Xϐ����<Vzz:��Ҝ�K��ZEEEu�܍=A��{�9�ͣt��AQ�vz�C��n��u�A�Nm�9�kLDDDD�Lkp#""B[����/Vנȝ�������l���yL��j��d�sf����^�۱��'R�ADDDTqZ}�ڵk#<�~���>J\}Jc s��lTU� ���ȑ#���u���-��.�S�N��EnCa�ǡ�g�.%%E�x����<��bѬ/��b��bbb� P�V���sjs��1�����1	��j�����꣣�a0lE����.�F�.22�>�[�M�6Nm���������:$&&j�;&�R���Üw�V��~��F��>� �o�>]c���@RR�S]PP"#�wCQ�^z�D��h4����r`` ���6f������JKK�<&�]��>5����:t#���\w�}�f�܍��Q	�޽{5����k)%t#��i{ݮ];8�q��!""""״�P���%֡�������sW[�s�Κ�8�~c<.A���w��ҥĬ����(�C��+8� �![��g�n�Νz�DDDD�5\��J���%r��t|�5:t����ĉ8s�ޡy�J�

4���y睨_����(��z�E��СC]4 !D��6�/_�����������ܹSs�����X��Ԉ�����ѨW��S��۷��7���e+��=z8V=�Ԉ������uTT����ر��ω���n��+Wp�������11�����Q�h۶�?�Gm�^��W7�رC�����%����!�t�/��hk2�"��W���2
!�	��Ķm�t�������lݺթ�`0����yCJ���1Q�(,,���9H
���I����ޡy�K�ϟ?�y�u\\7n�X�7݂�j�(ʣ ^{��={:�����/���whDDDD^���׬���wEEEq7w�gϱڴi�F�95ضm


tʛx\�h�$E����g[@1���^�Dǎq�-�85���y� """�	�N�Ҝ�ޮ]���+�2BϸH_&��1�>�r�~�4�mڴI����G&�7o�\Sܿ(��Gj\TTĵ�^*...�}N��k��������x����EDD��-(ҕ�� ��V�Z��W��ӱ{�n�C�*�������Ņ���cǎ����%=�"�X��p��۠A�w�}Nm��Ҹ�$Q%X�n�����}�Q���'�֮Q��p=�"}DDD c+?���pj�~�z��	U�G&� ��_j�2ıxWTTTg]"�DEE�0�V~��'������믿��j�12""""�t��e���N�6,�]1n���C#ԨQc0�[��K���n�ڵz��<6A�駟����T߱cGDDD�ˊ���g\T�Ey@M ����ڨ�����J�Ј����֚5k4��X������% ����B�I�����_b��ٌ�G���7���j����?w�B`ذa�U�cbb:�U���� �l�����N�:N�~��'�>}Z�Ј������ݻ5�V�Z�^f:�[�n���#:th0�V�����5ۭZ�J�����&� �z�j���:�?���hѢ��,�|Sǰ�
Y�֗ � @@@������������H)�r�J�kc�ؗ'Cq���'����N۶m�UU�l+w�����N�Ξ=�~�A�ؼ�G'����o��E��Q��z����rjH%666�x[y���hܸ�S;�ł��D=C#"""�	�ׯ�\f�Ν���I�϶m��U�����B���c�j�[�b�~�$��WGJ�v
�ӧn��6{YU��j��TU}�֞׬Y#Fh������(,,t9�����;yܴ��h�fC����uL����~�L&�v�.]r��7]?�O�Ϟ=����(x��W�"/_�<ʩ!y�������G�����;�ۿ?~��g=C#"""�)�}���(�w܁�z�^�R�rm$y !�4!D ��������[�.]���|]c�f��WGL

����nt���^�R��M��t���OJ�>�}^�6m���zJ��{�)�������,[�L�ڄ	l+֒R~�[`TiL&S[)島�SO=��͛;�KKKs��?��H������g�i^�8q"l��V��_�F��ҥK/���'M���;�۳gv�ܩghDDDD>i͚58s�S}���1r�H{YJ���d�glts���! p���g�yF��E�4J��yE�\E�x�S}xxx����L&���!L&S$���r���q�}�9�SUs���12""""�UPP�y��i^6l"##�e!Ģ�m�6�+6�9�z@[���^s�aw��A|���z���&A�����E�4��1�[����DEE��ݘ�m��!> ������[�f>�gxDDDD>m˖-ؽ{�S��`��o�	??���M
��ݐ���6RJ��p��{/�w��v�ܹPUU��|��$� ��W_�b�8��n�����EQ�	!����6���3���_y�4j�ȩ]zz:.\�ghDDDD >>���N��[������3�L�G�[����)��? F 		�ԩS5�nܸ			z��3�*AUUӦMӼIDFF��g�u�z�d2i�ڙL���l+w���>��f���x����]�����˗k^{��gK�%�X�F�1U;UUhe+O�<6tj������x=C�)^����Ç]�$�����;VM����G\Tqqqq-��q��٤IL�6M��Ν;�n�:��#"""�>��C?~ܩ�`0`���

�UՐR����t>+����d'�j+0 ={��l�K�.�����z�8z��S��(x뭷�) V��ĴrjLբu�ֵ�V�7 ���h��o��ڵk;��������������`�ԩ�����K�����_1p�@�^�Q�L&�}B��xdd$&M���v����b^��`�ĉ�[�7h� ,p\�^OJ�]LL���f�������� D��&M�Tbj��Y�f��ٳz�GDT��F#a4������`0���(^�O6y���D,]�T�ڃ>�!C�8V�9x����Fe���n-���֝׮]����<��ʕ+�2e
��z��S��d����Æ�K/��ym��՘9s�c������;w���%8r��������w9�}Æx��t����� +�R"!VB��u|�^�@! �p�^ßF~~~�m*BJi� ��j/;�QUV���ŰZ��Z�(**Bqq1�����*�����"�Jc0�b�
�����b�={���I)_NII�>���\LLL#)�. �W�-B�N���J)�������;L]�FcBBBQu�xy��(
�}�]�{ｚ��~�m�X�±ꇼ�������C�T�bbb�)��g�:t��ŋ��;q��|�Idgg�#�?!���`0��k{mK�m���$�f�L�^�lI~餾��EEE(,,���:DT��M����?�\������C�����UI ����?�3Fڶm[���p+�;�2e
�x�	��+W���ᘠ�v�����ЬY3�k����_Ɩ-[���_���m۶9oOU"::z<���r˖-�b�
;��������q��=C$�jfK�������???{�1	��i�_/UU�#�EEE�$>??(**��<���{��{�iޓϞ=���;n2�
!�2�͟��k۶mPAA��B�.��#F��_�l�w�^<��3�'ey&�:kժV�\�5j8]+((���?�ݻw;V���7�#�U/::� o��M�6�'�|�y�puM��M��
��tb0����Ѩ��kͦ�t���W���>_\\������#77L�����ѣ1v�X�k���O?���L[�U��l�D� }T۶m�m�Rv�����S�N��7)--��_q��E]���jеkW��_��|�����1c�`�޽���?�5�U'&&f���~}�F���'� ,,L��G}���U.[��� ؓrO��,ޞ��ǖ��F�

������|�E��n����?��Ci^OII��Q����c�R�7���;��M����'��Na?w�{��/�G�MAA�~�i$''�gu`�^M��4.;;cǎERR�c�O����X,�u	�Gt����ҥK�!\�ƍ�d��h�B�=7n�k���"7�(
�F#jԨ�+�/'�Z|=A/�-y�M����Evv6w"��>�qqq����ۇ�{�q_!	����9z��+bbb�"��  �VףG̙3Gs����?~<�mۦg�Ն	z5��?����������\�7��� �(��PRR�a]�rQQQ���3)�ö�f͚ᣏ>r9r����ѣG���P�8��l�S�m��q�&��϶���{vv�汪D�BBB�駟"<<\��b��1c����X��h4�v������ƶWU�[ �mu�<��O��rۜ9s�j�*�B�vLЫ��(�1c���y�v���?��X�&�����曨BL&�m��Y��s�>���s�łQ�Fq�v�j"�@@@�}T<   5j�М
Gׇ	z�Z�(((@^^rrr�����y�&M�����7BCC5�>|cƌAZZ�c����dBB�w/~�b��у ,h�<x0&M���ߠ����[��3A�f��୷�>�y]UU��Ǘ~jdB�LNN~Sr��u3�L	!V�k��С�ϟ��[; 9r#F�@zz�^a�4��`�%䁁�L"�����*��������v�j֬Y3,_���LZZ�}�Y<xб��b��lޭ�&r�ڒҙ ^��	!0z�h�3���V�Z�9s|o�t7��s��p���O?��o�]��ׯ�F�3|�W1QQQFEQf ���}�����믻ܙ955�F�r<���*��(D�5�8=]_LЫ��Ҿ�=++����Z���O���[�d��Izvv6^~�e�ܹӱ�@J9�b�,� Y�\[o�
@G[]PPf͚Un��{>1Aw��`���x�G\�ٻw/&N�X�h�?��O���l�� =Xtttk � ����F�?�v��`���9'�D��5j ((L�t��8Ҟ�������牨����bɒ%h֬��u)%�����w�-��p��(Ó��������� �# !����p,X� .߷l�2���;:D螘��EQ���c��.ۜ?/��RRR�%���x%99�J��Qڶm�_XX8�T8�wiҤ	�͛���(��MHH��q���&���#00��9A��ݽY�V���#''��ϯ��-�܂?���_\�ٺu+�x�dee9V_B��������%�L�fB�� J�<>���1c��%�RJ,X� ˗/�!J���<'Nt����j�G}�?���Ӽ�R�SRR��K�n.&&����C8l\=cq�ԩ�S����n޼���:�]'[B��5kr���`��YlS�sssq�������4P��R�vm,X� �ڵs�������?�����җ�*�2��,4���{V1@-[}@@ ^|�E4��5����:u*6l�`&�n�w�ޘ1c�F��6�����ɓq���җv������*ctW���a��N0��)G�Z�0i�$<��e�ɒ%X�p!;;D`4��xPPwT�PL�=��EEE��͵�e�x��c41}�t����eUU�l�2|�����-�o�������r>J��y睘5kn��V������/��}��Uu��	����Ă\\=�mٲeX�dI�#\T)� ������X�ATTT=!�KB�9^�ڵ+&O��ƍ�x�ճ�M��M�6Uu�D+((AAA�i�f��ga��}
����+W����KD.!0h� ���K.7��'Ob���سgO�K� ��h4~����[�������6R� J<���1c0|��2�
�	p�ԩ��c0Awsu��E||<ڷo_f�`���0�ͥ/X)��孉zddd}��P��ZӦM1q�Dt�̯֭q��	�?G���H�<���?j֬i�Ä�;1A�n����\�r999��[k߾=���Q�n]�mTUŗ_~���{W�8mu^1����#oMԣ���0@_8�� ݺuäI�V��X�n�O��%��0A� �����;F�U��Q)%���;,X� ��G���b2    IDAT�b���_���[�4`��L��E'�|@M�k5k��ȑ#1dȐ2�	 ��0k�,nG���Z``�=!�r��ݷH)QPP���l\�t��T]"ШQ#���,w�,++|�>��ҳY C񉪪o���x��B�L��/H)B�ļe˖�4i:t�P�����Ü9s��_Ve��	�����[o�����2��o���ŋK�f�`�U���{DDD@�5B� �ḱ��}�>�(Ǝ�������1{�l�[��
#&ro�� ((���

*��y'&�ͶK��+W������D�ئ�O�0���gϞ�ҥK��W_�j���\�[ �Z�n�y���N�Ylll��r���o Z����#G�_�~��E��~���8q�DU���{���`�?O<�D�����\|������O]%�� �K)�Pe��lv�9oݺu�x�b7!� � P�t���@���#F�@Æ���;w�����q���*��Ƚ٦�ےrN['&�䨰���ٸx�"��hݺ5�|�MDFF������X�d	���;�u 8`�����_��������~~~� ���)�ǈ#��#���f�z_��㏵�͢R��{�6m�`ڴihѢE�m�a��X�G��\���!����~_���cbbI){!z���[�9ްaC<��0`@�Ǧ٤��c�ܹX�~}��L����5k�F���&�䊪����222x�	�,����C�b�ر(����U�Va͚5e-�<%�ؠ����������fVj���d2E�)���> �Yw\\��nݺU�!bb"�|�M������b���0d��9AAA�W���Y��7o.��q ; �R�Z�V��;w�̻���u���/--�v���VJ�	@g w���uEQйsg���]�v-��p���f�,\������!???�(97w��0A����������/jM�%�zM�6ń	н{�
������͛�v�Z$&&�մXJ��. ;�X,Ǥ�U��$""�v@@�I�A�@G ��j_�vm������GDDD���ŋ��{��o��ҙ���4l�/��~��
w³���u�V|���صkWE��X���!, �I)�8�(�EEQ.]ڿ��M�m۶u�Vk����B�� �	!Z���!D$�H e.|B ::�z�BϞ=ѨQ�
�� �g�̙3���~�'���Gpp�=)'�(&�t#������ũ��ڷo��'�U�V~ω'�i�&lڴ��Y��r B�Rp\JyZJ�&��TTT�~��A�s�u�旑�Q�j��SU�>��B�B�Rʖ�:֢�o��]��W�^�ҥK�f Wg�Z�
K�,�&�7�	�����رcq���_WG+##;w����۱c�\�|�fC)`pS�h���p��w�s�θ�{ФI��zrr2-Z�]�v�LDn�h4�V�Z�Y�f�g����n��jEVV��Ґ��_���BQ���cƌ�вSG���;~���ر����rq��}SS�BCCѥKt��:t��eq�����믱d��;w�f��iLнPdd$F�U�u!�TU�ѣG������$��f�>}Z�5g6DTT����;��xJJJ�ҥK������;���,�|�sj_O�K��3=3����(�"|�B 1�D��̦��(���DB
Q	EA�BD�%A��D�(`p@�oc�3�����3�/�Wu���~�:t��z���S�}I-�]g���t�}��}��B�D�F�6���]ש#Щ������8��}�{DGE<��#��G>����c��b��W^yW�^ŵk�p��d2�S�t/I�099���o~�q���:-��J��o~����Glll�B�Å}������ ~�w~��[RZ���}�6������lnn"� �N�Z=�׏(�p:���|�����Ν;����C�廮��h�?���_�׮]���!�E� �l6�n��n����q0��ii4����b��{rXQ���_��_�>���-o9�sE�Qܺu�n������;�+��F8�N��a��������q������d2����O<���&F�]`@N��<�ȱ�:G.�C&�A�\޷��`0�d2�f��(���D��o|_���92���`����鼫�$DGŀN���H����%����x�{ރw���p8}�F��t:�B��|>��a��j��`�,�0��}m��M������H�)`@2�.]�o��o��xǑ���\.���������˗/�+� ����g>����	�H���*�_�λ��5��mz�SSS��_�U��7������/~�WF�YF�?�0���wᡇ�ۣi���xꩧ��o~KKKZ�3�Ї�(�x�ߌ_��_������:o�M�x�<�~���駟f�����_���eh&��ʕ+�я~�z�	tҒ�b����Y���}N�r�N��f��?�����~��v�]��R���x�����~7o�Ժ����N ���1<��Cx���7��Xc�N����]���^z	�/_���|WՑ6�1�g�Y\�|?�я�:j���0�S��V�H�R��b�!GM�$�w�}x���7�	�.]:���Ǳ���k׮�ʕ+�|�2w�i��Z
����_��?��Ә��F(:�7p�dRm�q��-���+�s�0�a	�F7n���~�#<��s��B���kEA�TB<G:�ֺ�S'Ifff033����i��7���c~~��������/��@�#�����2��v��r��tB�e�t:H���
 (�J�T*P�L�T
�t�LF�D���ɮ�4�}mm?������+cS����zY��@.�C$aC*:��###�e.�.�K�&�I=۞�f�(
*�ʞ���x\}ｽ��Z���o��K�s�z\�R���2����.����r9<��s��w��s�DD' �"j���4�����D�(�� ���8i����Z���K/���}�{�v��<u�N������E�P@$A.�Ӻ,"��ĀND})�J��?�1�����XL�r�����b��3gP�ױ�����-�%"� t"�����W_����=���|SHD�I��3��R	�X��刈:������k�ԤR� �#��\.kZ�e2�066�p8�Uu"�b@'�}�k_Ӭ���j����f�������v��
loosj�11�QOivv����""�/�SSS��jH$�F�Z�DD�Љ�'8�NȲI��.���:@��!�����߫՞5LDԓЉHSV��,�n�k]
�A�t:�t:Q,������DD-0�Q�5���\.�F��!"�.2�����d2�H$�uIDD=����F����rA�e���u9DD�!�N���χT*���mv'��ǀND��h4��v��p@��!"�"�n7�n7r����yN���:������1iDDt$6�/^D�X���&
���%u:u� �Z��z�0�LZ�CDD}�l6��ٳ�T*�����Ύ�%u:uD����^�׺"" ��V������Z�DDt�Љ�DDQ�������r"":z��P�@ �x��߉h`1��]�$	.�n��ى��+DQ�����E2���֖�%u:�9iMEx�^x<�R)lmm��hh]щ1�ё�t:5�sT���6Y��N����	EQ�.���1�сt:�~?dY�9����P�A�+�DԏЉ��x<��������W̉��/� ��Y��J�����z��uYDDGƀND{��������O�Z�2�Q�in}w�\H�R��ND}���  �\������o~�bQ�r���Nl��fP'"�e�DC�T*ᩧ��7����y��!""�8Q��x�r����F��ND=��hH)��'�|_��ב�d�.�����5�{<�b1�b1�K""�C�t�oA �2�� W�4�����Hc�Z[[[H��Z�BD2�_|��u WЉ���fC �^�g8'"�����066�`0���5�""�1��Ʉ@  �٬u)DDD=G��cjj
�Bkkk�T*Z�DDC��h��|>��v�K!""�y�.\@6����g�Q�1� I��v��v�yƕ����v;fff�L&9������h�4�z<���u9DDD}Ku4[4e�w"�
t��p8������5Q����`0�ǃ��u�r9�K"��w�D}�d2����b�h]
�����8s�
�VVVP�մ.��:Q��$	�n�[�R������bQϧollh]t�>#dY����9s"""���n8�Nlnn"�Nk]t�>b�Z`0�.���h�I����1����T*i]�9t�>������9Ϝ���LOO#��buu�FC뒈�O1��0A��z9Ϝ���4�ooo#�Hh]�!t�e�����.�����HE��ax�^n{'�cc@'�1:�>�N�S�R����.�;w;;;X[[��(Z�DD}�����\.vg'""� ��t�n�cmm;;;Z�DD=����L&�A�L&�K!""�E(�XYYA�Zպ$"�Q�D�$	�.��M������l�ŋ�H$����u9DԃЉ4�t:���!I�֥Qy<8����X,j]�t�.��t�iNDD4��z=Ν;�L&���U��!���N�E��@���DDD��u���X[[C6�պ����#��w�w�.�����Kx��ǵ.c�1�u�^�G(��bѺ"""�1�$arr�\����vJB�x����k�\N�g9�"A �2Μ9�pNDDD��l������Ժ"�WЉN��hD(��4""":2Q1>>�B����e��u�K"�.�
:Q�	� �׋��I�s"""�+�333p�\Z�BD]�t�2���DDDtb� `ttn����DC�+�D \.Μ9�pNDDD�\M��t���t�b�v""":m� `||�\+++h4Z�DD��+�D'��DDD�M6�333p8Z�BD��+�DwA��!�f�i]
Q111�L&���U��9��{*���� (�����������x<�������k���������Ѻ��ǀNtLv��`�$i]
1�Ӊ��Y,//�P(h]Α������|'����ŋ��ZG�Z���7o�ʕ+��w�����S�-������O�uzQswi���$IB0��n׺"""" ��?���B"���֖�����������?��:��.]¥K��|׮]×��%<��s�\)�vx���f3&''Ή����� �׋.@��k]�>6�������/��ἕ��_��W���~��h`q��^�^�W�2����d0p��ylnn"�J����o�6}��=�k4x���w�5�B!|��_����]?�=��#�x�"����X�c�K�Љ������j�"""�^'�"FGG�t:���EQ��k=fgg�|�$��|>��կ"��s�s��9��?�3>�� �Nw�����-�D-��vLNN2�Q_���x�f[���S	�M������>Qd����t�]DQ���,�Z�BDDDt":�gϞE4E$��k�c�=��s�5�B�=��y�D"$�I� �˅��<��Cx�[�����9|�A������?��ӿ������!t��Njss�<��e�1����d���HO6W!"""�[~�v�KKK]�+>66�}�Cm/�J��׾���A.�k{�O<Y��я~�}�{۾G���?�'�|����$���WM���A���A� ��nLLL0��@2�͸x�"l6۩��G?�Ѷ��c�}�Q<���G
��t�����mϚ;�N������j&��4�$I����~?Aк"""�S#�"Μ9�P(tj�a����w���c�D�>�(�����/��2>��"�Ͷ|�=�yϱ���1���2�����ls"""*^��Ν�$I��-�T+����˿����]?���>��O�|lbb333w��D����������$�֥u��lƅ`�Z;��=�P���;���˗O��O=��~�閏=���'~~"�1��PE�p�p�[ډ��h�I��3g�t�#�����������ޱ����������:�DZaw����\5'"""�A�.�F�Dϥ��066��󋋋x��WO�ܻ=������F0�����鎽�V��NC��trK;Qf����
��9dY�(�W�^=Ii�(���^zi���؉�:4Q
�Z�� """��5��_�5���o�կw8-?���/���#?�N���l��ku,�N���qȲ�u)DDDD}AQ<�����?EQ��k�Ng�����N��G"�h��v7	��:$�ٌ��ɖc>�����`sss���?�L&s�_�.����t�,U��Щ�1����e�����������n�R)<��cG��nU�V�u�, @�Ri��Ә�N�ML040A@ ��v"�k�F�z�F�F�Z���Z�BQ��u ��l
� A�Ǜc%IR�,����Ծ�$AEH�A ������!E�s���j���(�>��Oڙ���W�Zř3g�D�����Vv����l6[���Ŏ�Q71��@��t�v"���J�RA�ZE�TB�RA�VS?�ժ������u:t:���?߉�5�����R3�7k�]w�F�(���t�� A�͏�M��?�h�	��`0�͆������E���`bbb���v{�kj�����Щ��f���pK;�(��(��(�J�G�s�P^�T I�F��O�^���� �N��N�f��V�G�5� @���	����E�i���z]���j�?���fÅ�����z�+W��裣���UC:EQ�uf��1�P_s�\����&�hX�J%�E

���A��a�h4�d2A�e5��U<EQ�i�00{nvX,�FH���fh�����<������Yx<�}��jw��َ���9���r�_���Щo�\.�� �c*�J���j/
j(���z=�f3L&�v;�F������h4��
�H���$i�w����	�N���W��}�މ�O2�ć>�!�������^�x���}�������u:�I�022r*G��s�A<��!�ˡX,"���[���t0���x<�X,0��0��-Wf�w��u���5û�dRo�X�V�F P�5{��w"�M���_�*������^;;;Y��N�;�ڒ$�ܹs�>���ܑ�'�:�������Mi�^�cgg�l�l;;;����VEEQ��b�,˰Z��X,�X,�3څwI��2f���C�!�<O_�V�4�k7k����?������O���&Q�ַ�O>�dG^��a6��}�ƍy~"-1�S�0���y"��e5�7��j�T����t�j��a�d2�_�Q���M� �h4��)�7rv�T��j{{�R�6y"-//�O��O���~���w��]�������jG��HK��dYF ��{�.j�������A��l��f��nW9��PE�п�^�W���M�z]�ͳ�\i'�L&��{���'155����m�D"'zI������|�\��������0�S���|�x<Z�A4��,2������Z�f�6������gt�ժ��	���Ps���fS������zsϴ��J��O~�x�߼o� ����8���������k׮��;t�Y�("���HD��(
��,R����j��WǝN'��QOPE=��� �~����v;,��s��h�R��c�*�
WىN�իW��SOa{{��������y晎��Щ'��z����Q�4�=a<�N�3�wEQ7��}�~Q�����K��ժ��Z�0�L0�L ~���2J�;Q�|>�F���t�9� ^}�ՖgͿ���w�u��ĀN=�h4bttz�^�R��Vs�<�H �H �����    IDATN�m�՜U-�2�N'9��}��o@Y�V8u��؝N'E���x�����p�ܹs�}�vGn~E"|�S��@eD���z��b���h�1D�^�XD"�@<G2�l{޶��W�eȲ�-�44��:x}K���"F�Q�p8{��7W؉�x�f3.\����E�j5��!�y��3�N'�� �MQ�^G<W?ڭ�������Y�yt��gj��z���n����Q�l����(�(�(�J�OtDz��ϟ��۷�ȍ���\.�~?�9�!����h�D��9r��։�F�\F4E4U��7�H��N/hn�ovv�':�$I8w�������.��g1���� dYֺ���h4�L&����Q(Z^'�v��m�sȉNf�v���u��f88�N�l6��n��e�j�RI]]'��DQ������՝+D�:iFE�B!��v�K!�)�z�D�H�h��=Qa���r��v�y���5W�#�t:�zl��p@��z��z��v45�
n�'z���Q��D'D�	I�022�U>���V���b�F����m;�����	����ͭ�D��jH&�H&�{n�5���������۽'��;�B4l�~?�z=���;�|>��(2�S�c@������5z�J��ۈD"H�RmW�$I�����������h4���º 0��0��jX/
�Dx��^����҉��� ������c@��ǀN]e4166��_z4�j���(���l��\)��|�e������ ���w7jlv�w��(������4�l6Ν;�;w���A3���}�S'-�$��Ʉ��1nɥ��<S����X,vh(w���x<�D}LQ�}+�n��,�K�M�\.���^,�i��f�;w����~�˲�}�C�4�Щ+�V+FFF8hh(��x<���MD�Ѷo8���}>ϔ��+�$��m6 ���l0��������h����q�֭�}XdY�����GU��"t:u6��p�ᜆB.����&677Q.��^g0��z`4�X!i�^�#�#��`0��r�����v7����(
���T*WNt��z=.\����E�k����:�*�Áp8�uD��Z�"�`ss�����$��v�����tv�B"�E�J�H�HD����xԝ4�$�n��n��Z�"��#��q<4I�0==�h4�����x�{�˩?4T��Ը�n��~�� :�� �bss�x��-��~�.��;I���fg���MȲ�Nmh����eN�S�_,5���􈢈p8�����G竫����8�ʈN:�
���ϧuDW*��������χ��z�|>na'�ci4�u�����ǣN?�}^�^����ZM�ʉ:��h�3��{�1<��m�[]]ŗ��e<��-Ϯ�t�(A ˲֥u��(H&�X[[C4m;���Z�r��N�DDw�\.cccC]U�z������$��p��p�YUo�=���(�������?�<��C{c0�AŀN#�� ����8�j�����"�8EQ�J��J�Z��?���UuD����J���~+++��W��o}�[��@��:��E"����*b�؁+Q6��`n��gˉ�+v���\.���=gtw���Ed�Y�k���(
���	��������'�4�Щ#B��9��z��H$���ed�ٶ׉�Y�
��l5%"��ћd2	���׻�fa�z�VC6�E.���w�k�dn��x\�R�N:�� ��*Է��"��ְ���j�������`0����
��V(������-u��^�W��tp�\p:�����f���N}+ C:,t�k����VVV����
��v���zZ�ZE$A4m��]Eu�z�P@6�E�\ְb���P�("�jR�͛7�����kߍ�vR�a@��"FFF`�ٴ.���EA,Ý;w��d���t"��ru�:"��ؽ��f�!�;�f�X`�XP�T��fQ(����J   MB���Z�_��:� ��jպ�#���������
�B��DQ���A(ڳ�DDԯr�r��f3|>߾s���N���ԩ���H$�u)DÀN�"�"FGG^�/T*���buu����$���!�|9�b����Ulnn�c!%IR�}N=��!��r�4��� �40��Ț+�����"�ܹ�����`�A�=oT��U�V�����(�^/���y�(��p�n��A�����~�����-�K!:1t:��s�s�e�`���q�M���p8��@'"6�ђ�hT=ڳ�� jC�|>�L&àN=�����hp%��:����r9,--akk��`n4
�̉�~FQ��q$	�\.�B!��=�X�VX�V
d2��i���CQͺ�u:��z�q����|>G������J��r�a2��\���^,��dP�T4����@ �F��9�Է��@�p��z�������l6ctt�3̉���A�U�L���ٌb��t:�u�9�`�� �Hh]
ѱ1�S[�pv�]�2�T�\�����/3�9�]zcPo�������4ϨS��PH�:&�'贏 �p8Z�B (�J�}������z=B��� Ϙu��ު������KA@8F��@:�ֺ�#c@�}� �N��e�\.cii	kkkh4m���t���DD���L.�L���"���<��r9d2�Q'�	����1 `H����N{�AȲ�u4�*�
�ܹ������I��P(�P(�9�DD]�h4�F�L&�������l�Z��f����9�+Q7���rg�tR�|>�s�T�^���*�ܹs�RA���0::��y��Z����-�b1��}=?A����fS��AG��N� �����Ύ֥��  .��G�2hH5g���ϣX,x������,K��#"�vj��������r��<.�"�N'l62�r��F�Ұ7o����
&&&�.��-�$8�N�ˠ!�H$����ڵk�s�͆��Y���0���fϐ����!\�$��n�B!��f*$z}A����C�%�!g��
��.��P.��իW��/"�Ͷ��h4��ٳ���{9Y������y,,,`ii	�Je��z�>�~�_7x�n��j��'>���ԳЇ��jE8ֺ2�r7n��3�<�X,��:I�0>>���>����I�R)ܸq-�}�L&�B!��nNߠ�+����?�3
�K!ڇ����l���(R�4����駟�����͂|>��~���=M����(��H$��^{�x��56��p���恵��<������ݩ�0�!�����Q�s�d2�g�}sss� ��l��{p��Yn}$"�j������C>����(��e�P&�I�
iX��i|��к�=�І�^����gFSW
\�vW�\9�s��`��������.VHDD�R(0??����7ku:�~?|>t:����������h]��}�H����1�Lҩ���XXX��˗�*�"��0��~��~no$"�d7n�@4my��l6#
��t��u������/h] �A� `dd�A�Rh�E�Qܼy�R���&''92��h��u���#�ctttߔA���T�ͼ��]�rO<����7i]
9�! ��0���R�����Cg��t:������w�2""�U�R	���p��ݷ�]�$x�^�E�R)6��S��o}����nb@~���z��4����֭[��P��|�����B""�#�L"�� 
���k6�a2��������'���w���l�{��&�Kpn�.�K�2h@�R)ܼy�l���,Μ9�EDD�Vs�{:�����f�Ǜ���f3R���F�Ҡ�����۷=�Gt������Ӻ@�j������8�:Q166�`0�F?DDt$�\sss����B����r9��i4�*�A%�"Ξ=���y���c@P��P���:�8Mদ�8Ӗ���MQD"�R)LLL�܁e����t6��NE�Ν��ܜ֥Аa@@F�###��Q�r7o�<�	\s�_ �� �H�R��[���z122I��<���\2�d�/�(�^���iܺuK�Rh�0��N����}?��N"���^C�R9�:Y�155�q~DD�Q�x�Lccc�ey������t�ͽ��L&&''����u)4$�Hsֹ^�׺�R	7o�D4=�:�N#"��V�Vq���\.����"�"�n7�f3Wө��v;�� ����.�� � 	�B�:�ݭ��5��������̙3�FDD]�J���f1>>��t��χR��t:���q�l6�K:�\.���U�ˠ#�;�����p8�.�@�\ƍ7���N�$LNNrR u]�VSW������k��[,$	��SG����\.��BZ�sd����}�} 8x<�ˠ�Dp��T���s:�8{�,Ϛ�����p:��7�L\M������:U�}�9N��$*�
nܸq�YsI�011���DD�3j�n߾ݶ�{s5�d2!�Lrn:��(�H$��EQ�rh 1��1�^�qjtb�X7n�@�\>�:�ݎ�g�r�9��x<����:l�X`2��H$P,5��E�����.^��u)4�xۧO���qjt"�Z���
�^�z`8E���e8'"��V.�������(���qQ����v���I'R,9z�NW��T8��hԺ�S�L/��2
�י�fLOO�b�t�2""���D"�f����lys�f����� #j'�J�b���uo�!���W��������^84��|>\�t�ᜈ��R�P���\��*:�~��es9�����@6�պ �}F�e��n�ˠ>T.�q������ G�$LOO��ٳ��GDD}��h`}}w��i�y[8�N��~��v���C'��}��Ʉ@ �uԇ"�._��d2y�u���w���@I�Ӹy�f�Qk�qlf��˕� P7o�� ��>���0::ʎ�t,�zsss�v�ځwvA���(fff8ۜ��R�R��[�������f9����[tl�z�o�ֺ l�A@8�N��]tt�|׮]k�Z�d00==��ޥʈ����(
������099	�^����
�^�x<�Z��A�ԯr����
��.��W��@ `�.:�H$��{��p�p8p��2��P�f��y�f��^��P���ض������u���{���,�Z�A}��h�[����������V�V;p˻ �z�p����N�r��6���ƀ��L&����eP�(�Jx����r�uz�333�""z[[[X\\l�l6� �ґ)�r���v�{���qD�Q<��3�d2^�p8p��%�|%""�eggsss���-7���NGV��p���ˠ>Āރ���JQ���㥗^:t+���W�V����h4��qQ��zy���,��bssS�2��0� ���;�t�j���ׯ#�Hx�(�8w��nw�*#""�O��`}}�B�����kY�F��x�z]�*��D"��v6�#�
z����Rt�l6�g�}��pn2�p���k������$P.�[>n4�+�����ۼ�CGƀ�C�#=������{�b���N'��^�� ""��B���mG�I��@  ����ʨ�(�����ˠ>���#DQ���H˭TD�Ͽ�_�~�Ю��p/^d""�h�b�D"-�����P�R	kkkZ�A}���{D ��hԺ�Q<oNDD�����Ŷ��m6t:��8GkQ[�xN��C�R��q��8�����z��h4�9�)i�Ko75�d2!B��w�2�'w��A�VӺ�a�k��$j%��^8����f�ys""�SV(077�B���q�N�@  ����ʨ_(����9�ˠƀ�!�;�������ի��e�x<����{""�.h�KO&�-E>��ۘ��j����U�ˠ�d��`0�s紏�(�y�&���(ʁ׎��bzz�7y������h`yym��e��Ψ�D"�T*�uԃ�$N#�,��*�S�Vq�ڵ�w�DQ����^o�*#""�7�D"(�˘��d�8:���e��vNݡ=���ш@ �u�c
����Cù�`���,�9QH�Ӹu�V�#ilG���׺�1�]&B�ge��T
�>�,�����Y,�{ｰ�l]��������177�R����f�8m�7�T*<�N{0�w����dҺ�!�H?��Om�p8p�=��`0t�2""":�J����yd�ٖ�����ω+�O"�@.�Ӻ��]d�Z�r��.�z���
�_��z�~�u>�333�$�K��q��u,..�=�&�^/��>����S@ лF��!
i]�����#uj�8{�,�E�EQ���������Ȳ�E�CQ,..j]� �.h�;g�F^�r��u,--x� 8s�&''�Su�������>n�����x�T�|�hT�2Hc�]�r�`�Z�.�z@�Zŋ/������E�ϟg�""�>�Fq�Ν�[��f3�@�m4�666P�T�.�4����d2���i]��R����T���t:fgg�����h ��i,..�mk0�ӒT�6��O�(���ܺD���x����֜q�1jDDD�#��aaa�j���z��!�T�Z���Z�Aa@?E~��#�;;;x���Fm2������""�T*�����v��$I�|�H �T*�vd6�Sb�� ˲�e�ƒ�$�\�r�Y"�ł{�&��K�Q���e��ϣX,�|�9+�����hp1����Pn�hW�^m{��f�avv�w̉���@�Z���B�co�(���qG��h�Ν;Z�A]ƀ~
x��677q��u����s8���������u�vvvZ>.�^/{�����i�0�w�����к����
^y�C�$y<���p�
�j4�}�6��t�k�n7�v{��^���̭�C��v���8�z�---aaa���|>�����h@(�EQ��FcϿ���5�k4�.�浍F�F�$A(��NA IDQ�(��$I������(XZZ���d��.�� �]m��p��-\�pA�2��;(B�$�� �ܾ}����^���q����&�A� ���`0�����������^��Z��Z��V��V���o�{���Q��4����5_�Z����Z�k���{~/��C�[�!]Q����43��B��x<�׫u)t��;D�e�b�n�:R�@ �3g�t�""jE�$�F��z�F5���z��e��e�J�=��T*�T*�
�ij�����#]�(
�ժZc�ZE�X��Ύ��i4A�=�=&�	&���n�4����.�ɲA��d�\����u8��#�l��Ā�z�~�_�2H#XZZ:��`0�����/�hȉ���M�Ѹ磹�].�Q(P,�J��^.�5������v�����������34�L0���D]���
 mC��� �[���(
nݺ���Y�K�SĀ~B�  
�Mː�������ׅ�a����~ADCD58��f�FX,�=!�\.#��#�N�X,�T*�X,e����7��RE��bQ�s���{�� ꟱�d��b��b��l�y�Z]]E��h���p8 ;{�r�������!Z)
�Xu�	ɲ�9�Cjnn+++�^�pNtrͭ黃��b�ss�P( �ɠP(��ZMê�� �Jy�+�zp/�J{�<�J�Ҿ_o6�a�Z�|��5��[__G��@0l�x��;C�p���|�2�(������|Z�Ax�װ��v�u###�BED�十�d2�y�\.#�N#��!��!����ijo�����硽�g������X,����l6��+�Dǳ��	A�NbH^�(brr�H͉��0��@0�
����;R8���DG I�V+�v;,˾�WEQ����f����\.�j��a��kwhoޠ�������n�4C{4����6��v���O���.J��    IDAT�A�nwgH^f�n��dR�R����,˰Z�Z�A]���p�m��`��ډڐ$	��C]!߽��(�Ƴ�,r��:/�z�$Ip8p8 ^��W,�������������Ύ�2�\e�e���c舆���:Ah�k�n�CQ6�B�P�t�;���Nǭ�C�֭[G��ح�hQa��`���p8`6��]S.���d���%��#��������(
Eٳ���uN�S]�]jD�[[[� m��7o�1�Q111q����?��B ඼!s���#�9����sN�b��n��n��Z�j�L�t�L��n� �9�P(�F������Q��5�|>����&DQ��nW;�Ұ[]]� jO�7r8��/�cC��>8Џ�yn������p�|>�sZ�(�j���t��rA��ﻦ9s���y�/�(B�e�c|�\F6�E:�F6�U�j6uG���*�z=dY���,�\]�����Aڎ�j��bX.cccx���su@0��$Im�t�`Z^^������y�^LMM�C1�^�vdEQ����d2�T*��nԒ�h��h���Uϩ7wV�>�P�V�������v7��U3��\���˲���� �"��Ǐ�'�z�1��~6�"G
�.�gϞe8��`0 �2�N'l6۾���g3��,9�$Ip�\p�\��T*��O��@2�D2�T�л\.���}#����(X^^�(�p:�-�i���r]���b���K��K0w��`����b�<���M��۸q�ơ�9LOO3��@3��Je�s��z�t�D�L��d�#v�]m֛+��l�����lp���x<0���N��(XZZ���t۩Bn�[yH���^�_�"� �9�#�w��H"��+��r�9�ł.� $�NY��v�a���=��Õr�va=�L�k0�ﶺ�
��
�����m�4p�1==ݶ����QG��+���W���}�cZ�B'��~^��?؇D:��K/�t�
��l������@�$I��a��� �#�L2��&v�����H���ξ��ͮ�+++p:��z�p�ݼ�J�^����۸p�B˭�ͮ�X�rY�
��~����~7FFF�.���!C�N�4X��,�^�zh�0�x�"o���hn	n\*�
��8��(��QOEQ=�^�בJ��H$���m��H��j��@ ��k4��*p����!]E�|>D"6��w����Z�Aw���`�狇@�X�O��Cp�t:����\#�=�^�������^�#�H ��0�I���z��zQ*�ԝo�������`���E ��u�k�J����p�B��}�(���#��;B�'�੧��o��oj]
��8�ζgzhp��e\�r�ЕAI�033��ܥʈ:K8�N�|��[���<��(���S�2�L�����z�鍽E*�
677�����������ԗJ��z&��n���H$���C��'�����vN��C�mp��p�����Ozh�Ap�����R�zYs�������h4�N��F��d4���t4gE�\.��e�b1$�}+��� �� ��pU��Z>�������Z�h��t��|�F���1�j��q��_��֥�11������ l�5\�v�H�w���xV�������k��[*�����x<��xF������H�ӈ�b-gD�^Uw�\<�N}'��`mm���-7�x<���N���v��u�?���f3��^{�x����������P��I������v[[&����6��t��#Ҟ(�jS�b��h4�d2�o5QQ����dB0���gx��x���`���˅d2��ʨ۾��/�K_���e�1�.]⭳78s������Eܾ}����~?����P����zx�^�������:b�"�J����j��d2�h4�J���:I����
��>�����<O�ǛG;h�E"D�Q���i����/�Ę�����������~�p�r�p�̙.TDt��V+� dYn�x�ZE$a�^���z�|>$�ɶ7���:����D�v��ٛ�z���*C�ƠN��z��q��m|��w��t�z�Z�A�(���^;�:�Պ��iv�e��<[*��;�lDt4�(������ �� ��.�� �H �H�n�#��riP1��E��۷q�������n7j�wW0Q166���%�K�#`@�����l� �����k�m�b4q��E~-P�iv�m���r9lll�|9�	� Y�!�2r����������l6���yX�V�����r��.��F��;w�����-'y �����F��;|�X�VX�V��y�K�C��ϘL&LLL���*�Jx����;,I�瞶w��� <ρc���,677̉NI�X���R�ԁיL&�������=��ł��Ϸ]�h��T��U�T0??�u=��Π3�����dێ����?{w��v���Y{��*��z���X���B1�pl���X�L1��#�(O����`>�U�<�&����`��H�䥸_v��F7�{c-�Z3�Ь��}QyШ�s����{;��:d-������i�Z���~W��}�9e�0E;cԐ�R����J����urr"������X���ddrrRFGG	�a�b�(7n��x�^����&ǯ������)F�� �0�bQ&&&�����ߖ���k׮u<�S;0�|�r�r���}YYY�T��Y���	�h�1���err�����c��<O�߿�"�KL
�{~�뺜qc�?�
����	�a���a��������2s b�\N�]�&����Kj��,..����LOO���0uDjssS��l�������E�_�)�uerrRVVV��
:�� }ddD�ɞ��!�666daaA9n``@�^������ejj�c󷣣#YYYa�9`�\.'7nܐ��#Y]]�J�r�Z�&sss���&SSS244�L��s�Z�ѐ���g�0�J%��ڒZ��Tp��.qO��r��uV�c���@���(��r9y��7Y�Ad���err�cc�YYY���ݐg�<�}!T�M�P�+W����@H3�+�Lʝ;w:�8�}_�={FS'''277�4�aR�{O�SSSR(��.X�Z�o���J2��|�4D$���LNNv�^4YYY���-����ۓ������J��\�r��C�l6+w�ܑD"q��V�%����l6C�°��Ė��0)@�ٴa__�y�Z-����Ǒ�7o�#t�TJ&&&ddd������Ɔ���q�`���A)�����}��ߗr�,###2==ݱ���jU;vvO$222Bg�����$@7P��cccQO]�������i)�J!�x�ݐrbb�c'�gϞ��ʊ4F,�xE����ؘ��Ɔlmm��y����lmm��Ύ\�|Y._�L�w��\.���z�������N�3C�%�I�gϞE=��'�R��q�쵴�$����q���r���f<��̥R�S�����<3 aH&�255%###��0x�'+++���3�z�j�.��E[__�{�i����^�wl�{������0=�<�n��R�kooO=z����;�q-����۷��ի���z]����޽{�@�f�r��-�q�F`��^���Ǐ����t�Fh�<y"�j���R����j�s�\�>44D�V����Բ�%�I�}�6e��D"!SSS��k������<Y]]���~[���#�!�(�J%y�7dzz:�tpp w�ޕ���t��<ϓ�����Ǒ����`�R�Ա���H%�Hp�h̴�©��:�#�n�b�]722"��:��888�{����ʊrQ	@|������288�q\�����~�}��Z�&KKK�'	��qG�����~�������1s��}�p��U!��˝;w�ʕ+�f��<~�X<x '''���������͛7;�7YXX��]���/��������E%ة���D�!z&ZM��t펙��eY[[S��)��u]����;w�H__ߩc�ٯ��ݐg��bQ�|����D���}qq�*t���z`�P(p\q�8�#���QO�C����81R�TdvvV9.�N�]300 o��LLL���rtt$��ݓ'O�p�9 %�u������k�u\�y^����!o������g�^�����ppp�}�1��f���?�i����s��|1�l6�?��2�q]W�ܹCS@\�d2)ׯ_�X��>*�wޑ���f�f�\N�ܹ�l"W�����2??O9\�f�)�����rGFGG�>3tt�^O|�:5k���޽�����ի��<�7������P�ݻ'����)
���y���*�����6t���a�~�d2I�I�R2<<�4zZ����~��rQOdqqQ����𰌏��0#�T*%333r���S�2<ϓ��ey�wh�¤�i�}��\�z50S�h4�ѣG���#i4!�q���!������yʢcf||����}����H�S���ߗǏ+�e�Y���	aF�CCC2==������C����j��� 􊑑������]���R�T�ڵkd�pa���$��w<i`ppP����j��g�nH$266&���QO�'�:�>00 �L&�i�4����X뺮ܾ}�c �E2�����v�ک����� �-�N˭[����?�G��7��j���B�֭��a���I����[�8���w~��5���!�qW,���_�x<c�C��Q p�FFF���_W�Y��ݕ���tzǅ8>>���Վד�$U1�>F�m�^,;���.KKK����744DC@�2�uejjJnܸq��1��ۡ��� ���f�Ν;255��������YXX��t��gϞ.��r9������U����벂�JE=z��N��w�W���'���zǅ���Fth`�qd||\n߾������3�{�.G?�---n�(�J$�b�u]�t�R���9��K�ҩ�/إ�j�ݻw�+����͛79��dll,�!wggG�ݻ'�J%�@���>y�7�ɉ���w���Ȉsk��މ�82<<L��Y�t�u9�1&>|�MNN���@3B%�I�y�LMM�zj�Z�������� c��+׮]�����F��m:>�z��'��ަR��=\`�qdjj*�i���胃�dRc`ssSVVV��
��LNN�0#�Q�����xڍ��B �$�����o(ȕ�e�{�n���@���U9>>�x���_r�\�3B��E��*@'{�jU�y��D"!�nݢ�g�8�LNNʭ[�:n���ޖ���s| ��i�}���qj�ѐ��YY^^��g���,..nE���h?7!�
������r��]i4ʱ333�s�3K�Rr��-?�z�Ւ��9�����1 k��+���233؅��}Y]]��j�{�U����G7�G?Y���&@w]W��^������*Ǎ�����3����^{M
�©�ONN�wޑ����g �188(�����Ը]�N#L����v�V�l6��k1�8�\�|9�i����g���C���W�K��r�ڵ�O�266&7o��XҾ��%����ls ���f��^�����q�z]�߿/kkk!�q�����
NX������C��6�H�=���yr��]i�Zʱ333��@["��7nt�����,//���%� b�u]�z��\�r%�w������Sy������l6eyy�����k�Y�p�"@/�J��XnaaA�����8��2��ܹsG���כͦ<|��l��1::*�o�Vf3www��ݻTA���~�6�t:��~{�E�.�>@w���;88�'O�(�e2�z�j3Bȝ;w$�͞z�}���� �I�P��^{My[�/G�\if���������$�N�8#\4�qdbb"�iĚ���� �8�<O�ݻ�,�sGnܸ�{-���r��͎[!�������R��B� ��}�j_:�F8�V�%O�>�x�]���v+�J��]du�N��~�?��;11!!�6s]W�_�xV���
��@�i_z�m�}�sss�vB���@���:^O�R��[����eu�^*�hf���=YZZR���r255`�T*%�o���0��jɣG�duu5�����Ǖ祋<?N����������*����d2!�mpp������Wɞ���<�����8�q����\.'w�ܑ|>��z�.<�����g v(�J��k�)�W*�w��43����Rw���r��ȥK���F,Y��E�S���ܜ*Ǎ��K3������*�޽{rtt�� �.�\N�y\�V�w�y�EO�T*�����z2�d���Yd�kt���:88���E�L&#W�\���`���1�y�f�恻���c�����4moz��YH3�������$��溮���E=�ر2@�{��/�󎲴]D(mG�˗/�&��ܔǏ�� ��u]�qㆲ|��}YXX�ZtGoj6��Rw�I0���Y�fe�C��^O�<�:wzll��8��8r����Ǖ��MNN������{ccC�����{�����w��J�(u����f̺ =��K6��z8���#YXXP�K�Ӕ��T�dRn޼ٱS���277G�v � cccZm[[[���i�Z!�6y���4�͎�)u����h�S��tVh����ܻwO��}��5�����R)�u�VǦ��VK>|(;;;!� �T*��h;88����K�^if�E�ٔ�����9��nTA\,���t:��,
3����7��J%~��>�LFnݺձ�D;8�9  pv���r��m���l�utt$�����T<�=vwwehh�c ��d�P(p/�����������Z��/����Cy�(X�A�D;�j5y���r��r���f��r��c����ܻw�: tY>��=n��jr��}�J��,//6o-�J�J�issS���Cy�_��_��|�#��V�	�9+�^�=�:�jjjJ2�L3�-
��ܾ}�㾴�����T�Րg �)��ʝ;w���z�.��ߗJ���`�Z�&������K�`K9�#���������\�z5���5����s�����ښr\>�����f[���=�GGG�����j!� z[:��;w�(�6�My������flll޻��#,���Z/�\.'���#���_亮�J����3�<O�߿�5�ڵk,��]����]�+��<x�@�2 p�ɤܺuK
�B�8��dvvV���B�L���,//��tZ��'�'���O��O�o��o��za�"@���H�-..��ёr�����R��`S�Tdvv��|  b�D"�t�6���ѣG�����`�����E������u��>�)�q�Fh�+�^����V�Zg�'�I���aF���А\�~�� ,ẮܼyS���/�?����f�-//�ϋ�"��Z��}������^/�N�g?��X%s��_���߱A�u��}� �ʕ+����4e���<|��� ��UO��e~~� "�G���z���P�n������~h���?���я~4���6�t���y��lmm)�������h3��FFF;q���ˣG��f D�u]�qㆲw;H�yN@�mmm���I��\��q����}-���ԧ>%��㡾f��g2���QOg��g���ի4��˕+W:^/�����c�s 0��233��/,,�C|ߗ����1��d��}�s��^__�|�3�	�5��� }hh(�)������Í����2<<�9/��d��"g�)wG�R�����דɤ��̳��%������>�!��_��P_����_F��j5��p��fL�J�R��R��9 ��t��q��󡝛s�����Ţ$�g�W�8��ٟ�Y���������B݋dl�^,cՍ�<z�H�ͦr��Ԕ���fSvk?<<�[; X�,�����8����j5y��Y���(�2`������011!���'B}͋flLs8���eY[[S��d2r�ҥfS��9?<<�[; �@�q\___�v�T����ؐz���z�P���    IDAT �c���/��/Cݏ��233��^#t�V�σ��]�z�ʈ��������9�I$r��Me�i�����AH3�i<ϓ����1$����k"������^��y����J�R�S����J�\V�+�4��a�|^nܸ�q��Z��Ç��I  �L&��͛���y2;;+���!�����l6�	O�����կ~5������9k��g2e)��j�dnnN9�q���l6+7o���7���,m �+�N��۷���VK<x��U�Cu���� ǮY����#y��|�3Vn�0.@'{n���%�V��q###,���t:-7oޔd2y��V�%���Z�# ��2��ܺu������hȃ�V��43����H���:^�'�loo���z�;==-��k���*�t�q8�"�z]�<y�纮LOO�0#�&�Lʭ[�:�^�����  ���dffFُ�^����,۞z���Z�偁zY�����#y�O~�2::�k�W��+J$2<<�=>��pơE���n��.]�����ݽ7��t3??/�J%�Y ����/ׯ_����� ���X=z$����X���j���%ccc�^w]W��b`�fy����п�}}}�[��[���~6��}]Ч���o��o������<~���3�E999Q�y�A�|�r3�i�]���aii�so�G�J%�����O��;88���9�u���{����wL�
�T*TYX��jɗ��%���?�k�ʯ����_��<|�0��>c�#����-2;;+��)�MMM)��!~����I������F�3 �fttT.]�����+���ݟ��j��ǡw�e>���G�������D���aL���/9�)@S�\���M�L&ӱ4	�511��gggG���C� �T���Z�!777#i2�hmmm�������,Q5�����y��?�k��z�^�o|�QO�fgg��]�r�=c=fhhH&&&:^�T*2??�  ��r�
帧O����N3�)<�Std��U�8�O��Vl�1"z��7�IgKlmmi5����244`���>�z�j���jU?~� �{t������/���rxx��`������X3���r�g�W�n�7�|S>��E��gaD���/})�)@�n�szzڊ*\�t:-7n�����Z-y���4��g �A2���7o*O��<O=zX���Qeы�bH3��j7���o��o�+� }iiI��梞4lnnJ�\V�+
288`�v�#��nnnN���C� �6�lVfff���z]>|Y����|�H��d�-U�8��[j>�D��:"�ig���R�\����������L�MqqqQ���C� �V2==�w||,sssl��!kkk��ًn���-������O~���H�f�)��ַ��4���k������fLNN�ߛ����  �3::xH�����0#���� �gU*��|>�p^���_��_E��������둽�J��w��]�T*QN<�;��s􆡡��c�*��,--�8# @\LOOK�r���*��{�NGwz ��?�a��������&#п���E��д����xppP�f
�������F��C ��9�#ׯ_�T*�;??O��qpp��K&�����p^�z]~��D���B��,zdz�\���~;����V������yoH&�233��{��dvv�� �W�J��ƍ�7m����f3��!J���d�-��}.�����>fdr1� ��_���Z��^�VWW�V�)����3�t������=b  ���듫W�*�U�Uy��1�[=���,zL<y�$҄N�P��~����~'��0��y������/_��l`���������M���
qF ���jW.�i�#t��0����/|!�9|�c3nA'� �ɓ'4����ښT�U�R�$�B!�!J�R)�)����k @WLOOk=k������n3B����O"�n��|�+��~�X�_��_�t/�$@�9��|��ΞONNvy6�Z&�	,1l6�� ��q����d2������=vSut/��E�����looG:���������dC�[��|���eqF���ZQ�l���㺮\�~]�D�1< �-�JɵkהAW�ٔ��Y�</��!
�JE�E�?����/��~�T�~����t/=@��~ �r9���%{>55��� j��Ӂ7���5���qF �^U,�ҥK�q���l����ًn��~��QOA����&"F�����|����+�m���������w�^�Th� ��ĄV�������0#D��� ��3�J�E�@�Z�w�y'�i���Y�P����H�����y�qd��-���m�l6enn�}� �P9�#׮]c?:D�,z\����M�S��E$�$B����Q�F�/�3z��V�<��K�XaF�B��s�������ٕ �ޕN��ڵk�q�VK?~�~����<u(�NK.�qF8���Y�>�E�ע�D�:��̷���5����655X���ɾs @���b��m���lǊ�gϞ^�����ͦ|�{ߋz""�QD"m�Z�^�T�޽{a�Ρ\.k]�LF���B��P,ett�����y��i�3 �t���Z����u�����N`�n6��L&��e(|��z
""�E9�����zKZ�VX/�s���>11���1�J��;�<O���( �u]���	ܒ%������yi6�!�a�}_���ǐE7����)Ϙ�1�-@���l'''�� ��gJꔓ�NW�\	l������n�  �-��jm���벰������d`.��j,��Z-��7��4DD>,"?Ջ������Ç�x)�ӓ'O�3���+W�a�������rY677C�  z��ƴ�����*3��S��
<V�q�������~;�%���7�iBW>tP��emmM9�u]aF[:��˗/w��j��:  ���k[\\�赘����9
��&�---��-��Ed"�-@���>}��E�t:���j�D����E�T -�N˕+W��Z����͑<��F���,��|ߗ�|�+QOC��y��!��z����I��`�VK�����NLD���.���������d{{;� p>���Z'�T*Y__aF���R�P�ٱ���/G=��� "���������-V(�����-�Zǘ�.�\.p��hhw� ���ӒJ���VVVh|C���rxx��z"��|>�pV������hHD>��v=@�������+�͞_�t��3A�Ǒ�W��"/--��	 ��d2�U��y�,,,�H�!�\��Ae�"Ϗ\�qAW_�qY\\��K��������r\6��R������佽��n�  ��T*���r���lll�0#�i?�B4�NK&�	qF8��}�kQO��<?v-4]�]�eU�`KKKZ����٫3�l6�*��j�� �ڕ+W�Jݗ���Z��0#���}e���f�mb�O��b]Ѓ�B#Z�jU�P�uell,�!LW�\	<f��ӧtm X-�L��Ԕr\��񲽽-��u����U������[QO��߉�dX/ֵ =�HpΠ������FGG�񊙱�1)
�(;� `���!)��q����l*�\zB�����.�)�%E�	�źAS6b.��duuUk���x�g�0������d  q��k[ZZ�z,ft�ű��\���&m��������Z�Ί��666�V�)��E������������U��  �P-N��Z-y��i3BXTG���˳��Z�����?�zm�"�o�x���|�ͦ{���x)�J�e~�jU���C�  ��\.����-���!�aQ5�#�h�/|�QO�E��E��
���R�h�xR����$����F9O�<1�� ��8�\�zU��yqqQ�O찷�'�f���L&���ј���z
/�e	�Y\W�h���keeEk���({rb���˒N�;^��ޖ���g @����dddD9�Z�j���|ߗ����1d��U��enn.�i�%E�7��"�;�#}}}����Z-�f�V��l6+�����Z-�m  �lrrR�ɤr���:g�ǈ�̽���Ĕ�>���G=�����fq���y�����.�FC9�X,J6�aF���t�Mgyy��� ���H$drR]��y�<y�$�!�j�fq�w�^�SxѴ�|��/p�4%"��-o'{����[NNNN8� �S�����=��r�9ڰ���uttdZ��Ot�/�� ��v3J�\V�K��244�m��*����4� ��q�ʕ+Z%�KKK4��	����K_�R�Sxѿ�+���/4@O�R����s=i��ǝ�� zR>��JHT�U���aF�6������n�SxQBD>֭��Bt>�f:Ks��fb�G:�ܪ�y��  =mrrR�o���
�Zb�fq�Z[[3���7�����gϞ����.&���o0���R��B�  fI�R211�Ǣv|T�U9>>�x�u]��r!��|ߗ���QO�E�E�g��_X���\kkkZ�t�������T*u��l6�+*  ����1�����rtt�m;;;���e��|�+QO�e])s�� ����T�V�?D"�X���C��mjj*����Z��f ��t��<��---�0#t���^`��l6+�DW���9=z�(�)��"r��.,����L���Z]�����1�������ߓ����
qF  �Mu�l;88�صh6��'9�C�P�jմ��a����^X���L4������˗�<}��c�  x������h<���ט�_�b�Sxم��_H�ι�f:88�J���N�e`` ���T��*�����8#  �P(������ȳg�B���\.6P��hs�(ND���E�����d���U�q###)a�D"!���c�; @g�/_�zZ]]5�'��Ι��7f���2��RFD~�"�B���<O666��R�n���1I&������} � �\N������3̥
���|H3�Y��/?�я���������^9@w������-�z]9������r�dR�=׭�  ��MNNj�J���X"�K�Z�x=�H��l����z
/�%y�0�B�r���jf�]��h5�]�t)�;���#���!�  ;��i�g�V��݈�Ru�'�n���٨�𲔈|���	�a�V����� �n�tZ�Eaee%��  `���	������4�f�n�	���d�����ꇈ\X�;z�6O���L&�-�.]
�q<{���0  ��J����x�'kkk!��R�V���k�o}�[QO�e�("��kz� �u]>��-�"{n7U����= ���ǵ�蛛�Z=`.�����[oE=���rA��_)@�k�V�%;;;�q�����P3B����[[[<4  pgɢ���n� =���o�@QO�4��"��W��q��y677�����t3B7�4��y  秛E���`/����z�Q���H6�qF�qrr�\\��/��+g@ɠǌnP622�噠���Ǖ�s�� p~�TJ�y��<�-�
�HJ��q��W��4^��_~տ��z2����a�����*�Q�n�t:�|`�i  �Nu�iYt���l6K�������G=�Ӽ�>�s�XI2��֖x�����/�d2�������;;;d� � �TJ��.{���h4�e�4�6���r�S8Ϳ�W*3?w�Ny�y8�<���s  B��V֦�f����N�n�f�)���QO�ey�Ы��������<����;88��٠[���K������  g��d�T*)�5�M�d	̣��,� \���7���i^�����D"Ap�lmmi��
�;K���<�&5  \���	�q���Z�a�Z�&'''����Lo��v�S8�/�H���t��ͣ�bKs8{�8::����g @o��r200�W�׵+a�r�x��<+++QO�4#"�3���	�c��<����Ky�������� ��t��8���E��}�ժT*���q������t���eooO�h�|>�{g�����c�ժ�  p~���Z�Q'''�@f:>>�Z����3m���z+�)�&� �u]�_F�{!�s{���onn���!� �ޤ�fk#�n/U�;�.�|�{ߋz
���"r�<��t>����N�n�|>/�B���V����  ���А�R)�r�̩*�RU?���<���QO�4�<?�����4K�R	,�iK�R���p�T���� ��q]WFFF��nllty6膣�#i6��'	�E����H+�����ɠ[N�Sh�T�����ɤ��Aw�  xu�����G�����@f�}_�t�x�<���HD�|���t�q�@F���T*uy&膱�����r�,�j5� ��R��ֶA��!�,�ck�����|'�)�f@D>x����ʧ�f�da�h4���:�#�b1��"9�#��ÁchB @�FGGeggG9nccC&&&x~���Q\:��u��f������?��]}�����t��	�-"_?�p� ��"�looku����d�Lo5P*��8�j5�  \���>����Fp�z]���i�k�f�)���{o9�#�l�F���k�����Űs.�����g��T���jf9��s�GՄ��9  ��:�����8n�>�����~V���k;S�������X&�������}�� @����$�H(�����aT��I\��r`deiRD~�,��v�Αf)��R�ו���4G�YH�=��ۣ3,  r]W�����XT���qk�؏�.:>:�z
�����Y%2�Nc��6�9c���  ��n���֖V� �Eu��Yj5cO6�����)o7����8��ۧT*���j5e�  �\.'}}}�q�z]���B�.�]<�3����"2�;���Z����j"��fR��Q& �9TG��mmmuy&�h��H&��=�8�#'�Ɩ�k�C'@���ޞ��P>�go�e��7z�m  �ohhH\W�H�����?�����8��dB�T*�V��K݁Zz*��m���?���>�Uxn�  �%�Hh��9�	<0���R��D=�N.6@g��Y��K�S �y(s�/��ۥ�06����hu��
�)�0G�^���C�8�q�n�����-	g�=   £������h=��� =�Nkmq@8<ϓV��4N����$�n���]�c:���;��<��p;;;�v� ��9��u&�Yt�4�M9>>C���|�V�;t�薷���,��*��qC �\��n��`�]*�r�S��_�R�T�L�At�?'@�K�XT�}NI  ���rZU��FC�ec�B�F2�,+�Oev�a��8�?�de����ZMYb#򼴣P(�0#\�����뺕   :�����n��7	M��r9������o����F��t^���)tJ6̡� �P(Ь�"�DBY�@� ������q���]��X��l��I��]:M�v������j%8C��:ts���i��{�]TNNNL�a  �H�RZU���i?���2w���p�����������j�������!@�'�� ��}����]؇n����w�yssC>���?�4g�9Հ� �u]�5�l6��0���#�L*Wڹ� `�R��U澿�o�y�8ő��T*�S���bv����ߊh6�1*"ׂ~�X	2����֪O>��d2p��b�M���ؤ�  ��J����O9��<��B�^�^�Z����8$6rZ���ʗ�G�$0�������Ǔ���i  اT*i��=>fPe�In��#k��|���l��g�.�[Bw�� ��DB�~q� �>��������n����u]������|�{ʎ�!8��|ߗr��5� �����j���  X(�NS�Cd��r�ҥ��Y�ٔ{w�l��_�H���� �}f8::�j"�L&�a������v  �[����'''���H*�1�B�FGGO��Ǐ�<��ɉ��.vГ�$�Ay{�8�#�b1p��  �Ku�o���3��'hPU7��4G������s�U�#p2���-o�)�������ͦr�  0W.��z��o��+{��    IDAT���(�Z�&�J����Ӆ��?��͠��ӆ9T�ꔻ `��d�aU�Ne������� �"2�j�Z��6t{�n�4� �~�:�}{��AM��qN=nMD�V�|�}H�����A!�n�r���G"��J2�aFxU�l6�����D^v  ^Q�P���t||,�Z�44���c����8N�Fq	7�lާ$"ӧ] �n8��Ǐ��k�R�f��l  @���K�{�(�ccc��y&kD�{�>�S�D"!�D�
�ΤR�nU�}�E  `����q���A�8{tJ��<�S���� ��9tt2�vp]W���>4  ��,z��0���I�u�B7�i1R�4(�l6�ټ�~��3�Z-�@[>���lp
�B`�F��,�  �H��Z�/��8n��g�T*��{ �wZ���33��T�:t3h5��d24���j��6  �2�xi6��~Ad�������o����f�>�E�}��St>Pf�T*Z�(o���M�v  �G��� �:Yt�app��.K2s�f��y����z�)q7�n�Ny��ɤr�:  �300�u6���'�XB��x���������ʴ�����8��� =^T��j���  �P"��z^�}�,�%Ƞۣ��}ttL�����#�������/@O&�Z+|�.����P�nU�vn�  ėn��n��"�n�B� �DB����Wg��0����PZ��r\"����%T7f�� �/�B}�v�V����Q�l�|>/�����LMMG=���e�=���J��)�� _��V�NNN؇n�j�x� ��lV~��M���䎼��A7�n�~��~0�jռZ�J��i6   l�DB�,V��6G��*s'@7��8��ˉ���� �PGGGZ���*o�F @�鞇�s�T�}	���8�������=e���� �A7�Nw;��"p#  �؇/d��qr����ȍ����<�S~��tJ��d2��t�F @���:::2�$?A�n�jU/������=z"�0����t||����H$XP���ʡ�hp�9  = �Ji=������ѩ���gv�t34F��ϼ�/��	�̠��Ly�T���  ��2w��J�pB�u��1wΠ�2��EU��
9  �C��]�yѢ���׊z
A:g�	�͠����s;� �6�x���|ߏz
A
"2�����|���k��d�_�  �\.���^��~4D�Z�^'�2���͢�A7����82��S�??99�f��l  @�\��N���|� ������M�O�Y�^�V�VK�G�q�d2!��B��= ���6��M� :�*�u%�H�4�ՂS"�n�82���!N���gt  �2��h�Z�jHb,3��>֘ �T�N�md��@�  ^�[��s�T��Ƞ��� }�����dRǉf:x���#��(�Y ���r9���z�.����7C��n�F������?�'@G���C�:��o   ċ���r,�O��8�-�3�?@ge��%��棼  t����������6""2��!����q  z����T%��Yf0<@wD�t��Z-e�LM�̧*q'@ �w�6�ӭ�Dtt����+z���_!�n݀-�H��p��*Q�� лt�j�*��wy6x�fS�k�Au$^�&E^�	���Z}k#{n>Uٚ�y��J   ��鴸���y��3"��
����P�����:���l�t��3��R��  @7�ζ8�������G�M�P�n��P蔷  �Fq,�O��5C����+"����DO�|� �|�  @���� ��3�#"?	��,hݠ� �|�  @�z|����&q�"/舞�/M�̧ZD�F  t��xn0_���e;�<������=��J��]Y��
  t�f�iz�����kY��^�ٔ��� �l�r�F���^ ��r]W���,��T%��h���j��ϫ�XIDd�����H$x��Z'{  �t��<?���l����c�M�E��tC��b�R�T�g�W��Ѳ  �؇��y�l��}_���a2�P�Ŵ���:  �E��>�\�sG<��2��:�����ͧz��� �6�g;�ͧ
Љ���j�p��)t3�lG0��ً�{  �O�I��#�n�OD"@7�xpG��  ���C�����KJ�A��x�yt�k  �TJ�Q��<�gé��%)jÏ;�#@7�xP��7�M�S  �������,����n�K��(q7]���v  pV�e�<G�� �M�+Q(q7M��q  �t0<G��.�v0����e%'z��k� @7���a�  x�n��s��T��:��}��{�.+9�k�Z����Xt��n��| ���>���M'@'��^�E
��
�R�O�sc  /#�:�dѣ�yFg�	�M��c�{e>�
��]# @����}��f�m�ӭ\�H�e'z�?�����=�  �(q�U� ���|H���U%�n>t  pVd�� �|�gt��&�n �xH&��}E�X ��t3��~DT�#@���z� � ��ǃ���qz  �w����<�~6f�,t��$%���Ƞ�M��pC  �9�I=<O�MU�@r4z�7�#@7�n��{e6t  p^�����Fw��HB��	Ƞǃj7T  Љ�s�f�G�~�Ƞ�@7pc1�l�+:  �D���f#�n>��M.s'�n�2�f��  ��n����؃n�78�·$z�A�U�np)  ���s�fSef����8��ߣ%�����^�M��k�  ��n�F���Ƞۡ�2����	tK��ͦz�� �Nt�2�wB�n�V�ح"�&�ͬ�^�M�sC  ��A�����<<tp�Z<�A  ���ǖ9��2TĚ����'�",���=�  �t��x�0��0�mj�A7�����ltq  �E�x���|1�{D���Ń���  tB����-t�A�t  p^��y<O �7v��&q& @��P @'<��%�v0���:pQȠ ��"��?v�ɠ#t  ��F��?v0�m"�n�x��  �m��������Xi��A  �Ew <���W�:�  @'$l��x�~�j� p�n�  �t�#\��w�U~���� �z�� �NH���������	�  zM����ƾOU����Wf��  �E����t�C�  ΋��xPmi�}6����52��Ľ7� �NȠ�qc��d�M�m<�A  �E��@������d�M@=<���  t�z�h�y�l$d,a��T�nt��n��D"��   ېA��Y�����ɠ@7p�]YE4T�+�  ��V��5� �l4���o�s��p��?܈t  p^���f#@�����A7��-��؃  ΋z<���c�#t��ВA7:  8/���{���&����k��xP-�pC  ��&b(q7���!�2��ߣCt�A����L&C�	  ���s�f#�n�g�A7��-��� �y5�M�qg� �A����# �xP�?�P @'�:�f#@7���fg�)q���t  p^��y,��� ���"�n�����Ƞ ���}�=�1A�8�9�cr��1k&����-}B4t��t  �$ax�0���!��¡KV6z�TJk��Z���GW��  ��,��;Q'ވ���O� ��Ǉ�K�  ^�h4���a>2�60���!���� =>T7�t:�L  �-t3���SU8�=z�n?�}��@��V���R�`i�  ^F=�!@���g���B����}�ԆS�`�� ���A��~<�G����tʦ��H$�?(�_f#@  gE=T����Sk �5<@g���J� ��Ƞ���H�<N�$�����V���g2��f  lQ�׵��l�l�f�ܣ
��Z�A�W�
�P�?�  �e�:�fSU8��A�W@D��"|XL@��l2�Tv�  ���<�
I2�fSe��Zl�K��"?	���DO�Ww��h4ʊ�� �6�g;�u�ec8J��`��hW� ��A��� �.��H��G�n��mJ܍���K���T+ᔧ �6U��6�̧��$)j�K�	�M��� @  �Ƞ�{��J����t>,�#@�U���fC�	  0�n������wq�!�n��P�h�� �6��P~�\��}_\�� ݗ���a���y�_�S�h)Q  m��J��q��1<�G�qS�<.�H]� ��DB����9�Q�V���i�Kk  @H<�czL�4�Sŋ����W���L����q�ٚͦ��7Y  ��tI�R,�N�]���͞����1�n�F�n>��  ���C�A'!j��Ƞ�H�Ǘ �|�C  *�mqm�棃�m'B�n&��899	����C�	  0��y�Mw$��J�o�!���+��x��U����4�3��ˍ  ��t;����S�6��@�n2��ZD�F @o�}_;�B��TM�Ƞ�!�XH��F�����D�z|T����4\�e?  =�^�+O}y�̠
�=2�vH����� �M�t���籠b8�Uqt  z�Y�����l�*���="�2C:c�bt�����[��'��z�(s �w�>�Q�n>�����J�'�0�I��t�)s7���q�un�  �.�sB��S%�Ȟ���s�OD���t��Ǉ�t���/��   �薸�`>U��h4B�	T�.��⿼���1�n�3%���9j�u��1   ~<ϣ�{�p�\����g���A7��0�����rዛ.  ����XkOr&��d��=��	t;$���/�t��ǋ*�N� @���Ny���J{����n���>�[�{v&��>t  �2���,�/�L*���!e���"|xL�N��K�Ȣ�O�BN� @�!��#�<�#�f��@�⿼'@���������Q��|>O�8  z��y��B�����U����t6�)t�9����?���S5�s��q  z��ёV��l6+���{f���T(�#�XL�P�: 3�身���*���8  �C�\���Ƞ���}SODhH�s�E�M�[�N�nt  �F�/�:�ǉz
����{:�S�n �d�#���FL�;  �C��� �|��A������/�t�6�<O��z3«8>>�k��d�@ ����ֳ���f�t:���}���Ʉ���_���D��z]�i��,��(s7�N������f  �rxx�5�P(pʋhg�.g�E� �BwՔ2w;�n��  �_�R��s����c��t5GV�����$S��=^� �n}``��3�EP�$>͑Q�W"@��n�F�n�9��K���  �5�M��6�qX���*@�A�9�Yc3蔸�B7�~ttD� �ܔY-  �t������n�q�{�I|���3�EȠ�C7��y��j�f�WE�;  ����x�f���=�#�i��@?�ݗ�� �Pg)o�Q�T7fn�  ���E�=���ɤ=�EN	��0�C�����3�EPݘ���L.�  ��l6�Z�*�9�Â�%(o�G2e������EN	�)�0��4t;4�M�{�M ��988�����O�XK��D&�i�Lƞq"��"|�LA=~TY�b��L  @Xt��y�t{�t���
��VS�z��{f������ܘ ��r��5�� ;����m����ln�����EH?@�+������i��������y^��L��  pF�jU+X;�s��ʞ7�M�A6H*��z
�̝����d��2�x�}�n�  �U�\[�X4�8(�@���X�������ɠ�C��I�lMDOu�i&  ��t��K�R�g����t @7��G����i:f�)�0z��n�⺧~5 �E<��~F#@��*�N��s��Ήȩw�(��f����:�u���j�g���K�;  1ppp�{��P(H:m�>Y� ��� �"�~z��B�ȏ�3��+�BAk,Yt{���^��  �Q�?:�ϩD6G.�GE����"�V��=~T�йQ `?�q,�ۃ��v1�2� �f�:���qxx(�f���t:�Q+  X���X+X�ot{8�cr_������2�Y2��؃,:  ���������(�4C�#���+� gϠ����B!�E[��
l>�� ���Ї���<\�\.���<�� �L&�)tr,"�.v��y��
�A؇?�ή}}}&��  ��ժ���(�%�INn���vɘ����k"�2��fS+�J�g���y������PH�  E7{>88(��ty6�(����d5K>olo����E:2s���Ba��   ����i��>oU�&���}_�Y�3��|��Q,��V�U*,�*s/
&  ^R�����X9.�HhoaD�2�L�3���<��u]�;��?@'�n�D"��G�}��h�ZʪV� ����ָR�dr ����?�4%s��F�q:�{�ѐV�u����Q�O�28�� `������.�I����c�\�.�*t>l&�='�Fqv)�ˁa�BA��l�3  �Q�մ�ۓ�$������N�Y򊊇��Z� t��v�<>>���"ts  vvv��Q�n�d2�<������}_��?{w��X�݉�q�����L��խReW�Z��eIo�j�!)l�
�#�,G�c(�~�ǖ�c�أ�3#OuWK�*n��	b�w�^�H�S�	�{��.���Q�}H�*� �}�s�O���@o�0bА��n�y8���ݓ��ЭE������̏��I��w��Rl�K��e���ϟL�-G�9t�Y2�r��N�3���QmNBDDDƩ�j�>7;�N�ri2�?��R�����o�N�����jTtv$4���lg-�,�Y��i���Fͼ�G}�MR↦�
$�����/_|nt8?����3��errRӋz�ZUܑ%��R��7t"""�e�N	:Y��nWl�+�2w�M&�z�s�n������	�w?18�/y��@Sw
>���n�k��.�2w�-�Z�*ށu8��JDDdB�b�v[u������!"z,j��y��|nnnn�^�e������kՍk=t�-Ҕ��l�\��:����u�]w"""��ڽ=�9zl�f-�n��fْ$�/���\N����PW[�)A��U��Hk��t���r�="�����v��iS�f����1A��j����7�M�o���[M����:řG(�(�����:�XL��V��"�܉��LD��zO8��n�!"z,n�N�s�u��2�^�ggx��ѼGS������EELLLhZ�2w�Q+�����)"""R���ѥe�����ruu�x������ȟ��%� ��͆��GW�XT����z9�����ժ���.�KS�_2����"�2�ɤ�d2�ˋ�"z�㕸<_a6Z���E�ٳY���d��.<���鴦u����j1� �&���4�N��)g}��u��=�-��nQ�@@q&cO���,��K-A�F�<�FDDd�n��|>��NNa� �ϧ����h�G�)�˚ֽ}s<�H�?,4tpsƟ�h}�/
C��[��R<��N�DDD��d2�>G"�FcdN�PH�:���GkEK:�1�����v�	:�]t�a�>��vѧ��u�����~���p|��&��y���5��%���w{M�;&�Sd.�h6����Z��ǂ�Ţb��ǣz6����_�\֔���n6�� �өx����GK�/��t��2��w��EE��a�u�,sݢ�������	��R)M��>mMj7U��&���L��T����:�7/�S��t�a��hK�ӊo �H.�Kǈ���ƛZ��Q155�CD��X�n=w-��������N�cāzR����P(pܚu�]�r�gd8r���H?�TJ�g�X,����I��~�5L������H    IDATN�u>&z��u�t�OH���|�z���ݮ��d.jet��Ӛz��H��霫 ,o��@ �xc��nߩ���qqq�y���@(41�hޣ��9�}$h�A�2��̧�h�T*�.�"�� �ɠ����<�fQʉs!�i�ۨ�4oPc~aA�ͭ���;GV�V��%4dZt�Ri2/�]�x<�S$DDD�K�e�[ϟ[��FV?��C�d���e�t�u���Ą����f�Nw��<J��b�F�ۭzǗ����P(hj����8Z͢|>����n���L���Z�Z�͆��>b4}7Ax��lA��,���֕L&�����	��Q{�r$4,,o����s�kwv�*WI<���w��{%�܅5���iM똠[W.�S��T���ݕ�eT*�un��pX��h��ۙ�O���<bME|���rD���;������D"����j���[�,˪gѹ�NDD�������B�!GC���x�v�^�$���&���Y�'_�%�UǏ�N���=�f�	I���4$6��e�c ��(�����x<:FDDD4�����:����*���]��J:�|�ln�����M_�$�,s݄���sܚuI���A�݉����͍�u�x\��M��t��������`�����x�I�>I�(�BE�u�JE�,3�[:�V�`�F���JDD��ͦ���ݮy�����r)V ʲ�#�&$I2���p8���?�S�B�L;jxu�/b�>BDQ�TZ%�2��-���(�����DDD����FSYs<״IB��؏���T�T.��+�������䤎Q}�+ wn\p��^���	i-o�f�C���)�L*��MMMq����Z���Q133�CD4,j	:7&�)�H���N����:��?����t��K�\� *į�j�d2�hv�]���n\H��dgQ�N�Tj���.��ɉΑ��D"�i3�����v���%Ib�-�e��Ϲ����/⓯�,9*tzw7����Zum6�e)���R)LMM�P055���k�!""�#�H$�x����Իq27?������am}èFp���>_����j���/�!���є�g2&���t��d6��x����FDDdqw�=7YB@w������x�_�W���a(���}��A� �ͦj)5�orr�Cu]�VcɎũ�E��b<�@DDt�fSS����Ѧ��z�v�^gy�y�A�CPs�p�/|�F��f�<��⬭�� �L�.���t�����ڮ��5�4������q�ܚdYF(�����u�x��O\sb7��J�+Y������;�z]��s��ɳ�#@��97"�I8�N��Pc\��'�9��aŒ��z�Ο��u�]���(�����)"""�Һ{>77�����@~�_1��v�l�kRn�%6����_��W�N��V���oC��� L�t:=�hh�2����a$��"""�j����Q�˅��)"�a��u�!�C��'���G���'�9i�О�f9>��$I�.:�\]]iZ�����s���l���03�1/$� R��b&�#���#T�p�n�5�1&s�d2��FC��j3""�qT(P.�U�y�^LNN���Ąb��f��v��cD�� Vm��C��Q�Z��X�����e�A�����"A�)"""�e��ך�.//�}t��ݺ�>��!hq��v��tI���ݤ��2�B����#�T*�T*���xxn�����鴦YבHDSe"����P�9ʲ̼��B�7WL�A	���T*��qGc�8LMM)����d�d22����x��f��vu�����|��.���:A����CD4ljG��:$I�)����H�l��Hc�		��<b��R󚝝UMЁww���[_�^G&�A4�{�n�cvv:GFDDd.777�*gff4��%�cs8�
�ÈF�X[[Ó'O�g�W �Z(x���V��L*�*�y�V�,��DB�����\.���K��D*��h�n�k��C���z������v�h4t���bii���xP�8�t�]�;���fc��1�n�K�l6K���h�]^^j*�]XX�B�h�`PuaO�Ze�k[]]5:-t�`�>6���N�R<w3"R������lvCDD�T*i1��z��t���ME��v�2��r��R�i��V�1�3)�׫:RxWړ��t���M�e���+��""7�$i�������g�7N42�x<ntZ4 |��o�	:�����uZ�c�5��e�Ł�=���u�����X�tZ�9�h4�J��V���ss���0:-~���o�	:�'���b1M��J�o������ʖ��yM�"""�S���#�"{������;�$I���:FDw!��x<�xp�8�	�X�K�8�V�������EQ�\]ADDde�v������x�z�LMM)^�T*lgb���V9j������N��;P&��Y\:�f?��L&����(B����T*!�ϫ��z�V9�J�9������V�L�>���.��٬��6��ن�@DDd(I�T��w��+++V٭#���,r�$��1��P�:��e�R2��⢦N�T�?�R�T��f��q�݈�㸺��92""��J$��G{b����^�����8�={��711aP4��=�G)?J��j��j�xvǤb��n�j�r��J��߯Sd4lWWW�B��������!���
��z��d2����tZe��4�������.?�����}������c}��ճ���a}kz A47��F���tw�A���~Q�`��ˊ��d=j���r���L�����!he���"�6??��M(�͢�n��%�͢T*���t����h8�鴦Ϥ�pXS���áX
-�2��������1:-� �������z��;R&�t:133��N�$�\A���QyD���,��ji�"��UJh������U�UN,2�o|�F���O���e3��涴��i]2��͖�j�p}}=�(�X]]�1"""��uvv�����2oJ�A6���q\�����gtZ=Zy;0�������չ���dNK�w��L&���
��ş��,)��(�Ꙙ��{��D"p8�7�M�4�H$�`0htZY'A�$��*LNk�қ��!GBF8;;S������]""��V����K�u�]Z�Ñ�=�����G��͆����~8쇠��bp�\����2�ժ������\Y����ބMj��:�G���,���_�5�����z��;z���'��!�l6���Db�ѐ��4�������NDD��N�5��G"������i���f~;z���	��g�
���0� ��������,�ͦ��Ժ�/--��v���4�MM�����a#��r)��$�"������]X/AE�jgƎ(�XXXP]'�2w�GT��������6�kkk:FDDD��,�899�Ե}uuU��Y���y�R�)��e���atw���=A,wd,-..�fS:�R)ŝV��B��|>?�����쬎i�H$4��b1Ml�z�v;"����,�9�D�Qş�ɔ �|�o�K����c���c��v#����$	�TJ������h�Z����������j��iڌ�������"C�b1�ͦj����˿��F�p�x�'�.	� lgZߴ�˃FT�������� `}}�(�� �$���T��W��KK� Y��fC4U\��sk�P�v �������J�����~�����v�LF����JE�׀��������h�����h4T�-,,����!�*6<���h��:FD�����.��0��n	���fff�z8����sD��J$�T*�OMM�ީ&""�L&�\.��.
���Aud���{d�o��F�pu ;�o�k����/�hj�R��������(6\^^��5""2D����Ņ�:���)$#.��t��l69&�"�����]|
`(O,]t��[��٠Zf��u��m����.�"���!��QѸ�$	o޼Q��;w������U��E�"��������5:��Jy;�s�������9=��ajj
�`Pu]�V�.��+��]�}>ϣ��...P��U����!
�%+V�Z-M=
�x��+�btw�����������I�����iw�G��Օ�y���i�G'""]�r9M�j�� 7�� w�G� �ַ�etw��ٰ���	����-������iM�N��*_�F�,�x���b����ex<�""�qS���^�8�Nlll�ֈ���P���j�4UZ��677�r���.~`h��gʑH���z?,֦݃*�E}�NGq>�(�����|t""
I����[M��766�p8t�����{�����[��[F�pWC;���k�?�������Tו�e���r�������n��1}DDDwqzz��,�����(�=�Aņb�v�ZMǈ�\.�����F/A��9�a-@�E�/���Ql�FU�h݅�{OO4E<�!"2Ϟ���>��j�QZxW�>4�$�.���Mw��5�J%���3�]���EMS ���ԔJ%���׫yS��-*�I��uȲl���� �	fX�6�u�[� h>�~qq1�h�z�g;�N���k�ADD&�j�prrY����vlmm�	�P����uX��r��퀁	��'O0==m������h:�U.���8&��&NNN^�������%""�I�p||<�fp� V� M�411�X���sk����gt����~ �>=�����]t�\.���j�u��}���j�����cUcDm��P(�	=� ��_�U�ø��O�� �no}��߶ZS��5==�P(���R� ����A2�T�yONNbvvVǈ��������p�X̊�tO�H�s�G��ʊ�����?�MЧ�����mdt����]^^����qvv�r�<����&''u�����*��kj
9�s̨݌���?0:����z<��D����i�F�U��j5Y�qrr�f�9p���b�U""�Z����S�u��}N����$�n����fSq������/��/�}�+=��W�O>��������i����c���(vv��l��NDD�Z-C�$�u���v�]���h� p�|�|�߰�1�����@�'�N��v��0H�p8���)�u�F�tZ���,�NOOޘq:���؀(�:GFDDf��vq||��y�f�assSq'�FO4U��_�����|,8�x׽�����`�n1�����z]^^��	��R*�;��|>lllX�)�,�x�����^+++��>fl6w�G���""���a܇.���$�$qf����~��ͩ�k�ZH$:DDf��d�P��׈���F��RIu��⢦
>-�x�c��J�>��hs8@���It�w��fmmMS����Z����$	d�فףѨ��<DD4�����+zb�Gv�!�өxSF�$�E#��r�\x����a���C��4	z�\F��KY?=�ۍ��%�u�$���J���l����8���1==�cDDDd�L777����0VVVt���fvvV�S?s���׿n�c��R�3M�.˲�'2���U8�N�u�TJ��2=�����W���011�cDDDd�B����s�u�@�}KƔ��U<���vQ.�u����C�C�/�Ο&J���[�(�X[[S]'˲b�0]�μ�f�
�����##""#T*�����b�z������1�v�X,���,,,X�9���|@S��5�M�Z����~��\.�
�1��tp||<���f���|>�Α������Y�n���ۜu>������v��j��cD�~�7���� Rz>��t���V������\��9��V����#t:���EQ���g���F����C�3�N�O�<�t��F� ���B��'-��r��?6:�����~@�%�Ri��x2�X,�h4���R� ����Q�������g����p�\:GFDD��n�o�������1�F��x^��묶��o~�V�%�]�e�L����-M�x�9���:޼y3����rakkKq�)YG�������UQ���x�^�"#�E�x|�uY����u��������}�|����.A�|>������X\\T]�j�8vm�U*�}�v`���xx���ht:l���E�������Y���r��*[��ٱ�������AM��w:T*�à;Z[[�tf���F�͚F[�TR�I�z���ކ(�:GFDD�������H��f�a{{�`P��Ȍ�n��qII��l؂dY����C�^��4A�u�&kq8��I����3""3+��x����j�χ'O�p'���bz�y�VS\g�ٰ���䜰���xT2��s���b1����C�K#Դ	z�^G.ώ�V377��6�ϳc?�T*)����|����N:�EH��7oި���%��pX��Ȭ&&&Ǫ�Z-�U�����F��� ����M�����!�	����-Mk����k�P(�t���$���z;��rYq�s��l�c��Κ�N'��o�C����	���5ͦ�a�E"�.�=�z�DB����Ԓ�@ �3�DD&�K��z�l6lnn29' �J����U�U4�X�w���l�N5��s�����$I��٥�a�=lmmi:;|yy�^�.IWj���y&��Ȅzɹ�����-LLL�����������$q�ܢA�o��o�C� �;���	: �99gSr�\lGw�����v�^��|�FDd"�v�����m�B!�"#����W�a-
�,jgg>���0���2��M���\%�F�A������8���)��uwWJҟ<y�ásdDD�E�v[�(5Q���vk�[�pX�3b����e��e��lt���O�`�Ȑz�@� `ggGqlF���	�ҭr����#t:��׽^/vwwϭ��Z-�&������]�i������㖭kvv���F��]� �H�^(���d���!baaAu]����%��P��pxx�v����������^�Α��z�����2N��������Y8�΁�K�Z-ê��������S #�D� G'F�@�����ۭ�.�H�V��YE��P�������u���h<U�U�&P�{{{�x<:EFV��z1555�z��E�T�1"zL�`_��W��-o,��ߤ�(�kEv�]�ltY�qr�1�eje��(b{{�g����\.���p���χ���]ROjU��|�G-���{��c� ߜ���̌�Ӟr��T*�CDd%�N���ƈ����-D"�##"�|��Ǫ�S(���y�{b��bg�z��JJs:���w�kt��+���T�~q�@M�	���Ύ��Xggg<{D�������f�acc�x\�Ȉ�F[*����ujj
���EQ���*�N����$Ilgq��뿮86�"�=,��K����F�A��v���������ԝ�������fqqKKK:FED4����pqqY�����`uuU��?����7n
����d~�(�?���a<�ϟK�����m�Od^���ʐ��<�Yv����������`ccc��B�$�}�V�(�n����
�����S_����}b��&g�[�׿��Q�9Q�o��`���t�����0�z�ѵ������6���Vr�D�����X��NG�HQ��f���&���u����n�c~~~�uY��!cq� ��h5t���gl-���ћSvx�0�χ��5�u�v�����,+�����h��`0���]Mc�����n����ꎦ�����.��N��i)m�f�����"ƃu�ݿ4:�K&��Fg�F�A����i,V&�Q��O�Z�b`�W�ۍ��=�a#"RQ.����k4�u^�{{{���B�&&&^o�Z(��:FD��'�'F��`�V?������q�X2A���7�KȼA��ޞ�3�'''lB���6���P*��^��J�� -    IDAT2ꏈhe2���F"����yS"Q���8�,���>FezΏ~�#�ٟ�Y���l�^��pq�0:z�@ ���U�u�Vggg:DDV��vq||�T*��� X]]��Α��,˸����ٙ�����,p�&���p8��J%�Ե8Y����F��(���������ݓ^���\�]C-luu�t�bQq]*�B(���N��U]^^�V�aqq�����Yx�^�y��ވh�u:����>��lXYYai211�؛��j�~�#�����+��xL�Q�\�U"����C�{O�>ŧ�~�ZVwzz�`0�xG� r��VWW��aNLL`ww������DHDd�z��7oޠ�l*�s:�����ys��n�����k��ɲ��������O��ј�؎�k�^��,���|>lll��k��899�!"�Z���;��n���"����
�T��`0��O�29'͖��Ǜ�����W�:j��j3I�?S젯���m���5%ߍF�(Y���"R��jÐ\.�L&�h4�Sdde�Y�}�3�(bcc������2 B""�Ȳ���k��ܨ����X\\�1B�,�*NLi4����	�&S$���?99�����s'��A��g��7�7��ONNMU�B�%�2���Q�T�K���G0���1���H��y�5�|�;q�\���x]�$����z���Cf�w XYY�|`t�@.�[[[���.޼y�CD4Jr�����d�A��������pU�U�~�Z59�x<���crNw6�xO>����Ы¡�� ~�w������#���+�H&�:DD���h��� �|��u�Ӊ��LOO��p$�I����F�x��)�^�N�Ѩ����{T��V��Z��K��D�V3:��72	������������n��ggg|��;�v�899���e�c1� `yy���Eр���Wm6赮�7Bm}}����μ^/fgg^�v�����:x�\#�J�����F�@���p��ӧ��i$I���1$I�)2%�TJ�����$�>}ʒw"��^I{�PP\�+ig��G����l6��i#�^��ɟNF*A����W��U�àG�D������V����|��H��jx������.�;;;����92"��I�R8<<T�655Œvz����\��׋�"Gq��=��H%� ��	2"666011������Sto�$������}�����yloosr �V�����...w,{�%���X�N���	�Z-�E#�a��j<V���{e^YY���ύ�� x��)�v�i�o߾Um�C�$�����`�P(���.B��Α)+����<{��]��A�N'^�$	�LFǈhظ{���K���~��xWxDx�^���t:8>>Vl�C��������s��tb{{+++|�!"�I������n\׫���Q,I&R�k���y�����tt����Z�r��Է&������w��M����fff�N�U�ޕJ%$	�n�DjdYF2�D�R���R�בX,�`0���c��!"CT*�����5�z�X__�Ysz�x\�yj�Ze)􈹺�2:��3�]�$d��a>�@�R	���<�>"vvvP*�T�G^\\���#���j����}�����n7vww�H$T�=Y��J�V�|Q,���2+~�Q�����n��hĔ�e՛���F���n�9�E|���\jY�UK����$	WWW8>>���@���bww��SD4t�z����7�n7vvv��������������s�Y=Z�{n��~���h����Σ�Z-�gO��T*�իWH&�}��|>���aaa�U;D��zGo���Uˇc��={�J2z4� `eeE��y>���Ȉ)�J��d��N��|>ot���8���UוJ%���G��M?<<�;׵�������g@�D4���:^�~���K��i�5�aQ;w^�T؏e�Ȳ����W�l6���Fֳ���@ ��������U*���#�J��ޛ<��t"zI�pyy�ׯ_+vP���9C(R<w�j��6�
�;�h��n�kX�:Q�|Eu>z�<:��c�}pTn��D��J�_�F2�T<��;^����]sztN�KKK����h�$	�D��0��X���r9��1^�{{{����6ϣ���j5,=u��x��	666�p8������n���}��􈢈��e����r���GS&�A��5:��6	�,��EA���X^^V]W.�q~~>��h,�F�|�r`�_$��g���t����"���իW��W��0>���������͟R��y�#���<�G��t3)
��p�\F�B�hss�RIu�f"����C4�)27�v'''��󘛛{��n�cee���8;;�"�����JEq������2&&&t���U4U���h4P(t���rssêS���t:mt��A�W��x<յo߾e�Q�B��ׯ_���o�X0�ӧO�����G��FW���������s�͆��y<{���9���������N�LFǈH/l�gc��s�hr8��W��� G�$��$IH&�x�����h4��|�+��q�h��ݽx��TJq��W�>??�&p4t�����NȲ�L&��H#�����蟌ݫ}:�f��
���U]�l6q||�� ������o�'Q������=��D4��2^�~���S��Z^�;;;�����<�E�)�RC�\.��8#�Z�r�D�.Ao4(��F�AC0;;�8��X,���B����)��x�����>��������q��l6���[*�4w:�X]]�ӧO9��t5??�x��T*1�Q�,�����0��� d*�B `������r���4���>����:EF�n��P(`zz�����aLLL �L����k�,���"�H �N+��l6���`nn�(�!ѻI#SSS�7�E#"=��eű����L�;���<"��ѡ�#|�~��)�R ��7o��x��zu������D"�l6�����^�A�����(.//UϨ��H��t:����m� `jj
���p:�:FH��������뽦p|M�$�����0��O�>��8�͆��UvQQ�J?��Uw �N'�������v�����^o�Z����\R"�e�BWWWh6��kC����x���t:���9�3P��)�뎮ލD�N��o��oM�d�x���Ǎ��$�������U������C.���avv�@���z����K��Dd�r������@ ���Ł��DzE����cj���󙬫��`����	��,//��v������U�E"lnn���`0���ف�j�J(�J:GFD��J%\__�6����X\\d�72���5�B�����<�*����s��3%�c_�}ss���%6�QKKK�V��]�s�.//1??�SdD��J%�J%��ͽ����~<y��r���(
EJ4�*�
���U��ߏ�����X��6??���W*&�#�^�397��O�{c�xG{tmoo�Z���_^^��v#���`�r����@ p;���:�~�&�@ ���L��T&''��^o4���:FDz�e��Mn�K��n�cee��MFX��Ə�c�D�͆���Y�DF������|}���e\^^���hH��"nnnP�T��J"#��~lll�m��H&��#����<.//��t�T����LNN*΀$��j���V�����p`oo.�K�Ȉ�������X�S�Vq}}�frD�@�e��y��ܨ6�
�Ê����r����5pz�$I�c����.���y�&�&$VVV8nk��E��'?A��U\�v�����áSdDw��x0==�p8�w7��l����T�o�Dw$I�mb�h4��h�x���ȴ�v;���n<Ȳ�T*�:������l��0L�	�I��~6	�d����:V"�ɓ'�F��r����D��i�Z���ڍ)�q��t�N��N�g?���X,�x<��dj�(bccC�ǩ��V����C�U�	��-,,<�I����/_�T]�����.�dz�(�6��0Ȳ�l6�D"�Z�f@�D��h4�N���d+N\.������
�	ǩQ�۷oU{1�33%�|w�9�d����5q����j899Q\���qzz����"#��n��T*�T*�P(�X,�����R�h4���D��\.#�L����|���A4�[������X,29�R�ɹ�0A�9�V�\�������&����d2	�˅��Y�"#z�b��b��׋h4�H$򥛎�m�z�T
�L���hlt:d�Y��i�3��("�bzz����r��b��j��9�cB�$vm�&�}d�Y�A�+{{{h�Z�3����p8��,�V����WWW�Ø����㹽��x������E��y�R)~`��U�ՐN������=���X�N����^o6���1F��${�XϠ��z���ht��N���>�L���f�a{{{�x+"+����F�����{��Z�"�J!����,���"�˩6���l������4�~��=�`0�����G1Z��{��F����#�ð3�Ag��`vv��ؘh�Z���T���l6<y�sn��DQD(���d��$I(
H��<�N�"�2��*�٬�n������4&''�NA ��χ����}�:�wSǈ,�x��;�k��"�v;VWW�0nL��u|��g�3o�wϋ���I���v�199���ɾ%��FCә]"#5�Md�Yd2�iN��h�Xn�[������`ccc�&��'�������0,�	����aLOO�Z���>C��R\�t:����˥SdD�����D"��}w��*2�ˑ)t:�Ed�Y�cJ�("� �`bb���i�8�NlooL�%IB2�T�qE��������G�	������%�e#�b?��OT�2��n��찙 �$�͆@ �p8<�z�XD&�A>���F��ۤ�T*A�����l�B�D"���d5�$�Á��́�,#�L�n<�h9??g��;b�n1n����F�A:��r����;�;�^����<�H#MELLL`bb�@�D�w^=�͢P(��==�n��b��|>�R�4�9f��011�XB4*�v;677n"ɲ�t:�zt�FK�VÛ7o��r��[���4���a��R�~���ܝ�	x��	wgh,���v7s�w��A��.
���"�ŢbR��)�D"L�i,�l6���+N�d2��j:FEF�e<�pL�-�f�aee���PHG���x��j�>11���M&�4Vl6�� �� B��{���,�X,�P(�P(���j6��ϙJ�2���tbbb�p�P���4Vl6���'�d�Y��44z��$R���aX�����$�=�$!�Hp6������,�x��b�^(pxx�$��J���7���v#
!
���C���x�]���Q(����e�z�v�|�n� �z��B��uIcK���*��r9&�c��l29�A��x<�P(dt�����z�Ju]$���;�س����`��½�ۥR	�B���H��D�\F�XD�\x��t����W�A4nA�������5�\�JEǨ�dY���1�< w�-,�L���eA�iaa�$a_q].����1��י��X�t:��r��r ����������ׁw��{g�K�Ϯ��N��r��r��R�4�(���%�� �^�Α�� XYYQL���<��1��d���f�wԛ%977gt(����% PMҳ�, 0I'��z��z��d2	�����χ`0���ۍ������]�R�ę��n�Q�VQ�TP.�Q���gE~��P�@ >��G��XZZ�=.�O�P@�\�1"2�v�}��J��	�=�vxn�,--������Hq]6��(�XYYa�N�G�V��y�/&�>����X�v}�\F�RA�R�N��4�ۄ\�g�r�n+(�� <_�4X^^F$x��׃����9{��&���L&��z9�e���B�$���F���z�Edi?������d�����������w:�ۄ�R��Z�r�]�N�j�K�GE>��6!���<CNtKKK��y�ʈ�S.��(����:���4fff�����Qqxx�����s'��nzM����s8�z��|>ߗJ>[��m��+����F�?Z�j���&��:j�Z���v�����J���yD���tۧ��R����H/�N���F�AC��
���9?+++ �)I�e�����J� �v�����z<��s��x�������&��Z�F�Z���_�n��h4P���h4n����x�3���������8�#Au�e��M�e\\\��}D1A��������͘��(�K�ӐekkkL҉�;�Q/qw�\�� \.DQD���RB�l6�l6�h4F��|��E��@��z���7+DQ���B(����v����D,//#\����n��z��hb��@�v�T���clyy6��_�V\��d I��`P��+�w:���n7����?˲|����m4�M�Z��6��vY�o���������/�w��~LNN��r��t��r1	'2Po��R�v&���tpqqat4DL�A�P�m�C�iqq6��^�R,7��r8::���:�.��n�oG��#l6�v;\.�v;�^/� �v�m��,ːe�$����n�����������,��v�_�>_��v�}�}%I���^\v���z ��p��p�n���p�� �I�l6��� 
\���k:�z���ML�I�ԝ]�����<A�˗/5%�L҉L�Ir�ټ��J�Y�!����� �e�_\#I����ݍ����Qo����h��lX[[Sߛ�f�T����y�f0A$�N777���3:2���l6^�x�xw3����� [[[��M4B�����m"R#�"���Vaʲ�l6�QZ�V��D"at�~zxD�r�5	�x~��j5E�XīW��M���h�����u��<�N39'Ȳ���s���	&����	!�࣏>Rm�T�T���K�5�"""��q:����8�W�$�R)4�##3�d2���F�A:a���$Ib�	 B��?�ۭ��^���˗|&""n����p�\}�w�]�R�;�����j�pssct�#&�CP�VQ,��L��������z����&^�|�26""���z���	����z��A2�dexW�~zzjt�3&�C�W��x<x���bwV��觗/_r�)�
��؀�޿Gs��F2��QI��J���}HX�N_�r���G)�7ޕ��~��BA�Ȉ��h�&&&���6��l��D2���HT�בJ����}���:2���a�I8|��G���V\'I�L&u������%�beee���Z��T*��tK�$���1&�C�ٕ�E�(�>���:Y�qrr���s�"#""���Ǳ��A�^�T*�f��eY��ȬdY���%�:�1&�C&�2�K�� ��������7���k�y�o�DDD"������)���r|��/)�l6=映��ns<�gii	{{{K�z��4���y�����l6����D�^�e�L�I���j�����0�`L�uR.��BL�Ň~8��kO�X�˗/9�����677�^�$	�T���=�,��쌽�	��8z���D"x��9�n��Z���/_�^��i��x�������z��E2���,�����F��0����H�$\__��'��?V��l6�����y�"#"""5�`���p8}�7�M��ܠ�n�YA�Z��'��]g�F�t��0Ȅz�ҕ� ������	�b1����q���^2�O����ٙ�a��0A7@>�G�Z5:2!Q���3���)��e���x��-+2��� 0???pM�TB&��{5�%�2���y󆾄	�dY���5��@������ލ�I�R��NDD�3Q���������eYF6�E�P�92��L&�J�btd2L���vq}}mtdb333��_�E�\.�u�b��9����rakk�@���^38VK��!�    IDAT�F����t�j5�G'E���~�i4x��J��N���@ ���큓WZ�����n���o��t�e�Y���"�ۍ�}�k���U\��t���kVfA4UlW�V�L&y�����x"����n�"Q���S����f�k�k6r||I�t����h4�l6,//cqq� �]S(��f��Te2 EL�M������/�j~~~�!�N��L&�/^��l���q:����D$�{]�$�R)1#M��*ϝ�*&�&�h4�J���, ���O>A0T\W������C�=��~loo������j�pss�&��	睓VL�M$�ϣ\.Y�������177����҉���.�bccv����Z���椙,�8==�sҤ��&�H��r��0�����=��~<s�;�^�ױ���x����h������E����eYF�P��
�I*�B�V3:�~R7I�puu�_����2�?�ǣ�.�N���?�Qn�[[[��N��T*���\.�+�	tj6�H$F�A
���'� �*����x���(���� �(�7��븹�a�U��V��s�tgL�M�\.#��Y�����~����c`�wUo߾ś7oX�ADDc�f�aqq������E��i�gҝ�>oqJ�Ϡ�X:������3:����%��?����t:�j����́;DDD���vceee�1I���dإ��L�e\\\��n
Yw�ML�e\__��j
YLo۠st=�Ql�� "�q����=09o4H$L��^2���ҽ1A7�n�˦qt/.�}����;�w�]�䝈�F��f������&�,�X,"�Jq$�K�\��͍�a��1A��f��_t�A�����ϟ���*�e�w""e�[[[��b}�����E�#�Q��p���[D�Tb2�[��{<W\����BDD4Jb��bI{�Vc�vz6�����BR��ժ�a�E��v<{�O�>�(��I����S�~��������v;���0??�w,���r�d2<�E�&�2�����t�����/?=���,~�~	���">��s
�"#""z<�@ O�<A(�{��j!�H�R����t:�r�lt4"��[L�����%��҃x<|��GXYYQ���n�qpp���s>爈�l6�������uY�Q*�pss�N�c@�4JJ��ɤ�a�a�nA�fWWWF�Ag�ٰ����}�k��|�����x�G,���Լ^/���155��z����14����&�U�����y|\U�?�ϝ=�d�dO
݀���Zm����XE�VA@6iYd/(� ����RE�M�#�}�B��k�ɞ�2[f�{~��̝4)ɬ���Ws�=3�R�7�{�9�3����x�A) T@�`��.����0��,�BDD	E�$�����#���`P��t:����Bp4#� ��Ѭ��; :t�����t]KLt0j�.Daa!��x��F��v;�͛�.Q�v�aQ�����qd��Bۃ�`�C���$����i�4c
�r�JTVVN���t���===|rLDDqSTT�#�<2jr�r������fL�b;gb�la��zzz���F���>K�,�^���O�e��f�ٳ�����(��z=.\���j�T����`����>�f\?+�Ӭb���� :;;9͆fTII	�=�؃����v���q4���f�$I(..�QG�Ѩ�'4j�r�b����X,�x�A)�	z�������b�D3*4���/~1j��?���!""�Y����#�8������
�5���v�����0(0AO!n���0Ҭ(**�q�7�J��7���fL�B�dk͝N'����9%�<�~?�����	VqO1V��EEE��RLh����b�ڵN�S�_�һ�j�ܹs�NA$"":���,̙3'�,�@ ���a&�4k�� ZZZ���b�#�)hppV�5�aP����Ê+0w�\�)�!.��v�BGGGӉ�hZ�j5�����k.���fCoo/�s�5�,���~�?ޡP�z����V�EVVV�C��V��`�TTT`���R�'�@oo/���PUU���H��(���梪�
:�N�������&�U���X[�bM���aU��R�P]]=iq/�����?������q�a�M�}�'�N���j���(���Z��qd��z{{188�0(Ft:�nǎ	�ԏ#�)L�etuuaΜ9�j���RXII	
�����u7����l6������|�)�DD�B[����E��0::���.��Y'�����s�����^���j���x�Bi�n�c��ݰ�l��38��Ñ���Ȉ�(�dgg���*�l?�χ��a�|�GF��n����#�aP�%�:�4a00gΜI��"�)Btvv�����kM&Ӥk��(��t:TTT ??_�,˰�lp81��ҙ��BKKK�à8H��S�ӄ��Aww7*++�
�I�P]]���2���L:��b�`hh��މ�ҀJ���d:�tv���m�(�|>�:����4�������x�Ai��tb߾}]�e0P]]����EFDD�������ʨ�B�^/FFF8��b.`���|(��8�Nq322�Z����x�Bi�h4�_�"�w�^��n�~����GNN;�0dff�8R""�i������N	)�����9%&�ihpp*����s���(**Bkk+��ڢV���hhh@ii)*++Y���(	i4����d2)�B�יG[E4�dYFkk�A����4500 �Z�
�s*�
���Gee%ZZZ��ݭxc&�@oo/,���QZZ���DDI@�$�L&���B�Q���:s�7!�����x�
�8\���$IBEE�Fc�C�4�t:��܌���I��t:TUUE�!"�����Gyyy�u��###���B�l6�n��;J���	z��$	UUU\�Kq7<<��{�tK�ш���k��(����PYY���,��~�V�5j�X������H�à���Z�FUUC�C!B?���wЛ���\̙3������`0���,�~��`6�N�3Ƒ)����b�w�`��S�Q�՘3gt:]�C!B0��lF{{�����9VVV�KDC:�eee(,,T<�p8X ���bA___�à���F���9s��j�
��$꭭�Q��T*1Q'"�e�%%%0�L��;�p8���Qw� �5!�������P(A1A�����P]]��*Q<��~ttt���㠉zii)����&"�AL�)�Y�Vtvv�;J`L�)�1I�D��������<��<j�%%%�����DD��Z�FQQJKK��B����f�q�4JH6�f�9�aP�c�N	O�ף����%$�ǃ�����L:R��jQVV�=ԉ��I�V�d2���$jb�t:a�ۙ�S²��0�ͬ�@�����`@UU�tJX^�7<�}�D]�Ѡ��eee�<MB�R�d2qĜ����@{{{�à$���FFF*++��PB��|0��]����5�DD�i4�L&�L&��#G�)�8�N����;J"L�)�ddd����S�)�M5QW�T(..Fyy9��QZ%���Ŝ�N)attmmm��N�����tJ&~�f�f�y�}�U*JJJPVV�D��ҊN�Cqq1����˲����ɪ�4�n7ZZZ��Ӵ1A��������
&�4dYF__Z[[1::��$I���Gyy9�Fc#$"������� ??�$E�p8p:�Lr(���n����&蔴���PYY��K�(Q	!`�X�����:i���l���#???F��>�ш�����*���|p8�>�$JT����|�D��	:%5&��FFF��с���I�gff���EEE��QR�$	yyy())Aff�b��������f���L`�NI/33�����NI��t�������>���())��0Q�	�a^TT�X_C�e�\.8��	q?JtH8��f
tJ	,G� ���p��Q��T*���,�HQ<���pb���9��t���Vk����R��`@UUG)�	!0<<���X,�I�fgg���,j�%"�X���Fqqq���^��n�����Ӊ��v~�i�$R���w ��<:;;��Sғ$	���(,,����l�:���p��p@�ף��4���DD�E�V���&�Iq������N)��t���-�a���ӌ�H:��@ ���>��f8���T*U�S�,"��������"(Nc����4vJI������RP"��3A����QUU��3(���vtvv��\FFL&����o��f�Z�F~~>L&222"�!�v��t:Y��R��n��l�v�L�)e�t:TWW31���Qu"���x e������P(�1A����jQUU��&�(��l6tww���o�5����0�L(,,�"��V�Eaa!


`0"·�Hs:���|q��(vB\{zz�
�8&��4�������
Ѭ�e�������b�:�%IrrrPTT���BnQHD \���PPP�����!<FGG�r�8ŗ���� �����&��j5*++���*�ߏ��~tvv�n�G�V�QPP���"N�'JS���(((@AA��Ұ�����Ik_�!z{{144�P(M0A���R�PQQ����x�Bs�===��뛴pSFFFxT]iJ+������<*�2�o���Ugg'�Vk�à4��Ҋ$I(//Gvvv�C!�!�V+���������ohD�d2q�Q��j����G^^�Fc�yY��v�1::�*�ք��蘴+�l`�Ni����Sy)�M�{{{�y�$	F�1\,��划�F�ANN
P��r�������,�hoo���h�C�4���Vqq1


�QB�e�@ P�*.WXX���|h��GJDS��h������<���D���{<{#�L0Dkk+g�P�$R��ͪ)�a2��
QܩT*������d��z������6��$!33���(**�u�8��t���Cnn.�FcD�`0��ä�(�@ ���nH���S\��塴�4�a%$!���7�t�К���|c$�������pR>Q�Л�嚴�Q���|hii�:��(Vi�	:�MVV***�4�A8�b��j�F�3�BT�����E4CT*�F#rss���Q�Q���������DS�r����Y��
t������J��_�(R0���,���S�T���F~~>���V����pR�V�ǝ��z�ᤜI�Ԅf���f.�����h�V���*&D�$���n'�v�=��Nfff�xUvvv�:Y�t�9!''����B���n���e��������w(D�0A'�@�V�����(i�AX�Vahhv�]�_ht=��633�	;�%�^���ldgg+��x<��Gɉ�}}}�w(D)A�bJ�`f�eee�[�����j��� ��za�Z1888n:�,������*QO\_K�*�Z-�Fc���-C��C���`0N��!�fs��D�L�)a!��Ӄ`0����x�C���z}x7 p:��Z����p8a������0��!B����ٜ�BI�`0�h4��&.�
�z�ᤜ���f^0D{{;\.W�C!J
L�)������󡸸��n�fP(I������������p@��k�X �u���FVV+�SB
%������)롤�	9�����hii��D������� ��˙�͒�#�~�V�5<��f���������x��T����F�1b�0�l�j����DVV������9n�,��bn>�^��kȉb��v������E�(�TTT��(N<�v;�V+�V+�v��\�NN�B��e���R����9�kb�u����|�#�#�͆��Nn�FI�E∦��񠣣���7cD4�����t:����p8��(eh�]�$ddd�G6CN�rL4�F�AFF233��������l*Y�����p8���ß="�?!����P���(��p�����x�C��T*rrr"v[p��I���(
i����z.eIC�$A�Ӆ�ПcgL��~���p2�u�D�I�etuu�w!�C����,����FQQ����M��g��u�\��������Fځ�Dml��i��/��74#4"n0�R� �@0���?�	�>��X��������P��tJ*�����|(--�;Q�S�T�"rcML�C#�.�V�5��I��^?.����0��t�$��I�N��^������ ���F�}>FGG��D���^/Z[[9��h�0A��]���W����C��8��{<�p���x<���,��0���P�V�e?�$I�V������}�A�A��6�-|��p���t:�����D3�	:%%��.����͐�պ�!��z�{Y��l��|p�\�z��Z�F�V�^N(�Z�/�F�։�J��F�	�]���}��%IB0�,�����Ѩ���(u���a�NI��󡽽���҈$I��[�;��V���r���#�G�eY�Z��J��Z����h�����W��
��=|���^��qf-�ց�]�}ÉHI�.��j�w(D)�	:%��/���B�L�x�CD	$��fee��� ��$>4rJZC�}M$��,�㶔�$	�$�K�C�s(y�f��+����ض����Pl�?�.��fJ @[[<O�C!JYL�)%��񠼼��҉hF����~���G�^�#�D�h\.���x}"�e�G4CFGG������P����R�CCChmmerNL�)��|>ttt��p�;"""��&�2:;;����J�D1��RNh]��b�w(DDDDI)���6�-ޡ��A���u�DDDD�Z6�-�b�#��FGG������P���������LΉ�	:�<���ٌ���x�BDDD���� :::����P����SZB``` n�eee�}�����ҝ��A[[�@�C!J{L�)�8x�^TTT@���;"""��Boo/��%#R�	m�f�Z�
Q\�A���s5��tJK�,���.�eee�$)�!ń��A{{;�~�C!�	��SZ����z�(//�w"""Jy###����9Q��wJ{^�f�6�-ޡ͊P����.&�D	�#�D8�K���N��Uމ��(���n����J;Q`�N4�����AYY233���288���>��%	&�D��~��f���(��M[ @{{;�nw�C!�i`�N��� �n7��ʠ��
%>!�N'�f3dY�w8D4M\hK4���Q����n��;"""�Iɲ������39'JRLRYYY��ͅJ���`�N�p���t: N�V�5�a���/;�Ӊ��R�#""����z������PR�J�Bnn.���  ��ِ$	���{�׋`0���e��0AOPeeeX�`���QQQ���
���#??yyy�j�SzY�a�Za�Z��ۋ��n������������i�^VV���p���� ���C��h0w�\̟?���(//GEEJJJ�������)�����j���zzz���mmmhjj����,��P��jjjX�1�


p�1�`�ҥ�����������z��܌]�va�Ν���EwwwL~v2+,,DQQQ��)�ti4^C��s���������4I���s�ￏ:�(̝;7f5�����o�>��Յ�B3`)>t:�nǎ�x�0A��^�/~�8��c�r�J~���i���lݺ[�n�����p8�RB���M'�C����V�����>m�����r�J{�X�brss�R�,�ػw/�n݊>� uuu��cL�Ӑ^�����3�8�|�$u�`;v���o����\�>�J�Baa!
�
%&�Dt(� :;;9�:���8���q�g`ѢEIs͵�lx����[o��?D0�wH)�	z������;��r
233����}�vl޼��׿�R����@YYY�X�G���    IDAT�0A'����������$222p�g��s���%K��:k�Z���������pR�g4q�9����ϟ���###������ �V+����t:�t:!�2��ej�:CVVV����dBEEL&ӌ\�����W^aQ�ϨT*O���/&�D4U�`��ݰ�l�%a͛7���wp�Yg�h4~������Gww7�E�].FGG��Z��V�a4���.*WZZ�����-��ЀW_}���Y��1AOQ�����q�����p������CSS���g���N�Cyy9,X����Aqq�!�_ ��o��^x{�왑���hDiii�
�Qrb�NDS�p8���$�/_�իWc�ʕ�|M5��ؽ{7�������뛱����٘3g.\���#���G����Cz���A����ظq#���&�)���?����o|#<�=U6�۷oǇ~��;w���-.���r,Y�˖-ñ�����i��֭[�~�z466�B�Ʌ��Dt0LЉh2�`===L��X�r%���Z,Z�hگmkk�֭[�c�����e�3�Z�#�<K�,��+�|��iרr��x饗�����s�91AO&�	?��p�9�Ly_r ����[o����_����NB. ��$iH1�	 b��"@�$IE ��a��ϟ??\����� �������'�@SSӔ_��233QZZʵ�D�	:Ec�������`
�-[�뮻K�.��kdY�'�|�w�y���t���`0`�Ǒ$)CaP��W������.O'�tN;�4L9���Q���x������iz��'9�^�K/�W^y��Y�V�����?�1�f/�I�� 4Ȳ�[�Ѵ;�NsSS��Pb���ջw�P�T�!��@�$IKdM����j�y��ַ�����)�<Y��i�&<��i�DO�$��;����&b���*++q�M7��SO��k��݋���/x�w`�X�}�� � �j������^q�{�}��_Ͱ��K�t�$IG��o ��I�T*���/����g�1�����x�'���sI�41AOb'�p֬Y����)���O�q�F��������!Ŀ l�x<�j">]'�t�fdd�F��
!N�$� ��U*�/_�J?���v��ׯ�+����������B���;"J LЉ($��yOOO��/M���q�UWaժUS���z������M�6lP�O��wdY����v�ڵ�P��Z�h�Q�V/B|�� VP��k4q�Yg�.�G1��߽{7x�.;�&�I(777�p�?�����e��>6l؀���h�z�&�x��t�����3���/�P�gϞ�$}�� �)�3�L8���q�%�L�2e]]������p��E�$����7�Di�	:����l���w(	g�ҥ���1w�܃��+����^zi�ٛu 6ɲ�?�v�UB~0,�1�~v��MD,[�t).��r����!�26oތ_���lM�$s�g���o?h��`0��������~����.!�+ �����o!D�?"=�c� ���% L����`ժU��w����Ig����㷿�-�}�ٴ:���QVV6�b D�:���7!�����ۋ���`��7ߌ/���ɡ�!<��3شi���	��$uȲ�{�F�ߵ��	_ i�������?�����BFGy$���Z�p�	}���n�y���Of!���=I�F�]�_���'�'���o������l6G��$i��)����޽{��lZ�h�N�V]qL�'//�_~9.���D����ڵk�=�H+���0�LP�T���b�	:Q��x<0�͊	e�;ꨣ������������3�<��^z	O�DԠ$I�˲�����w�aPL������_-I��P�պh�"�p�X�|���#�2�{�9<��S�nRc��-Z�Gy�k���uuuO	 �$�Ѻ���f+�xX�h��J�c c�z���*�t�M8�S&}�Ӊ{�o���,F�4L&rss�
�t����ׇ���x��p$I¥�^�n�a�ݑB��ׯ_������� ��D}}}�,�S^x�z߾}�B��+ϟ|�ɸ馛P]]=���ڵ��r�t�ا&�	��s��ڵk'-Da���裏����Ҵ�w����O�$��_�5G���$���qY+V��]w݅�����B��{�1n#n�F�n����Á��N��(����}�݇�O?}�~������{�o߾��F%Iz6>����7k�&�%K�+�� ��o��t�������{I�͆5k�`�֭�jRa����Z-n��v�w�y��{��w��C)m��J��e�Ν�Z�	���f�$I�@Q��ݦ�`�5�\�K/�tҊ��1n���ߎ8���������q'JqLЉ҃��CWW�������?�8��S�K�����������:F!��*��޺���Y6���Ԝ-I��q`˶��s����t�xY���O��g�e���0AO@YYY��/~��+WF��t:�裏bӦMO�!nkhh�8�A&�Ϟ��
����-��?<鴛��.\{�hkk��0��N�CII�A�Q�b�N��dY�����Rz@�sY�x1�x�	���G�k�.�]����O�)��͍���g3�Dv�I'i(I�= 
B�$��/ƍ7�8�h�o��{�~B�q�=����c����>����Oq��O,l&x泋�s��L�$�jjj�� ��צRp�j��n@mmm"M���())�F��w(D4Ø��.�˅��N�|�x����<�L���Q��NRج_�������!&�&�ŋ�x�UcۧRp>7��#)�X�&�	��ÆPRR�ϦM��nݺ��F!�e;f=�$�hѢj�J����D_����ӟ�4�������[oŖ-[bfRP��(**���2%&�D�'���v�=ޡ$�.� w�qG�]ll6n��6l۶m\���$����>�:�/>�� �U�333q���3Έ����\u�UJ�w���p�B<���(((P<�r�p��w㭷��.I��������&!I�TSS�} ���^�h~��_���L�u~���v�}��E�8�(�0A'JB����kzbժU��曣^���݋o�qb�q+�����)1&�e˖�|� �j�$	�W��7��.T[[����c` ���1AO Gy$6l�uk�����G?�޽{�6;\͋��,Y��hY�782�VTT�_���X�h��k�� ֮]�7�|3Va&�ш���I� !����(�	!�t:���������+����_���-[�f�������h4����O{�����l��6 ���<��c��#�D������_��u)AW�W��;�0��7����777��K/����$�+LΧo�Ν�dY��$I���q�e�EM��j5~��n����N'Z[[���?��)ň��Ekk+��ۙ�O��_<ir��?�	7�x����i�Nw*���B�����U*�J ��>� �V�Boo���*++��3��d2�(RR�v#���������W[[�k��N�j�I��Ǭ��l۶ͭ�"��1O�����T*~�ӟ��s�U|������_���h40�LQ6Q��:Qr
�������p�CI�>�뮨׼��>���&/������;�e˖����B��BmeeeذaC�����p�W��ȉ4��V	z^^^|�Ũ�;v���O��$����{͘c�9�<!�d ���r�-���K�{<\~��hll�e�I%##�����Ȉw(D4ELЉ��V�===��6�<~��_+�B��G��/�8�y�9�����U��N��ǘ*����~��*�����_~9<O�+&�q������b��Ŋ�mۆn�^�7�pe}}��1
1����|U������t�M�������b���K.�:%�<���Ɂ�d�lDI�	:QrB��M�~�ӳh�"<��s0�x���ꫯ�mnW�է���6�,�4��L�� �j����3�<5I��7q�m��E��DJ��b�$IX�n]��|ǎ��<69�K�t�����аM�R �q��W��+�����d2a����`>	!l6ZZZ`�X�t����s�z�hkkCkk+��i*++ï�k�� y䑉�y�$I'39���K�K���  `�Z�� ��튯9��3q�u��0J�$A��+p�i�)�khh�u�]7v��_������6�,�4�s��]B�S�Y�.��C=�7�xC�����q���s�� �BKK�����'�L
��������.}�)���x��GQTT�x��'��8�}�,�_���k�I�i����!��㡡!|���GO�r���(�)��/_�?�я�uww��믟����uuu�"͸���=�$�` dY��w��(ܩ��u<�a�X���
���p����,����Ǟ={Ҫ@�L[�v-�>�h�s�7o��O?=��Y�ќ��ؘ~{{�ICC� �����k���n��+I��~̛7/�!���N�KJJ��#�(���l������p�$I7��ս�	���kp p��-�܂�&�N7�p�-[�����Gww7���'n]BDDD8��c�޽�w8I��sύ�;�֭[q����m2n�����	!�
���⦛nR\ʑ���_��,F#)���T*<�����ˋ8q��7�[o!�XWWW�xC�1���?B|�8���u�]���Z�Raݺu��ɉu�I��񠣣���\GGDD����v;��ۇ��n��x����̙��n�M�\kk+n�喱�v _۽{wG�����1t��Gaݺu�}�Ν�[n�%V����M�W�^�/�ˊ��q|��G�cI�����x�bg������:t��Ӄ[o�U��Yii)����BZZZ����D�������(��ߏ���x����j5֭[�8��r�p��7�]V�p^}}}C,c���,˗x;���k�a��͊�/���G���L�,Xu��;＃^��,vI��\�}�C}}���<t����'�T�{ꩧ⬳ΊUh)�n����}}}�1!"���v���Ԅ��V�|�x��2���*���(����;���>�$����wcE����s��!�kKz�!�޽[���wމ����ŗ�R.AW�T�뮻��j#�������[�z@�V_�e�f'	���a-�<�{����*�]�f


bZ�B�j����K�,Annn�C"""�����hnn�{̀�?W\q�⹍7��w�����꞉I`4%MMMvI���l/x뭷*�`�������'�1��\����~K�,�h�ew�ql6[�Iq	�R$!�,Iҥ �����SZ������o�9�!�!,X�'�x���w��<��׋��v455q˴Y�R�p��B��E�3��x��G�6�p8��,8�����I��7՝��x�G��}��8�b[�I����$���?���֝X����NL�i����$�b A �<����_�:�/_��R��`�7��M<�����X������~�?��9��=^x���X0�O~��\�PӨJ��n[[�/$����� �����͛��{�)�]�v-�z}�BK+)���x㍊	��l�����6�����ޘF�����}!D����o��"�f����Ŗ�F#.��<���8��y&"����z��ى�{�r/�Y����k��F��/�0n�$I?޹s��X�F����]`_���T��������bY�H�}�������E�!p��������l�$}��Γ���@���>��|޼y8���cZZ�����ի��SO�.��w""JHB�|>��f�߿�F�E�\s���f����o�6���Γ�޽{�$��g�X-\y'�+��eee�/-�L�~뭷B����7�xc\�1!Ě����X�F����ɫR��Ę��SO=����k���h�exi#;;\p�z�)�Q'"����za6��o�>&�14g�\xᅊ�|����c�j�Zy*%������m�6mڄ����~z��^{mLcK)����8�c"�].��'>�766>��hF�ܹ�# �ǰ/��2���#�����K.�ehi'##���7��SO�{����Ss""�X�x<hkk���������k��h"ڷlق�۷���kkkk�c� !ĝ�$u|�=z�!Ȳ��k_��Ν��RY�'�$�ꫯV<��3��b���B�	!"?Y���n� �EG~��+�[�j�
;D�v�}J_~��{,֭[��.���:ńhmmESS�Ng�CJK����g�����'Vm�mll\ё^cc�@����ݻ��-��J����ѡ�jjj���%��O>�=�XD��b�Yg��^#��MCC�rJ
�/�
��B�6lP�����O��'��h��#I���PPP �V�p���F�Q\�ED��̙��/����8�S�NZ��/��N;-����^�C=4�����w#:R�X�x�; N���2���[�ɲ���;---�qF�t:ݎ;��H���.�L�}Æc׾صZ��1�főG�,���P�?좋.Bfff��"�Akk+�����p""�������s�[���Ϗw8i���B����ų�>;��u&��O��[� ��ۋ�^{-��J���իcZ�J�}��Ŋk�{{{�y���$I����O-)�lܸ1(Iҝ��;w�>�藓��o}�[1��B��t����zHDD�D�Vc�ʕ��o�{��e{��w�G��j�*�T�)�ƍ100:��˸hv466��)t��3ό;��a2�bZ�J�}ժU�������B�V!��� �t����
�����]r�%��<(v�n7�������ժXX���h,�N��}�kذa���j`ӦM��[p�	'����v�t4�����~<����c!����������T*�] ��e���_"�h�Z|�;߉uh))i3���"�|���v����6=Z__?��h�I�t����Z�m*++�r�ʘ�Eʼ^/�����ڊ��A&�DD�h4�K.�����V�;�'�x"�9��w�}x���Z��7�����������c3�B��#:Q�ڹs�~ �����y�����??b}:M_�&��s������*\.W�Х��~щ�Z}}�� �:~���{
�� `pp��ͰX,����QYY��կ";;=������r����h���;O���_{�?����;R�B<@ @ww7�{ｈ>yyy8��cY�I�]�$��5�,��W�w �x~ǎ����f�B /[x��������O�Z�$�2�����ڊ��N�S'"JCZ�===x������	yX�t)�͛���'�`߾}�c!įb�FCCC=�-��_~Y��>��LЗ-[�������۷���'t($Iz"��Q���?
!�	�_��׈>j�g�}v�c��B`tt]]]hmm���0���(!� z{{��؈O?�CCC�������b�������E<{�$��>��c���>+V�@IIIL�J5I���q���6m{�~}}�ޘD1�m�6�$I��T�7oVL�N?����E����a`` ---�����w"�!����FGG��ك��A�G�D��(n��p8���vR{:fAQ��@7p�����_ l�����'�t�J�SO=5��f������B��ޔ2$I
o���ۋ;vD�9��QYYӸ���A���������c�IQ�e###طo����p8�}˗/G^^^D��o�	��:� ��X�E��e˖�����o��8@m0��&��e˖��� �����'�@�Б���ZD'J)uuu�����o��G�$>�KR�f�---B0�wHDD4	!|>z{{�{�ntuuqFT��v/��[o�=�3wNJ}c��ܹ3�OMM���bVJI���NPl�p�x}۶m�Dq%������VL�;�B�    IDAT�D3����b��������wHDD4�,˰��hjj¾}�8�=�H��c�=6�}ppp��EI����QJilll�I���7ߌ�#I�?��}�����v�}�Q�X��W#:Q�z��HV��|�	���/��d��FVO �������\�*.��j��j!I�EGDDS%������� �������#�<RqW�-[�������S)Um�E��,�k�F܏�\�7nTz-DR%����;wnD����ǎ����>:/^�	�e �u�ֈ]�VcŊ��P�^�W^y匽_ ���w�}����A$"�e�,��t���^�7��P(�����?�����<�)�Ȳ�Y�R� ,��ߏ#�8b\�+V@������%�d�T	��+۷n��^�/i��,A���p�7Ft`�>}?��O0�|�s�v���?�x.�4���+_�
ZZZp�M7A�VC�I�KQ�s���������˗G����q�W��eL_���͋/n08p�=1A�����G����x��Ԓ�.��c�Ql���T��*J�,��R�����fX,���XK�,�Kl�j����K��l6�{�1����͛����k֬��`@nn.rrr�R%]�"���[n��a�XX�-M��j���D���֎�iE�T*�^M?� p l۶W\qED��K�2A?Iu�t�҈���NX,��J��0i�1�L�n(>��ӈ>��χ�h�uhII�$�z�Q��~�����aDSw�g⨣����F__���XX��hdY���@[[��݋��&�i��#�DFFFD��{��uuu1��$I���W�N(�ntpI�����aΜ9�J����6�,(J[�l	 �:V��A�Ra��ű+i�x�X�p���_}⚳�"I~�����p8���DKK,�BM ����Fgg'v�ލ��v>�$ �z�TWW�^��Ľ1�Y�����bϞ=}�9��=I��/\�P�����(]�t�t 8ꨣbL2���ۭV+y�G3}�w���<�ߏ��!����l6�j�rou"Jk^�سg���a�Z���ƙ��80�b�����N����+Me���Ciii,�J	I�]� �w�{�aL��D�-�Mss3�~?�Z�,�yP�f���Q��?��Ӱ���s].���_g0���Ƶ�T*\t�E���~6��s�\���CFF׫Q��������":(��ﮮ�q[תT���eL�P�8
 ��ݫ�a�����eLI/it��J�e�����U*U��fJ:�ng�F������#�9�;�s������+���Ͻ�����{�M�u'�|2{챈���:���/�4B�v��v���ߏ��,dgg#;;��:������e>4-*�
��͋h߿��������X�D�EQ��<�s�p�B�����eXI/i�@��?������|��X�D�cǎ� �B�J��;�I�A�|�Ɋ�/��rB	ڲe���#��������N����hjjBWWl6�{QR
Ass3��݋��n&�4-0�MM��=5�, JD�ܫ��]�^Q)���%�zEEED[[[��áݻws�Dzk P
D|6  Z�%%%�f�G������a���q����x��q�=�D�;���m۶�M�}�N'�N'�����������b'D��Bۢ9�N���7�^�%K�`ŊX�d	


�������𵶳�{���G}��۷'�C�t�tO D�c1AOcz��q�֮�.~����D�QtI����zD�wuu��B�Dt��"�h�$�4 ���Q�S^^�=�h#�[�n��j�q4S��{��?�i��/}�K3���,�f��f�A�$dee�h4";;j�zF~ѡ%������z��i���L\t�EX�z5�����������_�2V�Z�Պ�7�^���q�-��p��ݓ�؎;/^l� ���L�g@R�����T����T��!SJ+�$u����c,^$����������8��Z���80�J����Y���с���C*pGDt(��z��������-9_�l������?�q��<���<\u�Ux�7p�'�N�tP�����������Fi��d2A���2���#�&�I�}�H��
?��6J^\\�`�MMM�b���_�g��㏱t��qm�$�#�����K����b��`O��XY����e^�V�###��E�V��s�=��	 ��믟�P ^x!֬Y����f����c�=�����3MUQQQD������H�X�e�S�c�#�I����¨�[)RR$�ў��=�S�DiC��i1<<��'///�!%�Ѩ� ����%MO{{�b��f5AB�����h�Zdee��X����CY��r�022��Y�?�{.[��s�⹙�)u���;z�$��o���ß���yO�������q�Su:]dFFiE���>���X���LЧ!�t���^��Y�*�J5������r����9��t�٥���B��i�h�%���ձ�3~�V�V��$!333������>�N�����x<3���w�b����k��6#?���>��Ӽ��[�{�n�����{�2�{�	5i����+��Pڐ$)<b�fȦ')���\�����JOZ�vh�2V�5"A��YJw%%%�흝�1���D�9�K����hxt=T>33�U��X0����j��n�ܣ�9�����|�ͨ�^ӡ�h�����ZS�J�x �s����{�		�m�ƍ�_oA)E��� ���	z�����h�{Y���Svv�u����Gi?O�^�!Y�#����+��~?FFF022�J�����;?�D�m�(���H̶B+//�:�h���<���q�a�����Gmm-��ك��a�t:����-���UUU�����?��33MN�w҄߷���v���A��1����HУM	�G�$I�U��bn˖-�ŋ�(>a����w|u�?��L:�B��nIh�� rT=�pr���w*'*��ʩ4��
(F��I)"�C��B�!=�������o���dwvv��|<|����y��f^�i�^�,**Jq��,oc6�QZZj7!QDD��*�I�l��׮]C@@�-�����z%�r�,�l6��� 999���/7~W-�&�~���*�
�O<Q�1�$�/���%K��%$$`����ׯ��ϙ0aV�XQ����9J��*�Z��q�l�l6+���:�k�$I����7��0@�K�_����z�'L;{����=h�'��yyy���Ê+�cǎ������t�DT	Y��u[w��n��(�o߾�%���ׯ�9^L&�L���;wV�9�ϟǿ��/�5
3g�T���۶m�q�T9���
�V�i���,��ֿ�������9^Е��PXw�_�&��B���p\�ҳw�^�ݻץ�Yo S�~}ԯ_����,˸p�N�8���t���o^1�>�/�e���(,,Dnn.���4ٲ�(��*�>�������m�yY�|������3�(��߿?�
�p�mw3N�GE��~�Q:￝�]�]@@@�ׂ x���-�)�bq������xӘ谰0�m&��|			HHH�u����Fzz:�;���tdffz��,����!����|M���Nbb��6I�\2#z�F�ЩS'��w�ލ5k�8���|�	���������ٳ'A����U��;�� �;�$Y[�q��U��W�Z�� Qm�eY�����.����zʀ��QWv���
		Q���K]I�ڵѭ[7t����v�?�Ν�dk�7��E^RRbC^TT�u�0&&F�<##�%Ø�w�8t�jѢE��\I���[oa�ҥv����ШQ#dfr	nw�BOD��F.!�b��{�Q@����^�x�8:���'e��*}I�B����-��5��t4�����-Ξ=���t����������NT���($$$�]�vhР�qO�Tc�7Vܞ�����ر��}ǎ��y~���;wNq�֭[3��Y&��7��`�����9^���ժU˶OE�i��o���[d���﷨Vו+W�7j�H�J�'>>^q�իWU��u�^��p}wg�S�N2d����;w'N�����q��)N>G~G�e����A�HLLD�ΝѺu�rC����V�:�zFF�K>�C��mܸ�Ɵ�u�V<��v�[�n��۷����1�{�
�V\ܚ B����ҽ7��I�}�WtG�qԮ]���  Y��Yi��l.w(�(��Z�w�/_V�ޮ];�+�Guz�:�JM�T:�+V� p�g�6mЦM4m�+W�Dpp0BBBj�������,�E�ƍѲeK$%%�U�V^5�FM8ZF��6l��:���?�������;j��T�7n��^�poӧO��;vp��+����`�kT5^q��Htt��gQ�Ui�,˱֟������B����!˲ݒ6͛7Gdd���Cw4C�+Z��AII	JJJ��E�\hFXX��GDZ ˲mV����o���_вeK��A�Q�VNNN�?��w/p�g�+��O�<���уr�{���r��BNNNm \Rďɲ\�zoP���q���?��k�c�e�;˒��o�b��	� ���� 33Ӯ+�(��ի6l���n/88w�y��_�U�j|�$I(***7?� 		�����`1��j�A�b��d2���������ða�p��"..�F�8}���׉�SZ��K�V���СC5�|�fO���R�^=�2��7S���xe6��ݯ��X�z��(���s�"�;GZ�[�,��T*�����Gc��n�ciii�c��ޫW/����m�X,HOO�@E�K�eۍ%AAA�B�5�3�Su�m/))��dBAA
mEDD�O�>6l���]o���شi֯_��Ǵ"$Dy/Wc��t����,�((((�kp�3�\G�)44��SQ�8�ri�!�,Wz�-�2�_��jM��+��q�e/A��Si�,�M�?;�4�3�:���?cРAv���n���k��nܸq��SSS9)�J�kCW���ܭ��e[���N@�^ZZ
���Ʉ��B+.(�"�v�aÆ���5K.IRSS�~�z|��wW��f����l:C�m���~W> U
�lAw?G�����.IR3K"m�t����ׯs�f'yE@/**Bvv�]��
AU�"-J���]�!Sv�؁3fحg+�"&N��Y�fy�2�:t�Ν;+�۱c���PE����5����m��!�b��$�b��l6�za���T1�+i֬��Ç�x��+W���CJJ���U�h�����Y͚5Cdd��>Y���o�����*-��������5�3���ۖ�!Q� �:�.VE[�v��f�{;�+:p�nŀ^a�8�N� --My:j���v͚5��YZZ�p91���O8p ]�t��7r�H��������LY@@ ^x��}�$a�֭*WD�2��0��(,,��'h�� ș�5@�$�x���R��f[w���b[˸u|��\م���?��֯_�]�vA��j�7���U�޼ys��Ue0�p�K'UG_PP��'e��U�k��L���DQ���DBB��1��󚻛����N			�u�� ���� l��Z�nmw̙3g��R㯾��Kŀ.�"�͛�x@3kf?��S�W�ڵ���\�nώ�*X��[��ҿ��L�+�%I��z[[�KJJl���?+�l֔(�0�6l��p���:~����?NT�(��jժF�����p���ѪC�۵�ȗ]�p&��n���r�掟Ԑϓe�`}pڼys�����vY^�k��S�춉��-Zغ����5�"m�$)���-00P�]���oߎ�/*vQjҤ	�ϟ���~�a�e�>&Lp�����Cc�B_���� ��X�g�kG��5�ڥ���֠mm�.��f�-|[�y�e�aÆ<x0ƌ�p�����Ŗ-[�j�*��,��2e;v,���AгgO��8��g:�8���I�������+<܉���	ǎ;�jq�	� �Z�+<������&�;�ӦM����j���������5o�q{�$����k�����G�X�`��y�u/5jf̘ᰫ�����o�>��"�+�"_�(�K�.8p z��e{8`6�QTTI�PPP`��e�*�������ѣG���&ϱ��-��m��\�;y����ۛ���஻���ѣk܅]�$�߿)))رc�m�ww��%dee�N�:嶇���W�^ز��v���ۣ^�z��2�+=p�*�ZN�:e�Q�!I7 ������6m�(��o�yM@?q�dY��坔���� � �璯�f�!))I�'N�V�7���o��@�WV֫W/,_�S�NU�e*<<S�L��Q�#I�ϟ�ZM���7o�A��db2k���_��	��M�.�C���rYgΜ�ƍ�v�Z\�t�EU����4�u�]v�'L������9F��pߕ+Wp��9�kt��X�?���e� ����1|��r�DQ�^��O?� ��U(�<���R�XC�����\~/W�����l�?M�4)����P_�׷8v�;���c��L@�С��1�,��Q.�Y�,㥗^�ʕ+��{�w`�ʕ���/�d�dee����� <�<�L�-6 �l�2>��s��d�V����c˖-~��L�0d��5Jq"!g�L&�ܹ)))��矫=	��8x�b@��t���{�~��*V\\��puZ�+c4��9sƥ�!e��HJJ�t l �C�,wA���`�� p��~?W��t 8|��]@OHH@�:ulA�� ��ȉ':�M��/##999j���N�>��s�b�̙�	����1z�h|��wX�~=>�.�ΎGMMM�{��s���va6l���W��Ξ=�6`ݺu�����ܜ�-%%6lP����m޼�'OV��1cΟ?�#G���sDQČ3*]{��o��Q�9
�lAWGzz:������W�$���h����zU�����[��t��U�{��y]@���Ft�޽���� >T�6�I�Zo:Z�h��s��!���z)))hٲ%ƍW�q!!!9r$F���ׯ�_~��C�p�ԩ*?	

BӦMѲeKt��	�Z���:�����׿��Y��iM�6Ő!C\҅�����]�v=z4����}ֵkװ~�z�^�ڥ]��ɥK���?*�����b���x뭷����𺍌�Č3p��w;<OFF�K�o4o�qqqv�q��Y���+--űc�йs�rۓ��j]eC��J�H"� ��=z�P<���ê��K�*����ϊ�{��Y6����t�iii��f�T#�`�ώf�ݿ�j���y��!22Æ���u������1x��	���q��u����d2�d2AEDDD $$u��ALLL�k��������p� ����8Çw8gEUɲ�#G�`͚5زe�_��6l�Ç�}�݇ƍ�賬k��Y�?����M~�EK�.E�޽[����1c�<��Cظq#�?���,�����8t��C�Ett�m��J��{���#G��e�?R��~���.]��� Ȳ<�~�h46`[�X)��رcj��3�*�gff�̙3v3zv���(Z�G
���w(�Tf4�-ܭ�a�X8�w5I���ӧ�x�'�����5�Yw�ܹs�4i[��)��t�FU\�v[�l��ի9C�-�'OƠA�n`%222�~�z�Y����.�����vӦM��VԬY�j�gdd`Æ�-ώ(�:t�⾃��<t{�w�ƓO>i��W�^��`XbbbȩS��w�?"I�H�þ:u�(���~�/�뭼*���={�zLL:w�\��},���,�c ���S�Nv�=z���j��3dY��ŋq��L�:�ұ�jڱc�O����<O�B~�l6c�޽X�~=�m��!.����͛7�� ��={6:t���(�    IDAT���seY����]�ӡcǎ���r7���~�Mq���}�b������ѡ�����o� ��֟���8$q��ݪ��K�6�SC�<�+g�����A����<�4�������?sڵk����իWc�����#//3f���O?�pN�����ѿ���Ė-[�kH�$�۷/��"���Y�f1���ƍ�<y�ˇb,]�{��u�g��/Qܞ�����4���*'I���c��nݺ�&�E�~�������nk0`��1�,3�׀������ƍv���뇀� �����P�ov�F��5�;��u�t��/��ܹsx�G0e��'�1��HII��aðn�:U�M�'??)))x�G0b�,[�������z�/_Ʋe�0t�P<���X�~�u�)RIZZ�|�I��,ۺu+�}�]�|�U�ƍ.���?�l6��|t{����{ɲ<:99���ʐ�x�z�֭[W��꯿����L���^���b�`�֭=zt��111�ի~�� � ��J�
I-�$Mn��_�>�t�bw����9>��dYƖ-[�m�6�}��3f�v�Z�ם�������]�֭���+W�`�vۯ^�8eI����T�_��~�-���pv{�9x� Ə�ٳgC��U�3dY�ҥK���|�����e]�ٺu�K�EU�w�^����M8p�@̟?�:�8�b��WS�Y� ��a�����ޫx��i�&5��9^Ё��yV� 0j�([@p�N�k���vZ��H���!aaa[_�1B�b��ͪ��O,�mۆm۶!..�z�BϞ=���l7N�&�	���ػw/v�څ�Ǐs��v��-[��24�ʕ+����.x��q��q�Î�,�H�:{�,z�!�w�}�8q"�4iR���ٳ���[��7j���w�⾢�"v�����Rl߾#F�(�=&&��sO�@�8�}�^�(�rS���p������j]��+�/����/�MҫW/4h� �/_ !  �� ��D��^�����n���4VM�$lܸQ���ҵkװz�j�^� P�^=�i��7F�z�P�^=#**�����b�L&dee��ի�|�2222p��i��%�c��{\�~�7oƚ5kp��IO�C�a�X�f��]�F�ݺu��`@BBbbb���<dgg#33����޽{q����ԵkW�������g������٨Q���F��Wjj*' �M�X�С�7onw����q��%U��5^�%I�ڵk1iҤr�EQ��ѣmc�dY�ضm�Y������A���ܻwoř^w��e}XC*�z�*�O�f�޽�6mB~~��K�)�/ƹs����ɲ�#G�x|P ����:tHq��.]��E����  Ȳ< ��1z ���x�������n�8�5k�(v{����f}�������� ��������)�|�2ù����D>L�e�{+A��C��t_RRR+�
#UȲ<�&�kԨ���owLNN�o߮vi>�k��+Wʎ7����.7vI�g۴i�bi�~/Y�������t��%������yk׮��d��>t�в��Ȳ<]��ȭ���Ag}��C)N���� �xm@��>�Lq��	ʮ�]'$$�)����!(���c�=�x����ْCDDD�B7n�P\�4$$?l���,�3mԬ���b���[C��ԩ��#G�SZZ��˗�\�o��~��!=z�n{|||�I,dY����bլ�\O���۵k�������|vo'"""r��>�Lq��<P��,5�"��5��~��'�Nl�q�F���"^���O?U���c�!$$��2Fŗժ��C��M �������'n-�^�W_}��DDDDnp��9�ر�n{XX&N�Xv����K���儛7�o�����a̘1v�ɲ�g39���֭[q��	��4��q��nzB�ӵS�0r)�N!«��]�tA�=�+,,��-Z���d�M�4���e��[= ��� �m}����l���<F���adY��ŋ�=��㈋���E�A�ɕ4O�W 4��3^x���>��sdgg�Y�_9u��m�f�=((�'O.���^�W�0�4-999F��y��mڴ����펓$	|�����:�� �c����v������O��t�N�S^��4K���&�3f����e�9�
�����]�t)�i^RRR�j��K�����>ps)�iӦA��ƍq��I���i>�eY�ܹs!˲ݾ���/����N�@����:u�$��2ܚ9�nݺ��?��x��ŋ����fyDDDD~)##)))��f̘Q�+t�,�o�V՘�`�(��X_W�SV&�	�󎪵��� p��l޼�n�(�x�W�~I�X1v�X���HsJJJf���pӦMCTT��q���;���+5K#"""�k��nܸa��iӦ�ey��h|D�ڨz�Fc8��qkb������l�-[��/�X�� .Dqq���f͚U���s�ĉ�j�F�����L���ӧ���x����QZZ�ViDDDD~/''~���G}�[����e�]�N�R�ڨz$IZ�����/������._��O>�D����O�/:�0n�ĉ0��ײ,�b0z�U9G���
��������bƌ��nڴ	{��Q�<""""�b�
?~�n{`` �̙S�k�(���t�`U�*����
������ދ�*;g��V�?� �}���D@@ �̙����& _q<��� ����f�^c֬Y�[��ݱ999�;w��ps�3g*�dlѢ�y晲������j�Q�%%%��6�<>>�����ݲe�o߮Zm�����b�+����%_���(�s}Fm���/l}����wo��o������*�����*8y�$>��S�}�ƍ�]w�Uv�?�z�C�FUb4�%IZ�ps���s�mش�����9s�.ѯ�d0�����7x�`�?��A��=U
�����c؞�$%%�駟V<v���X�n�Z���/Fzz��vA0g�4o޼�%:������2ADY�� �κ��矇�`P<���^�����*�/�d@��>��V���ϖ[*@���5��I5III=A��  ���Âhw�k����/�\!))))��i�`2�������7�@XX�uS�(�_'%%�R�H�c0 �����a�p���+�n�:lڴI�����tI�0m�4�u��`�4nܸ��Y��q�
�r�^��u B �V�Zx�wP�N�c%I/����yFFF�ϟ��/11s�́(��GI�6t�С�jR9��yY����NNN�̙3�=w�����g:psV���ߐ$�n_ll,>��Ԯ]���EF�q�j �֒��7׮�={6ڶm�x��E��o�>+$"""��X�j��!�}����)S�njQZZ�C���W�8������%�ƍc��egݷ1�L�2e



�,�o�t@��;w:\�1!!,@hh�uS�,˟�~�����(n��9N��_D�>�Òv�܉%K��Y"9��^É'�=���x���nj%�m��w�$�0�#�VZ�n]�������U<���^R�_����: ����عs��:`��-�
�;�^?B�����`h`'�&�m�'OƘ1c�?s��DDDD�����׿��p8��>�ѣ�uZ������O���/�%��������I�&�����ذa������eO��Z�j��?v�mz���2eJ���̂ <�����jE�����F q�mO<��x�	�㳳�1~�x\�pA�
��aÆ9r��� ""y���a�X<]�Mrr2>��C�nӒ$a������om�dY>e�X�?~���u����oY�_�������~�N�x��;0y�d�h>p����u ~� .._|�6l����ĳ�>[v�IY�Y���/�U�?HJJxk��(�G}�<���&�	�=��9�V��סC|��'�.���4�s�Ί3hyҀ0o޼����H��Y�fa���e7_�$龴��_T+�Ǎ;6��~{[�I�mQQQX�x1�z��{�?����o(**R�NO�R@��.�V׮]äI�������w��x�w�.!Ȳ���`�@��+�����럒$�;�
� `�ԩ�yii)�{�9�s""""/�e��3�����^z	�Ǐ/���(�?p��k$''Ǥ��[6������O?u�Ϝ9�I�&�M8��
�����q���(��ڵ+�.]Zqy��EQܫ��[�R�j޼y��h\"� @pp0^�u�7N�=���~��+%""""WZ�|9�}�]�}� ��^�/�P���� ��9cǎP�Pc0:Z,� Y�5i��1Z�P�5�/_�������?�T�L���: �8q���?.���|��nGA��Q��Ct:]����}�,O�n����G}��C�*����i�ƍ��IDDDD���V�����1gΜ��� /���o�СC��7�A���4�� l��K�.X�b��	�\���'��ŋ*UJJ�2�@jj*{�1�-�5�g�}����Y�S�F�gݻwS|#�c4E�0 �u[�V���_ 99Y�=�3f̨8��������o��E�9�?h� ,]����+�y@iii��h��}@bbb�^��J�� lCt��~,^�QQQ�����Ą	p��y�J%�6�@ZZ&L��k׮)���o��g�y����,?�����`0(� �����a�,˟��n<x0>��s�O��f3��y�_�^�R����H%��>^�uȲ�<��)))���;�n�'��:�^�^�6m"U)���{���R��,		��/��_|AAA����?0a�dff�U*U¯fqw�I�&X�h��� ?���O�^1̗x3//��?�����uzA���,�o��Ŕ)S0v�X�������ɓ���?�Q�W��,��|�𗪷z��ѫW/O���l6�7���3g<]�K5l�S�NEhh��KQt��,Y����Gyݻw�t�L&�ϟ�s�7�7���?��̔�Ug���ಓ�����B�͚���>|8^z�%*�X,X�h�.]Zq���� <�����*�z������2�c�94  ТE̝;�Z�r��#G�੧�r�f����,��DGGc��ر��c�������6m*�]��S�(>�����;z���� �,��E��7o���ի��?����tw��<�SSS1m�4���SEL�6����t)��f����ػw��Kq�^�9s�V�Z�.�����cƌ())�t).��3gj�d����q��O���s��q{v6�#""� ��`/#�2���}��/�ҥ,X��HǍ�G�ŴiӔޭ�e��cǎe��HA����
�ܸ�aÆa���~�lݺӦM��`@�,kG�Y�_����Wz���,�S�;v�mEj��hl,I�k� <�2�&���1q�D���wإ���;y�d�C�^U��c�*>u����t,]�ԧ[#A��q�йsgO�����1~��WO��V͚5�O<�J�bU?~���_�=�:t���R �|��G��ɓ�.ŭZ�h��{�Z�F"""θ\�3=88��P�ҽC�-�����Ҟ����X�p!����=�JAx[��>�WM�F��Y�� PnR���x̘1���R�,c�ҥx��w]r���5n���x��gv����l̝;6l��K�;��2=---խ�z��h�'�� <�����d̜9�7�V��ܹs}�f�������x!22�'[X����{�I� �������/)--E^^��o|�5Q	�u���f���9=t�S�NX�l�m��j@��p^��u�\dd$^����3�9t�f͚�����< � �=z�h��������, ����ēO>Y����|L�>۷ows�ޅ�$''c޼y�_�~��<xs��U�-ɲ�F�7RSS���PHJJj%��dY�' (�P�~}<��32dH�7�EEEx��W9\5���-� 7�*x�f�����C��+O���f3����]�CBBQ�1��!]�A�c�=�'�x��>/--�ʕ+����#//���� ,x�СC>�V� �^�,�Y��T�߽{w<��s�m;y�$�}�Y�={�m�z+t/��^z��R%I�ڵk���ҥKv�A�#��⼼�o�u2��c��8q��$I�A�
+ DDD��Ƅ	n�}��_�ԩS��Pjt�e��Xݿ��X�,rssU��έ<\A@TTT�=�|���\�y�3�{�ш9s� >>��㲳������o�Q�P"�W�$���1��ȥS�N�f�y�,�Oh_qbb"�z���<�e+V���w�t/3r�HL�2�O�KJJ��7�`ɒ%��S�)� V=zt����6 �x@B���j�¸q���#� ::��ϲX,��O��{��=�	wt���R3��{8�*--Enn�j���kkbYj���pn�LHwE@�~C�w����ԩSq�}����K�.��?ĺu��_�&�ǒ$}y��1�/1v�؀���> �����fRm޼9�x�	0��R�J�]���3gbϞ=�)�G0�{����*��l6��i�&,[�'�<`� ������c�M$VA����EQ��h �k���������_��W�����sO�<��_~iii.��?�3��&����B��\��R�Z-�|U��x��W�k��=44�j���Q1�{�=z`ƌhԨ�m��~�:���k,_����J�� �HE��#G�hff��ݻ��%I�}� �B�٭ڶm�|C��t p����~�y��!''�e�t/6p�@<��s�WO��M9�,c���X�jv��U�/�Y��
���$I�۵kwlժU�^	���Z��n� �#��  ��5
C��Ҭ��������bQ�?��+�3�(sgpa`Q������׺���k�&=$$����+`H��j�O>�����U������ڵk��7�T�P �����eOZZ�9W�|;:�.X�N ����]�0�UHH���1c� 99Y�;�O�ƫ���C���hǀ�����0q�D<��#U^��իX�n6l�p�/��L�pL��DQ����×j�-�C�q%%%��I��^�,˝A�[���ի��b�ȑUZ��9.���x��|��#�3�W�-�,�sWHg`��u���Z�n@Exx����5��k���y��x���ѣG�*�����X�n�m�V�V�L dY��QY�O����m}��	�r�J�(�w������?I�0�rY� @��c�С:t(����t�7n`ѢE����0�$tѨQ#<��:t�m��u��il޼;w�ĉ'�kip�5A�dY�`�e9G�ouY�#EQ�e9@�[�4P��ҍ7F�޽1`� $%%9����O?�w�awv7ru@gkbո2�0�T��C:�yո2��������v��w�]��	��T5�ާgϞxꩧЦM�*��l6c߾}����k�.dee9s��y��%�r� Y�yO^X�  � �ɲ\@AȲ��־�EF�}�����ԭ��d2��/�Ē%K؝���}L�f�0iҤ*M�Pѵkװg��߿�Fff����\ll,�F#�t�=z�Y�fN�����������/��qe@g`qNQQ
o`%X�#Irrrj�ٚ�W<���G!�ـ�Z���"ҽ� �۷/&M���-[:�^Y�����={�����HMME~~��*uL�q�HJJB�n�еk�*��[��� %%K�.e��b@�Q͚5��?�aÆU��{E׮]Cjj*N�<�ӧO�ĉ�x�˺���z��E�hݺ5���ȁ�7�?��>��S>|�%5��*���zj�X���-���S��.�""##�K�IJ׺3]^�ՠƄ��z�(�w��x�Gбc�j}�$I8u�~��W�:u
�N���ӧ��{q�  PIDAT�����`$$$ 11�Z�B�V�`4o��#���X�jV�\�`�"�>.66cǎň#аa���b��+Wp��\�r999�q�nܸ���R��~aaa

BTTbbbP�vmԭ[���hԨ���k\S^^���[�X���{�+:K�T'�3�׌�bA^^��,ٚX3���W��HUz�=\�;�_1�{7�N�q�ơ���n(+���������DVV���q��۲�'�[���Att4j׮��">>qqq.i�����_��k�ָ7�ǀ�'DQD���1r�H�����iJ��C�a͚5زeg?���t�(..FAAA��ek�k8�y���3!=   ����5T�%�*}�ʕ���U��w1�{���H�{�1b�S�Ե*??��=V�^���TO�㳴�y��F�$a���ؽ{7"""ЧO4]�vEPP���8Y�q��Ql޼[�l�իW=]��넆�B����&�N@@ ����4&�׺넅�\��v�:ù�X�����������>S�*�g���I���+Wb�ʕhڴ)��:=Vݓ����s�Nl޼�w�f���a������;�DϞ=ѽ{w�fiTÍ7�o�>�޽{��qv�KRAu[�X��d29�`���=$IB^^JKK��Zw��Z�EQDtt�ӓ�R�$IB�&M���+�_�l��}T}����%>>=z�@�^�йsg��������={�g�:t��\elA�sؾ};�o���rm���HJJ��`�w�ᒱ3U!IΞ=���49r�������o�%X�'$$�,�uwg8w됁��\���jղ���k9jIg8wQq��%�={M�6-�oɒ%X�|��*�mU�5B�#33�V�ªU��6m� ))	���h׮���U�4����N�Bjj*>�#G��A�l؂�Ahڴ)ѴiS4j��7F�P�N�'�2�L���ƥK�p��\�x�ϟ��ӧ����'t^��t�su�mIg`Q�$I�B:ù:�ο`��kݽj׮���z͚5�,�x����7�x�,�ǖt���-[�e˖hܸ1���� ::�鹤���p��5\�t	����x�"Μ9��'O"33��a��tt/����r_�u

`�X I�m�w���{�	� 0��������,*�e���		Ahh�������W�vm������z�jO��7�	���߂  ((aaa�$��p�d2��]�D2�CK�]ܽPII	�]��u�DQd`QYhh(���XT$"""8�@e��՗���Y�fqyS�����l6�l�Ľ;yHAA


p��EO�B>��U�|�Zc��<�׺g��]}�DD���������HЉ������4��������HЉ������4��������HЉ������4��������HЉ������4��������HЉ������4��������HЉ������4��������HЉ������4��������HЉ������4��������H=] ����h����v>�Ʉ��,�ΧE�(�aÆ����ի0�ͪ�Skj׮���0��WTT���l�ΧEAAA���S��W�\��bQ��Z���P���k���	:�Ո#мys��w��e,^�X��iQll,�qUϹl�2�={V�sj͈#дiS��w��|��G��O�4h����爵�>T=�֌=�����ٳX�l�j�#"�$vq'""""""� t"""""""`@'""""""� t"""""""`@'""""""� t"""""""`@'""""""� t"""""""`@'""""""� t"""""""`@'""""""Ҁ@O@D����&�I��y.��$I�?I�T=��L&^�*�X,��=���H�?���b��ED�i�D�VǎC~~�j�~��j�Ҫ��<=zT�s޸qC��i�ѣG������.^��ڹ�*''G�k=//O��i�ѣG������Ο?�ڹ��<�]܉������4��������HЉ������4��������HЉ������4��������HЉ������4��������HЉ������4��������HЉ������4��������HЉ������4��������HЉ������4��������HЉ������4��������HЉ|�$I�$��e�Y�QZZ��2���l浮2Y�a6�=]��1�����t~E�$X,O�AD~��ȇɲ����Ȳ���\��磨������Ʉ��|����ZW�$I���ᵮ����=������N�:�.�/H���"R:����H��½����z^XX�ࢂ��b��� ,o�U`,����B{�*�7f�<��3M�6�[o�Ő�f�$!//���D�*t"?P�\���b����Bz�*�W\\����r�,H����>�r���hL�4	� ض5i�,@ݺu=X��^��DDjc@'���E�t׺�Ï��"�t7(**��V| ��Q��\�k�=�����/!!,@\\��U�6��$"Ob@'�#lp��vdHw������yZ,vMu��`�ת�wG�ƍ���o�aÆ*U����AD�ƀN�g8��5�}�������W�V0�p6��Zwg�4h��rhG��i:��MH�T7��&4#�U'���H�T��)d�:=�ի���"~�W� "�`@'�S�&6��մ���dbp����ʲ�H��t��E {5�_q5	�� ADZN��x3�W�<�.&˲�*�m���^#�qUk"[ҝ����@�9�D�5�D~�!�j\���d2����!�6\938{�T���u9<^�+((p�z�| U5����D�9�DĐ~�jaQZǛ��;���^9w_���\έ8�B�ΉH�Љ ��#���h2�������f�,V�֕����u�,�Q����k�!]Yii)���x-�&1���5���fO��	j�M,))���e�3�[1��g���݁�:�ݔ������s�Z/���rNDZ����}Z�hQ�����7t���AݺuU;gII�߷0֪U�k�V����=s��������*_����5:�5�GEE!0�o��f3���ΉH���[���X����5�Lx��q��AV���o **J�s�۷3g���^�(������U?wqq1������ê���Z�n����#22R�s���x�����(��:u*����y�=��[;yvq'"E!!!�={6�u���RTժU+���	� еkW��?�App�G��	�(�^�H8���P̞=:t���=E��᭷��H8����f�BPP�G��	���x饗T�V�:��:!�9yt"r(((�f�B���=]�*ڷo�x,�X�y�~�EQĴi�0`� ����_�:u�hj����;w.jժ��:�u�Y�f�ŵ��3g�w���C�e����MH7���D�UЉ�R���x�WгgOO��V:�����x`��ҥ�Ν���PO��6���x��ѯ_?O���B��?�2��V]�v���n��{����R �OH/))a8'"�ÀND�e햩��KW�Z`�JJJ�ܹs��R\N��TPP^y�����ӥ���hĜ9s4wM�y�x��W��R\N�ה5����x���NGD�m�^�ǊD^�C���OT?oii)�=�Tk��ӧq��7VU^ll,�S���t��ϟ�իW�|��lƞ={�X��.]�8���N�:h֬��
����R���:���'O��ŋn��^���Ѷm[�ޣ��5�R}��Y\�~���b���n��^�N�Q���֭��M�����ӹsg��m��I�v�;�é������}��9����R��Q�8p@݊�oO"����@�'����U5�GEE�cǎ��O			HHH���EEE�����#66V�s�S``���Qvv��=66����M�:f���O�z�v���9�I�e�����L�$I>���Ȋ]܉������4��������H8��yMw�m۪6� �����/��v>-


B߾}U=��ݻ�~B����;5��.]���8y_��D�{��A^^��笪+W��r�=z�e˖���9����v�ȿp:Ո�lV�F���� `2�����]<1�]VVnܸ��y��y�檞��������(�ϙ�����l��KDD��]܉������4��������HЉ������4��������HЉ������4��������HЉ������4��������H��tD�4h0	���W�v� ��u>-��������lذ��7n�S�ZӠA��ܫ�����������^�z	 ��y�F��Ovv��j�Sk4h0�@Ϸ�j�������K=]�U�ѣG�z�"�]o���j� jժ����k�gϮ��9�u���W_}����Ւ7�|s��狌�������y�Z�}Ύ;�[�r�Q�ϫ%o���85�q�߯u"���NDDDDDD��DDDDDDD��NDDDDDD��DDDDDDD��NDDDDDD��DDDDDDD��NDDDDDD��DDDDDDD��NDDDDDD��DDDDDDD��NDDDDDD��DDDDDDD��NDDDDDD��DDDDDDD��NDDDDDD��DDDDDDD��NDDDDDD��DDDDDDD��NDDDDDD��DDDDDDD��NDDDDDD��DDDDDDD��NDDDDDD��DDDDDDD��NDDDDDD��DDDDDDD��NDDDDDD��DDDDDDD��NDDDDDD��DDDDDDD��NDDDDDD��DDDDDDD��NDDDDDD��DDDDDDD��NDDDDDD��DDDDDDD��NDDDDDD��DDDDDDD��NDDDDDD��DDDDDDD��NDDDDDD��DDDDDDD��NDDDDDD��DDDDDDD��NDDDDDD��DDDDDDD��NDDDDDD��DDDDDDD��NDDDDDD��DDDDDDD��NDDDDDD��DDDDDDD��NDDDDDD��DDDDDDD��NDDDDDD��DDDDDDD��NDDDDDD��DDDDDDD��NDDDDDD��DDDDDDD��NDDDDDD��DDDDDDD��NDDDDDD��DDDDDDD��NDDDDDD��DDDDDDD��NDDDDDD��DDDDDDD��NDDDDDD��DDDDDDD��NDDDDDD��DDDDDDD��NDDDDDD��DDDDDDD��NDDDDDD��DDDDDDD��N��]�Im
�(*�I���*�h��o�[��#ۃ��>_�s6��7�t�   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  ��ե/ �����~}}=l�|>o��E���ݎ<�i����<O��g�h���ӯ�j�cuY��acQ������ǡ�߇=??������,��ac &Ё�j�^oG�@��Ƣ>??o___�n����>Z������a���tz6uss�m�硛��n����f�rww7l�x<���\�_�   @�  @�@  � �      � �@���9�    IEND�B`�PK
     `+�[/�i�$  �$  /   images/60da03ea-f7cc-456a-983c-41a209708cd9.png�PNG

   IHDR   d   �   ep�M   	pHYs  ��  ��"篻   tEXtSoftware www.inkscape.org��<  $IDATx��	����k�E@\@���%7P�\A@M\p	Ab��4&�hF�#���W@��\PO܎(�: ��!QqAEAt&����XS�]��gzp�9=Kwu�{�����{/s�A���9����aÆAIII�	ꩠ����ν��ʂ���`���r�z���<*--u�çL&�~��X@6n�4h� �s�=�=��#hҤI��W_��~����5`뭷~��|�M����-[�v�ygǳ�>�,x���U�V9��dÆA���N8!hڴ������1�V�͛7j��/�����/�̝;7�f�m�#1 ���{�~��o0�e|Zh }g<��$��ҥK��g�5k�xެ��x�~���;l���ӯ5j�S���o��VСCİ�e�]����O���ĉ]�~L;�c0h� 4Ʉ�����^z�]����g�����{饗���q��$�Rnֽ{�����w��g�|�UW�ߺuk�p��U�V�7n��/~�&L�l���g�}�G#)�) `?�0lذ�'Ov�
�n�|����}���t���s0�/�K��իc�W%@0H��[p�1Ǭ9r�YF���ш/�b ���_9bĈ��>s޼y;�\��Ga�� �h~??��OS��������8 ���σ���;�1c���^{��i��v͘1cb�I%@0�F���c��?��c�S��󟕾��;�8��@�{�����x��?���t��0|�1�z����7߬t��1M��"�e��W6�����r�  ��^{ӦM���ٳ�U�������1���v�:�Ǡ��H�i��S�LYмys�Urꉀo���_x�۶m; 5�G�S�̚5k9�v�m�b�
��
��>��7_�n]j߻.j[���_/\�`��*��׿r^h3��ڵk��i���sQ6/��FA���8BJ�:�(Uf �m�@�����H���^߁��*M�Q \h���a�0y�W�v7P�4n頠��̓�u�=�g�}�=�E�jH�o��uG�$��c���ْY��W_}���(�k�.<x�k�9��{�t;B:dٲe��h6�e�N���M�"�,/��>��#�/\���#����:uj0p���C���s��+`<�g%B2<�����G`��n<�����w_�򥰾��٤0��uMMK,�#-b��v]t��6BjL�����+ ��G}4X�hѯM��M
+q�������o~�s��m.�Z��� �Z�X�!��A#�D�Օ15�Ĥ��o������0�J�bhïhү� �A��_s�5o��:��S��g1�i�SO=���={����;sZU�4L}����o~ݤ�O?��@@�������?��}~�%K�4iRl�CŐ0�( �(�oܸ�{qOe���+���<Ës�:�,���|���`��
^x�����Ο?�=���٫W/ڿ��q�=�[�֐,GR�)���	�<�v_�lϴ̰�|b⺳��N�w\'\9T\\��l��vYPI3zٴiS�rн�Ң�Q���r��܇{�R����/@�M J+9��lgp�m�}����ѣG�3v��)v�wI.��he�x�ʕ��q��Z�|_V@��
�����w��#�������:��:|�g�o]�"I`����k�IX����i)
,��� ��&�B�50��i��Z��g��S����+�o�5�
sF�*lԥ�}#�+�(5�馛�>xf�����O�*5������́�q�|���� �aǃ��͂'rC7·q4�#���u���%�%p�Qt�f�0�|���/051�Ɇ'F������S�),5L5 դ�?��#��|f�0�q� ��k��e�]�8��*T0������@Z�Ӭ�A� ��G��A��p`��S��F�� �T0��^]%ڎ*#=D��Pc����	���g`d�DH`��'��V�4OТE��MD�8dS�T��~���b�nݺS�L	�8�'A�E���6l��EaiQz0j�(���ڀ�1̖���`D��2�+^	��Ț =�L�Gӵ���=$��:���-@h�/^�U�-"�H�b$� P�sJ{�?3<�x��`�<C�����H��&B�� v�9t�f~��e%5N><�,_0�����#d��P�b3I�rY"݋��	��V~+�����l�
k=S��`�w�� :���{�ed��f��hV����:�$#��L�� 8� ��￿��/\a�嫮�Ԁ*O�PZ�	D�t�B�)���	f6����� �Ѯ|�@PuްQG�}�T�HM��:
��D��vm�(jL�0D贉 0�*�ݒ8�'�n8�L�/o@�1 ��҂��`T�\D���]]#[]�a v��#� R��E��0�XL�U��K^��8a�M�6C��w'iG��(�5?��H�D�!1���C��+-\�w����
>)$@����[Bp�K�k��4=D#�z*�}T`b[P� D?|A�����W$Bq��M����f����S��x~�x�`,j�;� �J��X@T<���%�!]P��E�l�{ME适Ѵ������q^P{���n��
O��``+ �d��E>��S��yru��ʖZ	E�C 
�*;Me&R�Gɫ�*���p�qf͘���8��]�PQ�R)�%U����̓�N?�٥!������ϑ0�w�%���">��
�|k��$�����ϯ�L�qyr�9� ��\F�Q��!E�|��DY2�i�aP4��=}@�H������� 1���a�夆�ݣJ����4���,y"�����u_�����l�6_U�C}� :��o^}�U�m��5���i�1E��
�|I�&�c��nV�\ρ����Q�i�I� ����K�|���`e�1�� �C5��D�>�\��4`�@�I4&mf4-�yZj� @j��?�#��8/����f���ZIU��d�_d��ؤ��WG�۴i�!�M4�~E/��� ��a�
�B��¸� 5�dO�X0�%%���~�҂��!�ǣ�-2�|��4�9�0���b��X������o*�; @�~��7;�0cƌ`ĈU@� D}>�A�a&�(���u ԦTĵ	["P`����D<A\}�
�y����x�M�<����"6������q���UEȰI��u�I<�P�	
ӳ��CR]�Mv�|�����w�S^[RRR�+͂Y�&�b1F}��|������tp�?�.$0D���MA�O� �����\��$�G<�`f��'yn�5����u�H>��5P�8Ym���C� H�`���I�Ha��c��I�q fΜY�]X�f<��>���Ft!�HZu�ån�{�Ə�w��+D��昼ޣ�I�Խ�-��s��	X�S΋�Lۜl�'�OF�<>��"e0����W�C�m���W�J|�c���� `���F�%��n�CIk r�s#4U�u!u��R��`�%�+���/���R[�p��^-�,�9�����g� �sF�������aC�5(!�Q�H	 Fk{��I7���Coa+N�ט��Y& �q�|'�x(B4�t��M�J1��$)��KR[��͒9s��{�;��{  >�Cb�X�s'�n��Ga b� �%���qS���&<���upj�S �0��yFK�����Y8@�x+d7ׇP��q̈4 �� $��ɼ�%A�C�:�fTC��e��xWx�Aռ�UBM�\Mr!-I|�~0�}��'�j��r@�qh�g���f��A*5�3i��
�T�Mf�'ϧX+Ɏ��n�&hfr��g|6fd�� �/�����J����Sو��+M'�E�n"��1�&��֙�յ2VځӇ��`���M+'�v�@%%o[�ע���2I���p=�����Bei�$H��I�p������65����kCe��N�Uf�:	�^��MA�s����Q,���t]���B��*(�*v�)�,�0��*�N�^"\�%��D�v}I�2[�����A�]��5MSP-��RH�ˇ��U�w� �|gը-�T��N��*�Y_g|���>��c��ϩ$c�:]8��A ���51/�*���6)�3\^���EW�>^&�"�GN3U%Ve|\9=�>�:��kW��F�z`����IH�)h��~����I
�;i#���:�h1줁��Q�>�Wee�.�_�D�g����n����-��O[ j�ɺJJ�'MP�4���|o
��^�4�S����Q ��(��ɨ����"igp%ͅ@�t������j�o��$D�:�A �=C|*T�ad��gMD�� I�<�����3��:�ƿ�3g��:F�]��e��8Bȣ�P[/$��(�,�*4R��~�
�G3h#�պZY5s����+���(��ko�$��K�K2b|�,p_�������P����Y��H��|*���s��w���{}�"Mb2b�3��&q�̈́Y?��U]��U0H����M���}�a��r����Gwq���9�����٠�dU����>+t�'�b�B�O�E����:$�gb����7h߾���~_�V�t�O�`��Pp�Q�	�� ��s\�h+k�}�w�O��q� 1Z���pl���1�b}�jY�ȏ#���&`�}\A�r #�w���"���4|��1�P�8 I}����	4߳�-双.b�:�扫RW5�!%�Z��^���\� �P�~��w��j��i� ��ԩS����r�'����HRP�dK��f��J�|�BS]���	w�g���G���`Θ���e����Bei/D�h�
��m۶�K�U��E����>��;�^7�"�~ppg$'���*�����͘�5����Wݱ�)A����3�RR(������ɳ��>�hai�.]��c�^ �Z��\��-'�����'�4����h��)��p��x>f0 ����.E>��!�8N��{�k��Y
 P ��o.��eA�>}�''��-��oɘ�(VH�.j�h<ҡ�aJm�?��*#K��V��U��;T����=�P���1l$ 9@x���w1�Td��v�^L�NgX���i6r���9��|�M)-�/�A�� �4����6��*=��f���o�s��U��E�h�D����f��8����]�Q��#!�=�f�9rȇtT�ֹ��;�)r~�j�*U�D"\��u��U�,�+�s�O#���̐���_�#Fi{@����Ӑ�����m)�@�gw9��j _�@{ ��J�yJ�T�ϊ[�#k� %���q<SS�<[���Z|<}OE�
*��w�A�w�a��bg|�cl]���0W9:(��|����Cs
��нT���$������񽰴�C܏�	@�����p�Ӕ��D�P>�pedw	��S�������uh��O��;�[���$��`Ӏ��鐐4�c�6����y�W9I��hZ�x���w��\ep��(�j�W$Z�髦 m�O��U�Ǎ1����
��u�U�o�U��N�IS���x����^Kj�1T��]�S��)fdx	��>W�$�  �ر4�������7�����W�7��k��4���2�m
EZdgP��򎠴#�>bk��:x�� wP0ri�(#"f�a踇v$ݜ��k���|�@Rⴺ��:aGF��xS��*B�HYc���#3͚�꒞:�ON�v>`�m���u�3�4O���j��`�ʸ���5	Px݊�(Җ��'U�� ��TO^��	�S�fkUH��k�Rl�T���q�(�
�QI�b�>��H�[��y�c(���cS�9>O��a��t�dxp��/���F���u�@E��!y������WI�P�S���!�]�P�و?zo������=D퐊�$(�V�5�f+C��)6fKDI=$�����ZQ���i�:�?�]峲v 4��߯iA �@M����G�+hw%yk>'"T�O�txJ�\�1�������q�[o�̛7�]+�ܾ���et���3���z\�#�<�%T�c�h���5d��{5�ϮKPV@�ҿ~ϵH���S��0�Ƣ��[�nݩw��ʱ�4R#��\[�'� �%I3}05|`$�}����'�����ȢE��X�d�b�����^mڴ�}�!��7}���{�9�s}� �d�r�!�����7��z��I$�m�������7�xՐ!CF0�K���" ��0؃�5(�D�A:�@�(ݻw��g��s~��i��g<Xh`�8x��ۯ���q;��l'��F3��!�{.��?�s�9#�����_t��w�yǝ^^�^z�)��0iҤ�v��ѣGW�$W/���IYb��`؋l����6�!V6��	'������
C=��;��E6x{L�0a������_�� �~��6m��A�F0F�D����C�?�x$�O=���;v,~�7*=L�
 � ���h���B���(�
{�&퀄t̞={��ar�'v5L�۷w ]t�E��~��!=z��RRRRWrZ�@F�������kݔ�+������ߵkנ\L�����U�+*�&� �j׮]йsg'9�[+yO�)9A)T���q��-fZv�M7=A-}`�F���v}����m�nSLAH��X�@�����~�JZȈ�Q��f^p�_Y�$:w@PY���/�믿>0�v9���̢Nj��B#RM� ��I����:�(W���3�Ğ�&@��϶{����\Px`&!آ��u�̹����o�!�&fC=�0�`�����u��&�`n0Q-�x饗�hw��ͥ]h�,�?餓�Pq�00� ��Yj���Z���y�Fx���Ql�ǝ��{�]w]��%�' �{�`�x���8R��@���GUl�=��=d[�ar)�ax`�ݶ���ٖ���"fR#ý�q�#Q;�4��D�;n�8�R�����s++��S ��?qO�d�����ĉ+F��(� ��C*��n'�<3�Zy_֖f��gy���0��\��D@��!M?����Ix)�cz{�M�ш�Z�P�5��j�^%��.(��D��4�ei�"a<��/t���>���&9�F9@0�G�� ᚰ������/w ����(f�ۻ���O�ҨQ��~����&��8��Ӄ�����q�{�΍��<���Nv��� <�2����R�+2����xa�%l�B��4���R\`���gt�����|�1V	�(1jqA�^$�gR��U�����K.�i�<�#^�ڄ�ô7��gϞ[xЍb¸]�*}B�a����:����<�Lg�Ѓ��CPS�A�~�W���fG;N#�j��`���D�NbDX���h(��Հ@z»��7�	'1i/�8FصH$�M
`y&�g߾}�d��ƣOz���B2�=�X��ɓ36@n5�ؐy\� 4Q8��Y�f���� �H�G�� ��[�<��W����(�{0�JOy)���u��ô��|�&U#f��}�k��r����� �c��#�<2y���gϙ3g	jRg�����n�m����>��.��Ӫ";0�w�=�d,¼�D��uv�ٓ�&!�L��t;v� $0���S%�D���r�k$4ʠ�t�*�:ˈc�]:>\I.U�7�?�^E��}"�;����l!.���O<�R��n�i<���3�~���� -̀w�ǆ�����JeUftc	#�?�i��iR�.�5�����Lz�M��و��`<+�$��d��*���|�V���ɋi�/z�V��(�/�ÓO���I���iչ�D�b�Is��>��Y4N:�̾����90<�'��i]t�8���<���ۉ1�qJ��ngaï�D�`E}/<b5]�f��R6I?01�cƌ��.�6�ŵ���Q�Ǡ��EƧ��2�T8�K�T�X�*��{P�ǀ#Eg��Z�`��Tr�	�\���ۅ�'�.0T�	q��ۀ����j�4@��9[imv�{l �4j�Q8D�0݋w��a �@J���G���g�q�Ku �C�U���x��;�&Mr���Q�.��.rȇ�0)DY+��D��s.-�g+rV%%� d+���q�\�H�?�3σ ls��@�zZ�A�\K1[)�\���0GF{�9WH���͖��ҨNiPM�&D�@@����@��0Ɠ�ɖ0Du�N��N�YaybR�xY�آ��D���ǹ������M�:E~�h���
���~�(F-I�p����� �q���)�:'w�~`�,&�`"��-��{H����k��*!d��Ue�Zp	Y?�gkR#��«c�Z�� �ֵI���"�FBRޙ�њ�C��(�J6u���$ �������o�Q��)�LF�E�������&-�٨��$b�/���]�}��E9�7��իK�֭��=����M�6�>��L�Z�t�I��}�֬Y�м�'�>�Poq�Yg���~������ꁕ+W~����Z�h�;���|�$�y{o�}�6�ѽ������~����XB��������w6P֔���΢��I$�m۶�`��]��m�y�����&}��mk`��{me�Sbjh(�:�d��,9��ka���;�z�UW�%A)B}��\j�� �ر�X��ǒ&�j��ך��qէ�vZF�`Tt�-�4�ٳ�R�j�c`T�NS'�`?Pe`���Nc�� 1��Z?��W_ml������W܋�A�ٍm�<�m@�}�Lm=8N�7�xc�5�n�쇮C%e��v�����j`XO�TH�Q= F���R`TH�Q= F���R`TH�Q= F���R`TH�Q= F��m)�����Tk��Zo�Ϧ1�k���_�mbPk���k�ƍE�5ڪ��Aiii���.kE���>+
���R�ImU�����mT�hK���V�ZUԲeKݫ��E�������:�+،�??JD��    IEND�B`�PK
     `+�[�c��f  �f  /   images/c88b2895-5e8b-4a57-9f9a-b80dd50058b1.png�PNG

   IHDR  �  �   ��ߊ  TiCCPICC Profile  x�c``RI,(�aa``��+)
rwR���R`����b
����>@%0|����/��:%5�I�^��b��Ջ�D������d ��S��JS�l����):
Ȟb�C�@�$�XMH�3�}�VH�H�����IBOGbC�n��ₜ�J� c���Ԋ�_PY���Q���Tϼd=#CsP�CT�%���X�}�����ߍ�������k'BLÂ�A�����΂ĢD�33��10|Z����� |�'�8��,������z����j��N��������.j���p  !e�2���   	pHYs  %  %IR$�   xeXIfII*            (           J       R   i�    Z       %     %      �    o  �           a���  �zTXtRaw profile type icc  x��S[n�0��)z^�8~$R��b;^eW�J�ё"�@`H�n-|DI�D��@ȴ�v=L�"�	�s,`�ۮ��z����"H����pz����3�ͬ,9&�h'�tN9#���(���d>CQ�h�|q�k��R�R����mOi�q�6�Z�ܶ=���C�>hrK$>���U`�͚t3�s;����%�S�T�c��\���~�y§b�_"%�G"a=}J�H����|)�Ni����2��yl�c���r�E��|�7$��8��s���.PJ����
��wq�8��P'��j����[ܞ�c2����g�+��|����RM�=�c2gҥl��ϞauTh���҈�\�z���줡㜥   %tEXtdate:create 2020-01-31T21:31:09+00:00��y{   %tEXtdate:modify 2020-01-31T21:31:00+00:00	�   tEXtexif:ExifOffset 90Y�ޛ   tEXtexif:PixelXDimension 1391c�   tEXtexif:PixelYDimension 800�요   (tEXticc:copyright Copyright Apple Inc., 2017���   tEXticc:description Display P3�y��  a�IDATx���|SU���M�M��ޣ {��Dq�����~�V*�~���(���(�"{�Q6-�-�M�{�'I�M������K��{onn���cU{�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!@��-[a츱�aC�5?�q8�^ݺ"���0�
�"���l�a���>C��p���Oo��vn����"��mE�9F�1\���?ۛ�����(:���c�X���_wlP(�ʔ{���=��|+��#}�Y��mo�w��k��]�o�������?�O�0�?���'�Q���W?s��3��"Sڶo�dՊ�}�I���i�f����gf^�t8Z������^d�g`���>�n�q�0K���k|=Ϗ���5�1��}���I0�p]�y��U��'3r��~'_{���G���ߢ��h������1o��v�#�����޵{�I��z�}Պ�ged��x0'""��!;;�߁�������t8�ADDDՎ��4���N����E�l4"""��L�����QQ���ԿTP�UK���	���sn������BDDDՓ}����{�������H/�=��|!'""�c�4a��sh׮ݔ�#F���u�}�?_+.q��p8PPP��o�O���m+�p���DDDG�}ǎ툯0;+k����C���PA܉��\��+z��I#<r䑓�\y���O5�Q�?�^D��R]�]R<�5k����q֦=11Q�s�*Yǖ�Ull,���0�C�Y6'"�`V|֠g�HKKS�o����T���Ύr���������GXd$���(T�:����=3+Y*��D�~2+3K��H�h#"���sx���_����`:͈�����O��;r��"""
f����6.��p�)�ggg��oDDD�����R�7Mgx�'�����"""
n�Cii����p:M{�'��]��QP3��SSѼE�8���,�3�:gOݟ�F��:�������y�
�DDD���";+;ơzI2�kff&���(��j����H�4�L��at""�`&��:���K@/3�^�a�Љ����nC����E��J膻��0���(���*w�^���(@VV���(���*����:��D^^>���(����p�Yo`� ��;w@/;�����FDDD�Mr�0��mPP�ϵЉ����iB��'ԭiՆ.������Q�V�%""�Qt/w���^J�&�΀NDD����m6È𶁴�{+�Qp�/^�T���t""��g߾m�*���6�Q𲧤�H������]��1�'���i��*w""��g����m*`��r���/��Ä�m�����NDD���3��G@g�;Q�S%�Æ����˝��(��3�����G����ΐNDD�Lس23��i�I��S��)U�ge���'{�3{NN�
����%�;Ճ������zdDD�i��K�DDDA�T=&&Ff��Н*�;Y�NDD�L{xD�t�S�:M�~Q��l6;|T�;�&L�Љ����=L��*w�Su"""
^v�a�ax�&�܉�����0�QN	�U�DDDA�T�\J�׉e���U�DDD��.K�|tV�3�|�i�̽t�U�DDDA��%���F��8tV��rK��U�DDDǀ�����t�K���˝��(���K�z���X���(��E�{	��7���t�,��ʝ��(�ٝO	�:��:űʝ��(hI����4�r��YB'""
fv��a�iz	�n?7�)���(�ٝ�sm��NDD��r���SQ�n��^�n��GDD�쐕�L��T07Љ����)U�J8|�r�Nq�DDDA�n+/�K�g@����<����@=?""�F��0;�*��乸ҵ033ii��k�.$'�@jj*>�����9	�QQ��S�ѨQC4k��6���\���1%>�|��%rpq��+�*3��?V�Y�?���Eb��-طo/<���<W�C=��,|��\`�!6&u��C�V�ЫWO0 }��A�&�f�1�Qȑ��i[�I@���p�{�W�܌���X�z5���;�:��V�ޯJ��(��Q�w�{�>)ͧ�Ė���/s0i�$t8�#�=�\|���ܹ��v��D$<�����pU���Ʉi7`��r��s�C��\�U�^�x1�����n�n٬��E�ۆ�)����`�E���Oq��W���GR���yv"��\�g.~��w|��g���;п_?�i`7нN��¹�}�\�-[�b����Gcǎ�p�W�����=轢������i�O��P\p���������O���u����拓�'�S��o�T!����>���2>�͘����3������_��p���T�Y���tf������ذq#��nԉ�cP'��'������ix뭷�|�2]�Y�^�z���'��2���V�{!�Pz^�0���*RS�µ��Gݷg��g'a��Mw���������{���#R�۟���#G���x䑇Ѡ~}u"
Zy���7o&��f͚���8��yHo���;�1��&��ޔ�y~&M�\�f��`�
���hܸZ�h�:�E˖z8Z�*UGGG#7'�z8ۆ�n�:lݲU�TU�[�Z�QV�a����HOKǨQ#� 1�A������K�,��߁�����Qi�tn��lC�C�����g�><����!??�oF׵kԸ1����3���&M��v�ڈ�{o���b�ʕ�a�:�~�:w���Gf ?/~�$��'�@LT�:�Ca�^��,���eʐ�0���or�gf��_�G*��`���9Q'>�>n��V=��v�Z�ϖ�|/C:�5i�H?�~n��L�<S>�\��S�5��s���[h׮n��z�~Y�(�2+&K�"��n�f9U��W\�Á�U	x���s���Űa�p�9�v\-�_+Ƴ�L�׭Kg�;��|2��֮�ù�J������ѱc�ؿ?K�DD!Nt�s����!�{Μ_���~�2�M�!����#г[7�_+O���/�	u�b��aX�l)�36�6��ѥK�� "�P�c�i7���*w]-̀^�n�ꫯb�d�z��L����p�Wb���hռy�Kƞ��u�@����~�H޶�����{�	�_xK�DD!ɕ�۝�i���q����0��)���_Q����p�����FTI0/N�}�Yg�����ǟ@���(�/3p�@*�y�m�4` ��cP'"
9�����rg��#���,F�9Y�.;ѵ[�G�M�VG%p��,2����/�L񲕁?���?���%]""
I�L�곛�k�Ԛ]B����i_c�jo��L������ރ^=z�R�'�N݃~�os�o�X��3��0s�L�{�DFDT��y�"X�X���x�����X]��:Ne��.��� ״������͞�}���[8�2{�u@|�ٸ��K�ɲ'8�w�{���O��������m=�c���xbP�p�ٟrss�����f��u&"B=�ߞ��y�v����y���Cn^���OV}���a+���N�[�8r��!�1�(ǲ��V�Nq�|����EFxȹʵ)p�>[u�rm��ץ���u}]�����OC��:����9�?���"��\}��ˌ���^��Пc�{�hU��)}>޶�R�5RT�y�s�C~J�@~�V�,�[9C�����57"��_@��U�?ϙ��+V�ۭ%cͯ��zԍ�?�7�/&:�^v	�M��C�0���-lطo�-_���Y"v���X�vV�Y��6`��]f��S�P�,�B�Z�ШQ#�n��:u�q�uD�����JZF233��]ۺ		:�*�>��)�f���X�x֩��s�N�I�##"�{hѲ:v�^�{����k�}^ŏ�r�*,Z�k�5۵k���t@����36o��{�@��]о];Ԋ�����u�8��W�3K��t�	�H��r��!���Q�X������u���lչ5m��}ջW/���u�9��a��5X�p�>Ύ;�q$C�����M�4E��ѭ[7$%��k U��{2��3-=[�l�K!�9n۶�))�����C��(�OL�3A��E�ΝѦMk�V���~�:��.�����MIJ�)���+T���6mB�>y��zK�D��f͛��,�u���㐘X��ZT��gVvv���}<p����_�X�����)�T��21g�(��t���k�8t�(���S_om�&���O<�R�>}�]}�������֊����m����ޭ{w�P��螛�J|���f̘����[�nEzz�����u^��t ���x�s�98��S�P%���w���x���٧��U8r%���5l�/��2ڵiS���C�o������
+T�g��>އ�";4h����õ�^�A�����8;U��n�����/�l�2���w/�k����(u�p�)����N>�$�R�ؑ^�/���<iR��r]d��_��*Hz����ᇙ��/�x�b��>>_�͎z�����5�\�s�g[O��J��`��F�ܰdrd�$���q�#T�T�9���u�	�$xUU��\�M���5�'���X�d����Hp�uT�.�6P�]O�ё"��*�W6�{�U�~1#G�ҁ�0��j�L�#�<Rbd�<������ս>Uw�MNNF���zoR����Z�.�1�sp��#�}{���� ���'��o��H׌2*��ґ��,X6�����?��v��#����.�С�)��^��C�`�l�R������;�ޱ�A.ǭ���*�4h�=z�K1�tP���>��U�ɫ3U[����{����z�g����t��.��c�JXd:ܛo�Y�ʮ'� ��%�ϕ�X��$�9[�
y���N��r��z�8�ޭ2�|��~��^v)U�gR�ve�]�b���ٳ����:���q�*w{�6|���0�Ǚ�Zɇ�J�͎��T%���_��u���<�+�ȿ����_�sGvv�_�+�lʾ��5�����y��ǟxݺv-���I�����B��Z�'_�.w�ځi_}�9?��ŗ\��{I����'g�k�|���z9ϕ+W�i���-�����nՏg�T���p�������KGb�*����?�{���K���Uk���̾R�����'[[��>'�dIAa����G��o֙)��L��M�����Z[j�֬^�u��T&��ge�ԯ���(g�pKU0߽[� �=�%~�q�I�������5�گ�GZ����[=�m؀�^{��9N;{$�6%������/�E]�r�Z����5�m��֩��,ǘz� ^U��7����}(���\�;=���}lٲ�����]J������7'��^��=�ܯ��5sm�?5o���ά���:v���)푆V*4u��p����N����|���f�?c�u�!�_L�[�n����|��"�>� /���]ŏ��VJx�n�\��cǢo�^��r&�9�UeXe�sU�-//��<{s][ɠIFsŊ�駟�裏�_����2��-�S�-��⟩��]x��gT@��&��̊ٵ�̮Z��?���H,���>��I����6��x���r�#����D�Х�2���>���:wB��m�Ӗ���[*J>�9*Q{z���믿�^�)��2�J(2���ч�R�J�H<�!C�v'T�%���'�x����d�k����~����@?���B����3�{5j��4dee��2?E�q80��oUf-�Ox�<�$�*�9
o��ffT�|ſ���Gzo�3�up��8���J�/�_R���>������O���$}�+S%57�F���Ƕ-��f�x��r��0��iذ~=�}�\tᅺ�_�SXO���/�£�<Zl�)��m[6]��������۶n�NjA@�����:lM.��t�t�2[�зO�׉�:�\jf���C����໻����m���WJ�Y��d��bX�w��_�h!��^�����_���*ڋ�	Z�1�w����a�B^���t|߁�'U
�4q�Q��-,���1a�J�=U�9�����NJ��= �r]���1��W0��	�ζʼ�������yx�����K/�Nco��^;i(��?��@���u�ȑ#�h�#!����F����9�[f��zH��������|���ū��s��z�
���zg㪫�
�gYڌ�3K�b�c���+�������Ǚ?⥗�cܸ�������eR:����ǝ�Tk��g��Ѝ�bz͹xť��`Ϟ�^����B�.]t5o(]!OR4��Y:t6o� ��ê ^�~��8ӻw4k�u���UT�h��]z���˖��]	��=gö����Ï�k{�E��T�ק�~��%���#"Ѵi3�B]Su���7';�R��Ҕ�n���VS�JЎ||�ɧ8���|�
_/�]	hLl��h��m�"11QG����uo�;v�;�Yg|�T�H��E_�.�W����=u�4LU%9W{y���D�=M�4Vץ�>o�$��RSS�a�l޴I��[_W�2L�:_r�
��0�L0w]���u�4G����u��n2�Jz��]�V]�dx_�X����(��N8�_�������ȑ��v� ���N��B��I��K�.�3�����Qڵ7oެ۶�'|��C�.Fq6=���=�;�^�I�$��t�2L�<����\ރ|O۴i�{�K�HG�C��r�򹦧�y9w��LӁ��}s���c��A>�G���}��/��\=�7mܨ�[�d��%�ף�t�S�֭[6+��)s���2>�����ak2�H!�ک��H 5��_�|9�?5��`�Db���T%�W^y��#פtu���ԗW��M�:����k�Nx�;�oÓO<�F�h�8Ce�Ru tu�+
�R��ۯ/���J�v�ih�����̈;)q�P�9����oM�R�1�f�Ϟ{n֫���]7�
�u0��3p�:N�޽Ѥq#=��s9���6�k\�����}{���#Ìf��:��^��"�>R�s�v.
�a*A�ޣ7�P���[�j�;W���W�dΤcۤI�����e�	�34t�x̘�طgRS���v":�N9�\}�U�qӦMu	�s]dH�֭��ݷ�����W`���"C�O���}zW����3�ǘ����yp'��o�駝����,���!�1�S��߅�����Y�,2K�s�{]VN����y"����}��ΕΠի� g�u&.��b=�q�ƺ7���zA~>RTfm��%�����H�Qِ�o�}�]�pB=����m곸��{p�-7���]���;u������gj��Q#1��u?�Lɐİ��?��kf@�R�+���D6Х�P������*p_Ub'�|*~�a�q�@Ĩ���'9��x��W�������6g�l��X��mX�z%�W	�۪�Ѩa�J't�P�\��T%���;q뭷��JPQ�L�p))�҅<������>V��t�Q%�����[���x��Gq�E��P��8R"�ݳ�w�'��?��*SeyUR��N�m\�а�8T`�*�G��"�*�ȃ�Եi�Jp�+c�\��-[��u-q�
�R��
�e��B�u��l�kޢ�=4LW97�_��K�jת���ҹ���N�ñ��?��IUb���{�͚4���^֬߀ѣ�ww����'�n��s�mh�2c��:��&������Izʿ8�E/�(ٰr�r�S�O|�Mԫ�P�{]�냅�Q������O�Ї���멈s�m�y2��|�q��aʔ)5r�:�����$C�j�9��nE�Bf��Gq��Յ���2����4��>A�I	��zg�'�q��ϬH�Zž�b���u���1}��qc�}˻C<��&g<�[��c�=�i_M��8B�)�|�ɧx���T�V�6j�Q�G��7�Ꜽ���R%����믿�vxz���T��^��K�DwZ�VaoǑ`0d�`]���۱g�.��lܸIWG׫�$.֊�K|ݺ��8����I����[Ǥ$<���X�n}���H&�ƽ8�{��1ͅ-���?U�1c���nƖ�-�c`��d=#�t���a�ĉX��[�թJ��1b�H]����ɞ�V_]O�II��V�	V��3f`�*9ߦ2��Q��J��u�_��T�3�9?o��!�Ho��]Z��~oSKK��|��:��^��X锸��Zzj|j^�9bz.w��멚�)N:rI��+�['P2�HL%&�6�i�ܵ��.2K5�u7p� =L+�]�#z�����J��t5���H{�|�ǨK/��\gW{�C���]����ݯl'��I�ᤷ�*wk�.=��`^ѡ���:^t�:�D�g=6X�z�J�+��;�w�q��ů"ץW������1F�t}��H�[O<�.8�����{��N��T`�>��C�aݺu8EmW���]���-��V�e��O>����+0��g���L{����t�{�+6��hˬ��z(��g֥〥)�|��a�葅����h*�I��K/�K�,յVs�H��c��	�N���Ց]���g��m�vM_d�p/SfVWs~��ŋ�[0�j��숃���V�ǞxLw[�'�([)�l~��ttx�� u��8��tӍ�ڸ��A�L�������mE��ύ7݄s�����9IIpР���O�x���1t�=iK'��֝�RʖL�ۓ�Fj�>x���J\~�e>k,���*�O�4��C("7JG+����S�#S�Ju�Ν�U���|�M�A�n+̋�Ƌ/�Pw}a����$C}��1�����Nt�p�Zb���W^#�j�G�)S�m�U��y�f�?p $k,��Ͱ�۳�&��KG���l[�V��P�i)��~��7�Y��~i�'�T.��SN�|;�����}�}�a���k�������s7�p�n���qM=%�u�]W���:w�&M���`��G'Z�l��.��2:$�~b}��f���A]�&"#�����)�Oj�V�Z�:�y�xm�>C�u�Ǒ���w�5)P����蒤�NS�*	����2��:wŭ�ݪ�D��.���o���f��.�+K��e:��^�\���0��$��a�k׮���B�{��]��Cꚻ:�ѱbJ��M&a.GMkC�_:Qe����B�+�ۄ�y���$\q���L��OI�.��=��?�:�X�b��5hr�9�<����uĀJ�엨J;�u@_�u�SO;�U��� �p��z���L��U-��V�[a���+���ؼE/S|��s��ǣg��*�JB����m�uQ��^�s��Uj+�2�aa�ͼC��z\�ަuk�{޹z� ��ҿ�.�M���[�5h�Hw@�L�kO@�*yw��	�M�n����̬��б�>k��]/�jb�db��[J�6�`�=D���3�:�[�
h��Kz��w�y�c�UU����0�!�^}UB)=g+P"UF�a��^����r�#��.N����72C��- �>=z�@�J���u��$��ye�лO�J��/���KH��uY�C:�z��(���3o�<����^v��F���,u��x�	i�8p &�5�G��ۇ*�"�Kf�c����(�;YAN'���*s��"1tL�v���u9�����M�>f��ܵL�*�W�L�b���:2ɔ���B�F�4i}�7\�c,XY�K�}9���B:]�t��{��_�׶BSO��1 �Ԇ���qb�>/A+�g��IV�mV�5�ef�U������U+Cw2S׿V-�m��zQ_v�ك��Vx}�k�nh߾j�Hr7M<����J&ϑ9�s�n��^r�ש�������"B���VMcNgH��Ւ����yU��n��sTt�ϭ$G*������٧�`)Î��z�Y���j��ڷw���n٪�l.=����� �+KWT��{�ԓ�4k��e�����H:�1u"ݮ]�J��}]t3���A�?�l��%ǩlgTڶ�ː@���;�`0���I����K[7o�|�y�w53+���m�Fe
7O�d�$3lU�.�Ռot4�_˫r����$ш�Yb1��4W�Ȕ���ɬ�i�u}TsV��]R�����<�b�0��;v�eJ��(qq�t'�ʒ�k�')=���y?�u*�픡��&ޛD\%t9Ve�U��쨌M�7##����=\��[Uj�_��d`�e|v�ڭgᓀ~dLDFE�q��Nz%�*ڼ-��b��/�$t���g���3�I�!���*s�I[]%�Ƃ��͝��Y��4C��I�oU�	��!+�Ig$�6:�t����W+N=j��IЊ�=�Z��k\�V2TU-Zer�t��*S)&	�nݢ�}�H&j��=���_�HaS��L�*�Y��?x�S�W�8��A�@L:TD������YCg&~U���JJ2��M�����۷O�U�w��`���4�eɼ޲�CU/BӴi]��(�8��;��[��.�?G��X�(U:�N�H���Q��H�������܇�}޷G��YO�����Ǐ�믿T�o��ѽ��z�����d�1�F��(8I	�^4o�L��]KJ����MWz]=��i�suj);�7�����/�yJ�99e�2�:Oα2w�T�JG��&�;F5J�$�v42 R"=��M��R�&��x#�k2��q6e�&5��؏�d����j�k�#�\m�5�m�Q�ƈ�]���:�i{�w��`&��[�M�*>
U��1���Idsr+7,�nS�+�����]M��W���e<���X�����z�Uѩ��jH	���n����dLm�zu�o���.;�Ɂ������O���V��G��*@Ib���C���l5s��J.�J�*��<�f"W]HG���e��@u�*��d�;Y����r{��jh@o�X퓒�F�3^�kv$Y6P��7o�3e5o��u�`>?��>�P`��+\��U���Q�*��SNUC�1G9��qk%�Nӽ�0���pk���a��򎥚�gϞ�V�;���˗/׳N�`��ʒ�F^}�5|��7�бz��޽{��%�KOfo3_IU��`)�hf��0HR��g=9�!c��5>�'
��L���C�v�\�3G�f3u���@T1�Yn���5��^*�K`?�a=fu��eض-�:f��#%g�/%EO��c�6����l��ZĐ�3z��K/����)�N�p"	��(�H�`)�W5�s����OT͝Oǎs��
M�?��$&�?f��:U0��8ӟznC�u:N�n[`��(�mHNކ�9�]�]��7�B<�*=Ʒmݬ���ڷo�zi����A�p~PzȘ*�gdT}�_��Z+�و���Ы��`^+�{'O�0J�\h�8��TT�Mu�H�ʽRU}'�zY����?���_�e��]	؇���%����t򓕮�ԫ[O�Ѷ��(��Ν;u�۪v�59���v��1̍f63�٤������Y����mT�:1������]޵Ls������U���v���_�d�R8�rF[�nÌ߫�J�̭>RS�v*���� Q�������*K:ffe!.6�J����]�N�L*Svq9������m�2��Uږ����۷��~�]���R����ft���;�-^��k���Æ�;vbʔ/зO�c6C��gb����|�z���#q֠Az-i�O�^�zhּ6m�^�e�Mz�}\_s-������6��u2;�$x�����BNN�I�d�����K.�Z�%yd^�#��n�Ն^3'��%k�r�U)}���^��u��]vN9i�Q�b��yr2>��s���d6�����mZ���O�܇gq����1��_,�"��u�֣e��
[�n�ƍ��mXY�֭u��(ڨ�^�nv�*��|#d	S�z������H���.���R� 'AIa�������������t�m6\~�e��/�q�:��ٰ=y^z�%t萄���G�)�L@1y��X��?�7��s���0{;�������`�1�Х��Qe
N+LtE�i�쟱{��>���٫�^~��ߊ �y���T@�a񬁕+WaŊ�8픓z\��������s�~��*cQ6@�&MФqc�h���:�����N~3u�	[yU�5��]�}�Νqɥ�`��qz&'+�&M������ȣ�e�i�l���{((��L&�hּ��'A��9���[q۱}�f�*���]wމvm����ٻ3�NG>���ckšO�����}'R �=$�����s����>uON�2����.\�_���Ԕ�أ�d/:��]�>�p�'�se6s����巽BL��:/l�
�W]}��6�[��e����+HHH��s"�ë얔m�*�?�̳ػ�[�z"��.��{�*w�R��ۯ�;��f����0u�T64`S�����|K/���ŤI��úw>ё����3�w��S8�����^ݗ�^���k ��r�ÙY���U0���;��2�UI=�S]�h�����z�I�YN�l2����~�m�a�S��p���؟��}N_��o����W�|�^�/��,^���dNt��7�|�.e�:ݎ^��?�|UZ����&m�'N���N9�J�/9�e+V���^Cf�� ({+JO�s�=͛5�B
$��ڧo�4�GX�1�=9/�8mޜ����W|e�Q���o�nW;g�uV��i��ЭÏ4�y�d����Ə:sJ"\݀7� ��*O��+/��6]���O�^<p?ڵi��	D ����3Ĩ��x��`����E�.]�>�Yg���y�υU_��[6���c�L%rmZ�:���j߇^��*�[�V�hѪ.��|]�
���O��UW_�y��!+Ӻs܌�CR�x��'sd�Lxz��^�cǎՙ~o��N���5ADd�^��j1���<�Kܒ%�ωe@p�v�����ª���n�{�X6d��a�oa��ŸM��SZ������6�I]6mقw�yWW��L���NJ�W_}���
�۞eY
��oT���*�;�����J4�0t�0�ya:�kW�DN��c�.<��p|�ŗ��l�$,,�^{-�w��`NU��s��_���V�z~~�|��G������n|���ҫ�ɧ��?{�j�v��|��hP�~���ccbi�?��}���3rM����t�SB7ٖQ��XRU7��0l�CؽSz�Z}A}����O=���'�����y��'�u�V��c^r9��,lܸ�~����5V�Ҭ����X�W<s }����}���~��3>��S��e%��_���}��GqҀ�^�&��Zi..Z�J*���7��/�p��	'���E�������{J��}��WGw��.:s�����q�
�����"G%_��Q����g��Y::{�ٺ�����w����<k�̾t�����z�T��n_���N�e�U�Zn	ݕ蒇L6q�嗫l�	��jއ��Ds~�	���;Z�j�~���G�����84i�1��:�K)\������{�`ٲ�X�d�.�oS9��Y�|��LO��1ϣm����}݄x�Y�իWc��%�J䤏��ٳ�f�\}�5�����!)Ig ��N:mڼ	ӿ��>�[6m.�WYN�l��?��^�`NUi����{���#��]z���eMM����q���~-[�@���}f��`��ǧ�->��l\���8ѵ{<��Cz\zM����j�ɢ֭�z���];q�}`��i�ԩ���9����ߥ�q�1��+�ak�r���6`�ZD����_�uz���F`�~�+odC��v�����٧vĨĠN|��)�H@�ǲT@Vw�����}�߳|�I'�ŗơO�^���ӫWO�5��s�^��[-Į�;0�����T/5+��e<�L#����g��)Y�p!�'o��᫆����`��0���@T��b-*(�y�ر};�y�/C@��z���xRe�'O���w��4j�	ut'���=m�r����زe�*I�.��{�F���SO���WMIg�}Ʃz+U��s�^�ru2���4���as��2q�i������G��T@/�#�蚢*\����$��z��c\r�˗-��Jg�[��d!�Çӽl��J���0���{�y1�Yt��9 7�9C�F���裏b��M�ԥ��k�v��~�=�UxD�c����<��Ư��M�5�SÇ��T����hеR*0H&2?� ���C�v�m�#遽i�z���˯��uהφ������3#��y�&x��q�X���d������u2
���X|�\������{�a���HP����z�Q^���ß�Rsx��e�^�6mZc��Q�q��ɖ��\+o�:W�L�ÿ��[q��w�I�FKdH��a�����ß��E���^)z����I���ʕ[�ҵ�J܆�63���&%ntlɽ�X}wF??J��ߞ�6�I/k�Mi�W��*�+�[^F���mݦ-�����
�\�����G��X����f
�))ػo��Ŧj�
��k����={b�ĉ��������H�|=�ze��W��SO;��s7�W���$��;g�^Fv�8���-2����U�9�s��:�	���K����ݺu�Čp�3���^��:�=��Ӻ���W^����aZ� X�E�ʻ���=22��q�}�����DU�]N_�#�=���{?v�H��A����HNN>f+\)���ˣ�����?��ުґCf�[�j5������G���!O�[OO[y�5W��s��OH�۽kL��:��x������,l.�H�M���O���O9�]w�^�F&�����^!N����5Z��W�������@�S�Z4���q��^��z�Ksp�	�>����*�e���G~y]lt4n��z=c�dοV���7��~?3��C���
�Q1�ر��Tw���6jРR���Ɏ�{��^�Z���bu<��qD��Is�|��F��}\(oi���9nӦ��=Opv�A�Н�����Ti����õ�K�L���m.���lݲUw�������HH�G�vmq�	'b��A�ӻ7��M�[�*Ty_҃]ޓ�������3�`�?ر}������К�fG�
�mU�\f�2dN:i �={+}��^�[�e�v:�zᜰ��Wmʾ���t�ֽ�LWr��I�V�!5r���֭[�kWu���Ǒ��S�Jur��=�d�%�v��!`��ʔ��{�,�w9���� ̋.׿Es�믎Ӷm�A�Hy�:��2r�sz����9?��ʕ+�����ɽe\
Oa���Eb�D����w.NS%r����Vi�٣�
n9% ��e��/=���tb릮yZڡ��/Sjk���W�\i^�fK��|���i�Oزy3���c��B��Zj3dTP||�����K����]],�J���մNG�s��gC�t�8�3t�;v"y{�^&TƖ������Y���HH�ڵ�PO���5k�\y�W]�fw���[�9��&w���ur�v�Y�F�N�e��Y%#=]�Ws�$*�j��^f��ر:w�W��#d����׫�	Z2���$�뮻���V"""W��+�I���>����QQQ~�ŕ��qϊ]�#>@���S�/�r�p��}e�#������-7�d��|b��+}lԵ�N����6m�ڵk�z��}�����lnn���bս.�=˒��ڵC'��v�{�Z�Z�
��s;��S��w�-kO�\�����S�|��/-�%� _��C�:�����Sqݮ

�����~%'�:u�ѨQC4i�T��1�2�S�
Ԭr�"�W݌�*ˣg����ِ\���5���@$��A)J%J2�Qj�����_��%�o��>�]� C��2w�zߒ ��� ��Ë����}�u�Dӓp�:�ʪ���qU{�o�VD�=��������"�LU}��qq�Q��)�/�I���&=ⳳ���ס�}��$�(:yHf˰�O�H/����r�;P�7��aUu<O�Tc��Q�9��k������΀^)f�K)C�\����b?�w,��#��L�im/��;�hݥ��8��|��8ގ)�ňp�z�����<��58��0K���0�~L��6�@;�\{u�yy�PM����Ni��f7����YB'""
f�S\�[y:�Q�ѝ8�)������^����3�-ӯ6�|v�#""
b���������(�ٝN��ֈ���7=S\�[�,HN�Љ������W~	]�9:����T:v���3M�r'"":�����,�Tn�7+�O"""
�K�ݯ8-%tFt""��d��m�::QPR1����DDDAKW��UBg�8""��e��˝Et""��U�:#:QP���U��8t""�`&U�~lU�?"""
F��ΈNDD�̊��3�)݆ι܉���;��~e/w""�����,�NDD�L��YB'""
jXm�m�DDD��"���������r�z�DDD՞S�r�5""����U*�}�k�r'""
ZR���VN�f,'""
fz�5?7eX'""
V�ߋ�0�'��,�U{�˧2�5?�r�܉�����m�r'""
b��U��DDDA��Nq�����(��~W�Q�b�;Q�Ǚ∈�B g�#""
~�C�˧2�+��^��DDDA���2DDD�ʏ�\�L��NDD���ΨNDD�����*w""���*w""�`�ʝ��(p�8""����kb=S+'�܉��B ;�U\m������K�p.w""�����\�DDD���X�U�DDDA��Q��LqDDD!����,DDD�*�˝m�DDDA�ɉe�������CgX'""
R�
T�Q�͉e���B��m�&�܉������6t"""
F�U��Gk��DDD����܉����
t�#""�`���WЉ����Dh�m��(񃈈���aT$��UBw8�HKK�!�p���� �`PS
Q���c�=�l����j���둓��ז�n��0l�C��Wæ�5�������]8
�������p����*�&6���e��-�8\yS~U��^�t1����h2�g�.��6��sDDDt�I��f4��&��� ""��JJ�:�烈���+UB7��͖n:�� ""��Hfsأ��ege�U;6�-3:::�^�n��������{�g��0=""�I&������K���;w$�Өqӻ<�t^^^/�4cTD��u�ƪ�3*8���c:1ϑ��g�#|���g��OF��x���$�����jժ�y�����W�<l��k�ŧ�O����;v����LP�F��]mn�G���E��l6�&m�v��0�æ�`ap�4�����rd��ϫXf��Ta���
�+����ſ�F�_JoWl����l�	�Q�k1׉x����󇢿B�8*�g�J����b{/���}����(:f��Qxn(���.u��{�`[�~���0T�.b�ҥ�{v�
/���G���NC�&M�T�^n7TWr�֬Y����[f�������=��ILl�o�Nɟ�f��MX�<[Q��}y�~����1�\4%�Y�wϮ�����,�{������vW��3K���yxv�c?%�l�Kb�R��\��W���)|q9��,q%��[����ĮK��}���n�a���{��_�]�r)�'�z_/)���N�l�b+��(�-6-�Y�b����J�-��ڨ�9��G�}{ΧԖ����t��pJ�e���%���-:�b�G�J�JM����.rџ�ݠ��:IϹ��\�������0̘�hg|BvIIs�����Saw���ʇ���G4�΅�Ϡ ?W?j"�gY"P������Ӑ@�p��ÐB�l�S�t8W pr�����T$u:�Õ��p?����w���&���\]$�b��$�o�^ܙ���kѾ����m6�����u�]o�ٽ�ً\t�Ÿ��[Bnn�;z��͸�λt"Q���N���on���'�<�������OOL�<O�EyUw�g��&�%�f�L������õ�Y�I�?\���u����hY<u���	S�,�;u):/��s�]6
ӛb�r�����
_��G���R�����̰�^����kc��4�ͦs�6Wy��-5�0�\�����6�]^cs[�e�._�CA��o��0RB�zHٿo��>�S?�� O�l٪UH��7�

���Vtx�is8t��4��J4�m�j��m�w��/�(5�_�O!_ega2�J%J��#��X�]<�g�إ{�i�'6�^�٧�Lexb�Y��Z�;�'���|��������Jl��2y�.�-�܌Ȉ��Zu#WD ��x���\���j�ژ��~̯s~Y߿}���E���[_a��p�2�mW|�ҥ�R��(�P�F�s+��(��/��(]�*��2�M��x�k�9��?ós�t�<�t�B�{��#�?=�Og^�{Tx6�k��F��'�����ܙ��r����w��=��M\�C���x�y0e[��|�}������vU��2��pU"R��Ɂ�
��c8�Զ��r���گ�S������r�Jt�ܹ�ug����e�,���o��� ����W;����"�#

�eF���e���سgZ6o�/S�T婌���o�c��-]:�mҬ�ks�u���'`��u���+AD,Щ���T<�$$$����J��ʬWr[�l���kt@�`.�;���*CS���f�^��?�>��t��6��{�Q0a@�2ڷh�ǞxR�����v��V&����a�?�`��A�>������_<��sػG��R���Jn߱ø���vh�] "
F�d�q�&�ݧw�_|�^�ڵ����������:��m;����x�駱j�
������f͚���/s�~y��6�w�� "
6�d)-��p|n���V���]*�J[�j5�nۊݺ�:ҝ���1f��y�l�i80ԫW��O>��/��Lꐄ�cǂ�(1���N�#:&f�
�y*�G��¦;�-Y��������λ����(�	N����h׾ݘO?�$%'�0���:Y�6�6m�ʔ���#���5*�M^n6����\s"��Q����{���K���@��0�=�Q��o��}�'�?�fM��;�"�`ŀN�.��b\{��6�#""|Wf��Ȫ/���K����^�jӎ.�bي�1b$��މ��\�����g��w�;��>�Y'>�G<"�`ƀN^����۴9�����U��Uv[�n����t@�$������ѣ�d�b�	�JtTTr��-�L�655/;DD�:y����`r�ڴi�Ff�*;ͫ��b�e8���Q���㭉1��o`5���W��k�.���� �n��O?"�`ǀN^}�~.����j���s�yyQ��q8�p�"���"*22��g��oLx��ٰ*�׊��ѭG��Np�����޻o���:`@'��M�ݺ�@TT�&e~^nS�v�U+Wb_J
Z4k�`�i75r����`��y���ϛ�����C��޻Љ��`@'��z�\vŕ��Ď�QQ۳27-���m۶bÆ�A�u��~w��b�vs�ݞݰA��+W,[8��G�Գ;n��jU��S߾}p�ק�<{�Z〭�%�:tK�.����`$����˒�����|�)�ߓ���mxi� "�N�ɧ����
���e�Ͷ��뻗�t`ѢE��ɑ�AՎ.'+��'�h7���]ٮ}����-c��� "���ɧ_�͚�D�:�W���g��^�j;iG߻oZ�h�`�״����p���n7���hܴ�����)_}��K�aԨ "�n�ɧ��.B�=l˚ի����Xt��۱~���	��SRS1z��^Ǜ6�,����\�պ�k0�|���K "��Щ\	uиq�ݪ�%=-�M�-����y��y�5�fϓv�I����v��:uz��/�ʱ���)�����b@�ru��I��9�U�a�Q�c�t`������Flt�1oG�v�7&L���[��#���7o�r�/?��y���ؽsN?�tUW�T.w�8�{�^�򚣠� �j�U+Wa�޽hӪ��x�#Gc��vsy6���s�͜�����O��3O���:c@�r͚5]��@|B����������e���ؾ�֭?f��<�`�E���_{�����/���w'OQuǀN�:��q�7�t:��/]�+++�n٭����v��:��(���y�EtL̎�mڌ�����0 ��Qv;"����_�z����/��?x�`�mLӡ�S���BlL�QoG�����7����`n���7i������3#����`ND!���Ҹi�rӍ��:���l��]y�e���ػwڴnu��MB�Ju\�j߻w,�����P��'�<��AC�1۶m��oL Q�`@'�<��Ø��iG_�J�9y+�Ihݹs'�o�p��������`���n��]�v�g�������q��_3�QHa@'�HǸ�I���Y����J,�v�e˖��AgU�9I0�/(��＋iS�I�?����#�7i����[2���ѳ[Q#��ÀN~��q=��t"۵�߅�2�3,�V3��ѳ��sƣ�4�g���k��΄U����s/�`J��]�v�Z<x߽ "
5���m����n94��S��`5��X�z��KA�U3�g��u6�y�w��˪vUX��]��Ν;��釙Y���� "
E����Cҹ�ٳW��av�� ?�2��x�M7VY@��JO�ر�������n�ڢeˑsf��)�a��_����Q(b@'�=8t(>��+ԩS{UDDxFA~^�	f��Ұt�2�y��*9��~�?|���0M'���e6���Mz��W�r�x���0⹧AD���o���Z�i���M��ѻ�23�Xm�׽*�G����ܹxy����̀uU���s���Mxz�3�5�[��ND!���ֿ�?^Ƥ����/������m�5�Wc_J
Z6o��K0߲u+F��m[7���m�ڷ����{�r���_���?Q(c@�
9����1))�s�n+m6���Hޖ�M�6,�K0����K/��彩�-�����4m�t��?��9���дi\q� "
u�T!��ɨ];			K#""rsrr"�n�jG_�l�vj@��0M|��g���>���U��a��~�ĩ���K/3���1�Y��Q���N2��3q�"22r}dT�����&V������%K�������J������k>^�"2��[���ۻ��*�<��?�����n4$kBGMk׭�bv�r�s'k7��f�v�Y�j^Rlk�Uh3#l[��dE!0�&"��*'8��e7��s�[�<|?3g8����w��9���L����ܶ�3� ���~�>*J���k������%��8m�F�Y�Dz򃴘מ���5k��\���G�|}[Ǎ�� ���T�|~�3y��' ���~�6�f��ҥm�3�t��_`�Kjj���ٳ
����Z:;e}F��������zWxDĎ�~����
� ?_�n� �pB��oK�zJ[`ƞp�m%��e����A�%-�-RRR"���;�jQ��y_v��]v�����	:���cGW@@���1��v:��Ç%.>ABCCK||}�m6k�����V)*:!]6�x�}:��W���Xa��MY+��f�����	�����Z�N��M*{��:�m������gŠ7T;v��J{{���_�|%M�&�w����74HRR��*+�^Q���ᆌ=|��W^����አc@�B�d��Sr?ʭ���0�Ӹ��*����	z_h1���ƍ�$���<��
�?w�?����/�k� W29�$��ϲ.%��*�~���p3J�su^ZZ*�Ϝ��s�ݷW�l�"6�U<͛�Un���o�ަ��RXX(��� �pE�1 ?��DG��M�'����X-���q6[�?^$֧�b4��禥�Dq�$'�H���t�����=>�Ճ���; �.\���x�ጠc@���f�~��������k�X:�=]Mk����-�q];��,)�k�d�	����N'QQQ{�WO�?c��v����+ �;��������L1u�
�k/{�$?w��������&[�n�?�#�}��Z!�!E3�e���hjn�m��  A� ����c�>bޙ�uZ���{ڨ���(��e2c�t���ҝ��'37HW�7ڢ�r�K�Z~:yrʮ���t�3R[^..  A� DDE�,0��_�Sl��~�����(/���EEb�Q����{W���%yM����Iϭv7��Fo׍��;�צ~x�;��Ȋ�� �_6w�,���Hxxx�ȑ#-�W�~�o�����XZ��亠����F6��Jj�:���/�Ӽ���ZdT�;�ߙ�>����%9�� �w:L�"uz\����-��dn�����R[S��o����)ٻ����i��%A����3��^{�g5���*� �C�1`�G����>Ѿ^��Ω����t��_� {��S�Iz}O���]��.�X����s����s�bc7�d��ߕ�P�1���y� ��:eF|��
h	)3��6���8m]��۷K��Y2g�,�8wN��$u_�WK/��i���_�Т7W�|�.�,~H  �"���ks��y��t����ߔNj��%=-]���$c}�=rD<=��]�GFF��=gv�ƍ�N����
 �cP^߲E��#gΜ)�;엺�����򤪲J*����Ԗ�u?o8j��֙�fnX���g�!�>yR  �t��%�n�Nʻ�|\z��t~�)�'��MR�e���i�L�]���훶lq���ɯ�<)  �:�d2ɒ����������ں��tz�~���w'L�X}Ͻ��ݺu���ݻD�d;A��tZ��J�:m��/>q����ā��%�GZܽ s�����j��u�̝@t�'��˧G���;�x�iʦ���X�V����`0J\|\ުU�v,8䊈���� �aC��?��{\Ǝ���?���b}�.�K��`4��W�Ǜ��j����pF�1$��^��:f츎�G������q���>��K:�n[xT��i�ؤ���[� �Cf�Ν��ޮm�r�������T����C�i�+��<�����-�  ����2˖,��/���s�J�ط���w���-���*<!!��]wߕ|������� }G�1���ِ������l�X��m�I=��������3>m�^9��ŕ���*/���  ���cH͙3Gv��-oeeɁ��"_�$�ݑ�]�Qn���z�;f�y��g�9��ӈ9 Aǐ[�x��d2���D����t:&8�UN���|�����`4�1��Eǋ���ʤ��V  C��8UZ*:�QBCB�'LL375�X::��lA:�����'wtp��u��wZ,�z�j1M�$ ��!���86ih��^��������dn�:V: `�:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
�O��Ր���    IEND�B`�PK
     `+�[��EM  M  /   images/d3694a2e-5bba-40c3-8069-8db85c4c9209.png�PNG

   IHDR   d   d   p�T  TiCCPICC Profile  x�c``RI,(�aa``��+)
rwR���R`����b
����>@%0|����/��:%5�I�^��b��Ջ�D������d ��S��JS�l����):
Ȟb�C�@�$�XMH�3�}�VH�H�����IBOGbC�n��ₜ�J� c���Ԋ�_PY���Q���Tϼd=#CsP�CT�%���X�}�����ߍ�������k'BLÂ�A�����΂ĢD�33��10|Z����� |�'�8��,������z����j��N��������.j���p  !e�2���   	pHYs  %  %IR$�   xeXIfII*            (           J       R   i�    Z       %     %      �    o  �           a���  �zTXtRaw profile type icc  x��S[n�0��)z^�8~$R��b;^eW�J�ё"�@`H�n-|DI�D��@ȴ�v=L�"�	�s,`�ۮ��z����"H����pz����3�ͬ,9&�h'�tN9#���(���d>CQ�h�|q�k��R�R����mOi�q�6�Z�ܶ=���C�>hrK$>���U`�͚t3�s;����%�S�T�c��\���~�y§b�_"%�G"a=}J�H����|)�Ni����2��yl�c���r�E��|�7$��8��s���.PJ����
��wq�8��P'��j����[ܞ�c2����g�+��|����RM�=�c2gҥl��ϞauTh���҈�\�z���줡㜥   %tEXtdate:create 2020-01-31T21:31:09+00:00��y{   %tEXtdate:modify 2020-01-31T21:31:00+00:00	�   tEXtexif:ExifOffset 90Y�ޛ   tEXtexif:PixelXDimension 1391c�   tEXtexif:PixelYDimension 800�요   (tEXticc:copyright Copyright Apple Inc., 2017���   tEXticc:description Display P3�y��  cIDATx��]	xLW~��d�(%�J"��}�%(�Z���B��_[y~R�R[u�E[[����J����ҿZ��j��B)��'s��;��Ĉ����>���=��s�s��-�37:�PTB��A%DaP	QTB��A%DaP	QTB��A%DaP	QTB��A%DaP	QTB��AW÷&��z\I���7�)I*�Ev�Z�:d;iJ�3mtRɲ�������V�$IY6��"a[�d��$}/����~�l���99��t.��$u0Z��d�M��(��5D��a�}0�*�
��?���h��dY~�`ȫq+��L��yY���@���[���������ƍ����0��`�Aк�C��"�|<B&�������r����t�PQ:�;w'N�{˧����a)y���3�t>���ʂ
E@fB\yyP� �f�3b�1�(p�3!�<ÃY=��䫄(�d���?0��&1A3vH�JIi�	�YCd��c,�p?��0���g�Ж���lqtws���%b�G��ɒ�2d'jaxR�v�Zl߈s��S�����_C���2Js;�i���8�f�ɒM>�Q.]�����С�x�g/�5J<����зO̚=�g����f6.:6lX�t]������B��5�D��;ѽ[7���s�p�0g�,�n�=_x��(���E��~/���u{���F�m�6�2�h��!����v����;����dX�i5�7�}�����ٿ�2~޳?��#n������1p�@xV�$��u˖�Ѳe��H�zi��|��u��,�Ν'�����ԩ3�/�5PP��7o���,�_���C�޽ѵK���ǚ5k�t�:>�,^|q 4�XȺ����7!&&�+{�_�~��d��ǎ	SԥkW�o؀������A��n��B�p2�7n����Na��>$3��ARLN�G��&����~�� �����QQ��wq�������Тe+xU�ºu_ lQ������͐�լ�K�.����ԙK�.��9����(�QN4|���X�p&M|�����5�OLLDu��x�"�.Y�9o��&�l7ww7�b�rD�c�)��?��޽E��jO����[���a�0�?B��ۿr6n����o�Y�}��E�E�:uh@lAZZ*�i`5]�ر�u�9Ǻ��<s�4�V���ի۽��1�Q�n�:AƢ����D�?O�F�g:b����a� i4puuÑ�#������W��u� ̜�iL8^<H�Ȏ��ʕ+Bui������®�v�u�zS����u>l�ФΝ�P�U�@.��+��������^M�5c�L�L��S��nW",�Y��e��'""#�|���'B�B�FMТœ8���	�R��ӓC��w��t�b�_G�R׿ƛG߭~=L�6U��?���קў��ݻ[��Z���\�rLd0�q�	��o@Ey.D<kI��
2^U��~�zB�!C^65V�E�6m�W���$!-^�j� ��溃��������͂�٤������m׮j׮����{��l"��e����G�fg�AQ�%{ΫbM�6��F�흚6m"�.\@�ƍD���]P��	��g�ΕG���e?h�V��\��ӊ�����ٳq"m���`1i.�[8c:fd��Y����<P��6���׻�2�sq�{dDG2kd'j	h�͛��)2;U�jW��%�=z|j���)�b~b����!JcӁ�L��+$3�i��ߪ[�Fc�8����2�F����~~���dG��?��%\�9���ɡ���3lw[wGDD���Ç�6�V�Z8AQ?��6U_"���YԢq�0��$��_M�i������W[P��@�nns+�F*Z��@'����!����ǤI��`�<a�CI�>��p������<*T�[�Cɩ�1K�,>�>}�/�h�M�vhD�*��89�-�aq�֭�M0m�t�jQt������5k?C��M�ۻ�Mk5���Z�e����ZSVY'�����L���������'����F����g(4�Ŷ��P�^G�>|<(��p������_�R�VUDK</`9rr��WhI�6��E^��9��~��΁�ʧ(��K�c��K�^���}Ѭis<���b�s���J�efp �e
���,���5��<�5o۶oD��h���%.�sab��F��%a�ȑ4I܍��u�Ȗ-�!00�==̤?�9@���������A��"���K�T����J��2
�������r�̋h���C�Шn+���\�t	�i~`�'t�dA�����Ӄ|�'���GEDCQ��z�5{zP�gA`�@��?�h����\�h*��5���]�r^^^pbb(��1��[ޒbo�ػ^8�s4�叽|�4�@����4}�#0(h�my
?A�#����Mg�<��7��?�il���_ �2Eto�����"����j�37-N^��4g��)�8����&��'�*JBCLQ�JH�C���=d��,���}X5D�2`�����0��g窆(&Q#,���!�.o���e�TF��[���9ʲIQ�[�<l�M�V��|/="D�xOR���vG�_G�3˚��7��aj�gE��s�6��ˋk�Q'I����܊�GBEiB���j���QCG�h4Z�D�$ݢY�-R��By%�V+i�T���I|3����4����ĉؙ}���2r����)���Om�fk\]�zH�|�R�iO�l�Mۗ�I6_dْϜf4G��Fk-匷�ݥe�k�\𛍶���V���_�3���X:�-�b(ڴ#ݾ���KĤ����h$�v!VI~}��+s�^����xg��p�h4"�E@�Ӈ$^N������1���	�����ǁ=j��������o��qbZW�?��i�1��wI�t�G��v��e��^3�x޹���k+�t�w��`-;q<3��rJ�r�##���Κr$55G��޶;�a�±c_�ٿΜ�V�{J9�Ԕd��=�(B���}�\�.1�7����׭w�^v�.\�[��"{x<����̣������{�"o���]�|ҵ�"#��[v��n�ٻoޚ>�Mۢ�̛;[�A���(Ks�#�����@�V�s��I������׸��������gn�fV��8\��@�*e	%F��#�n�����8v� �2�Ǎƙ3�2+yV{<6���ܜ����#d9�¡��ȏ ""�z�ז-_�M���^nzjJ�QNk��i�܇��#��~_�Z(_��?���&��2�G9��ɡ�=�gge|�yx�fY$�Q�/R~�'������ll���<����� ~�N�z�����t
s�PVQ��<^�q�s��mOrrJ@�=�t-���K		粲24x6�;�;�%JHJJ
*�|D��-KKMN!p5�olI�x��ݺ�Ge�F��kǏ�H�"A�ռ!i\�xzz�/_�<�R�u�7�u�����U�F��K0��N�rx����̬L�(B���^b���x:y9��}���E������k��%u����QTB��A%DaP	QTB��A%DaP	QTB��A%DaP	QTB��A%DaP	QTB����Blg���    IEND�B`�PK 
     `+�[ީ���|  �|                   cirkitFile.jsonPK 
     `+�[                        }  jsons/PK 
     `+�[�rՍ�  �               %}  jsons/user_defined.jsonPK 
     `+�[                        �  images/PK 
     `+�[�:��� �� /             8�  images/c7631ad6-ed21-46e6-964c-e953ba5165ac.pngPK 
     `+�[�AWv�'  �'  /             FN images/97fe1122-b934-4e82-b9ff-450ac31bc7af.pngPK 
     `+�[x^��_� _� /             v images/d5d3b89f-59ab-4c38-95f7-2948dd30f8f5.pngPK 
     `+�[/�i�$  �$  /             �0 images/60da03ea-f7cc-456a-983c-41a209708cd9.pngPK 
     `+�[�c��f  �f  /             �U images/c88b2895-5e8b-4a57-9f9a-b80dd50058b1.pngPK 
     `+�[��EM  M  /             ʼ images/d3694a2e-5bba-40c3-8069-8db85c4c9209.pngPK    
 
   d�   