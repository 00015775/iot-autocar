PK
     ^�[;�9:�  :�     cirkitFile.json{"raven_core_version":15,"hardware_version":0,"pin_to_graph":{"pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_0_0":[],"pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_0":["pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_24"],"pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_0_1":[],"pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_1":["pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_23"],"pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_0_2":[],"pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_2":["pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_27"],"pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_0_3":[],"pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_3":["pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_28"],"pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_0_4":[],"pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_4":["pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_10"],"pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_0_5":[],"pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_5":[],"pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_0_6":[],"pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_6":[],"pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_0_7":[],"pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_7":[],"pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_0_8":[],"pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_8":[],"pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_0_9":[],"pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_9":["pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_11"],"pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_0_10":[],"pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_10":[],"pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_0_11":[],"pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_11":["pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_12"],"pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_0_12":[],"pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_12":[],"pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_0_13":[],"pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_13":[],"pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_0_14":[],"pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_14":["pin-type-component_ac90f49f-b705-4887-b642-1d6309412ac1_0"],"pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_0_15":[],"pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_15":["pin-type-component_ac90f49f-b705-4887-b642-1d6309412ac1_1","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_22"],"pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_0_16":[],"pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_16":["pin-type-component_ac90f49f-b705-4887-b642-1d6309412ac1_3"],"pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_0":[],"pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_1":[],"pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_2":[],"pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_3":[],"pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_4":[],"pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_5":[],"pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_6":[],"pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_7":[],"pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_8":[],"pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_9":[],"pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_10":["pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_4"],"pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_11":["pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_9"],"pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_12":["pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_11"],"pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_13":[],"pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_14":[],"pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_15":[],"pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_16":[],"pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_17":[],"pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_18":[],"pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_19":[],"pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_20":[],"pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_21":[],"pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_22":["pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_15"],"pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_23":["pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_1"],"pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_24":["pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_0"],"pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_25":[],"pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_26":[],"pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_27":["pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_2"],"pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_28":["pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_3"],"pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_29":[],"pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_30":[],"pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_31":[],"pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_32":[],"pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_33":[],"pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_34":[],"pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_35":[],"pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_36":[],"pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_37":[],"pin-type-component_0767d6d7-c92e-4635-8656-1d8c21f3772f_0":[],"pin-type-component_0767d6d7-c92e-4635-8656-1d8c21f3772f_1":[],"pin-type-component_0767d6d7-c92e-4635-8656-1d8c21f3772f_2":[],"pin-type-component_0767d6d7-c92e-4635-8656-1d8c21f3772f_3":[],"pin-type-component_0767d6d7-c92e-4635-8656-1d8c21f3772f_4":[],"pin-type-component_ac90f49f-b705-4887-b642-1d6309412ac1_0":["pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_14"],"pin-type-component_ac90f49f-b705-4887-b642-1d6309412ac1_1":["pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_15"],"pin-type-component_ac90f49f-b705-4887-b642-1d6309412ac1_2":[],"pin-type-component_ac90f49f-b705-4887-b642-1d6309412ac1_3":["pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_16"],"pin-type-component_bf25649e-fc18-4b24-a9f2-ca8f731f26d1_0":[],"pin-type-component_bf25649e-fc18-4b24-a9f2-ca8f731f26d1_1":[],"pin-type-component_98bc3cb9-b170-4d4e-9899-7363cce84e7c_0":[],"pin-type-component_98bc3cb9-b170-4d4e-9899-7363cce84e7c_1":[]},"pin_to_color":{"pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_0_0":"#000000","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_0":"#010067","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_0_1":"#000000","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_1":"#ff2600","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_0_2":"#000000","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_2":"#0061ff","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_0_3":"#000000","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_3":"#77bb41","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_0_4":"#000000","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_4":"#a800ec","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_0_5":"#000000","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_5":"#000000","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_0_6":"#000000","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_6":"#000000","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_0_7":"#000000","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_7":"#000000","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_0_8":"#000000","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_8":"#000000","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_0_9":"#000000","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_9":"#007DB5","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_0_10":"#000000","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_10":"#000000","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_0_11":"#000000","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_11":"#9aa60e","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_0_12":"#000000","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_12":"#000000","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_0_13":"#000000","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_13":"#000000","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_0_14":"#000000","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_14":"#91D0CB","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_0_15":"#000000","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_15":"#95003A","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_0_16":"#000000","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_16":"#6A826C","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_0":"#000000","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_1":"#000000","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_2":"#000000","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_3":"#000000","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_4":"#000000","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_5":"#000000","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_6":"#000000","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_7":"#000000","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_8":"#000000","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_9":"#000000","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_10":"#a800ec","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_11":"#007DB5","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_12":"#9aa60e","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_13":"#000000","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_14":"#000000","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_15":"#000000","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_16":"#000000","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_17":"#000000","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_18":"#000000","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_19":"#000000","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_20":"#000000","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_21":"#000000","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_22":"#95003A","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_23":"#ff2600","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_24":"#010067","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_25":"#000000","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_26":"#000000","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_27":"#0061ff","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_28":"#77bb41","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_29":"#000000","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_30":"#000000","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_31":"#000000","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_32":"#000000","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_33":"#000000","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_34":"#000000","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_35":"#000000","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_36":"#000000","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_37":"#000000","pin-type-component_0767d6d7-c92e-4635-8656-1d8c21f3772f_0":"#000000","pin-type-component_0767d6d7-c92e-4635-8656-1d8c21f3772f_1":"#000000","pin-type-component_0767d6d7-c92e-4635-8656-1d8c21f3772f_2":"#000000","pin-type-component_0767d6d7-c92e-4635-8656-1d8c21f3772f_3":"#000000","pin-type-component_0767d6d7-c92e-4635-8656-1d8c21f3772f_4":"#000000","pin-type-component_ac90f49f-b705-4887-b642-1d6309412ac1_0":"#91D0CB","pin-type-component_ac90f49f-b705-4887-b642-1d6309412ac1_1":"#95003A","pin-type-component_ac90f49f-b705-4887-b642-1d6309412ac1_2":"#000000","pin-type-component_ac90f49f-b705-4887-b642-1d6309412ac1_3":"#6A826C","pin-type-component_bf25649e-fc18-4b24-a9f2-ca8f731f26d1_0":"#000000","pin-type-component_bf25649e-fc18-4b24-a9f2-ca8f731f26d1_1":"#000000","pin-type-component_98bc3cb9-b170-4d4e-9899-7363cce84e7c_0":"#000000","pin-type-component_98bc3cb9-b170-4d4e-9899-7363cce84e7c_1":"#000000"},"pin_to_state":{"pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_0_0":"neutral","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_0":"neutral","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_0_1":"neutral","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_1":"neutral","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_0_2":"neutral","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_2":"neutral","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_0_3":"neutral","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_3":"neutral","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_0_4":"neutral","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_4":"neutral","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_0_5":"neutral","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_5":"neutral","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_0_6":"neutral","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_6":"neutral","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_0_7":"neutral","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_7":"neutral","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_0_8":"neutral","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_8":"neutral","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_0_9":"neutral","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_9":"neutral","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_0_10":"neutral","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_10":"neutral","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_0_11":"neutral","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_11":"neutral","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_0_12":"neutral","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_12":"neutral","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_0_13":"neutral","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_13":"neutral","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_0_14":"neutral","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_14":"neutral","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_0_15":"neutral","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_15":"neutral","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_0_16":"neutral","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_16":"neutral","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_0":"neutral","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_1":"neutral","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_2":"neutral","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_3":"neutral","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_4":"neutral","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_5":"neutral","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_6":"neutral","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_7":"neutral","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_8":"neutral","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_9":"neutral","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_10":"neutral","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_11":"neutral","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_12":"neutral","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_13":"neutral","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_14":"neutral","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_15":"neutral","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_16":"neutral","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_17":"neutral","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_18":"neutral","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_19":"neutral","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_20":"neutral","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_21":"neutral","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_22":"neutral","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_23":"neutral","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_24":"neutral","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_25":"neutral","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_26":"neutral","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_27":"neutral","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_28":"neutral","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_29":"neutral","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_30":"neutral","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_31":"neutral","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_32":"neutral","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_33":"neutral","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_34":"neutral","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_35":"neutral","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_36":"neutral","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_37":"neutral","pin-type-component_0767d6d7-c92e-4635-8656-1d8c21f3772f_0":"neutral","pin-type-component_0767d6d7-c92e-4635-8656-1d8c21f3772f_1":"neutral","pin-type-component_0767d6d7-c92e-4635-8656-1d8c21f3772f_2":"neutral","pin-type-component_0767d6d7-c92e-4635-8656-1d8c21f3772f_3":"neutral","pin-type-component_0767d6d7-c92e-4635-8656-1d8c21f3772f_4":"neutral","pin-type-component_ac90f49f-b705-4887-b642-1d6309412ac1_0":"neutral","pin-type-component_ac90f49f-b705-4887-b642-1d6309412ac1_1":"neutral","pin-type-component_ac90f49f-b705-4887-b642-1d6309412ac1_2":"neutral","pin-type-component_ac90f49f-b705-4887-b642-1d6309412ac1_3":"neutral","pin-type-component_bf25649e-fc18-4b24-a9f2-ca8f731f26d1_0":"neutral","pin-type-component_bf25649e-fc18-4b24-a9f2-ca8f731f26d1_1":"neutral","pin-type-component_98bc3cb9-b170-4d4e-9899-7363cce84e7c_0":"neutral","pin-type-component_98bc3cb9-b170-4d4e-9899-7363cce84e7c_1":"neutral"},"next_color_idx":12,"wires_placed_in_order":[["pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_0","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_24"],["pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_1","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_23"],["pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_2","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_27"],["pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_3","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_28"],["pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_4","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_10"],["pin-type-component_ac90f49f-b705-4887-b642-1d6309412ac1_1","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_22"],["pin-type-component_ac90f49f-b705-4887-b642-1d6309412ac1_1","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_15"],["pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_15","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_22"],["pin-type-component_ac90f49f-b705-4887-b642-1d6309412ac1_0","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_11"],["pin-type-component_ac90f49f-b705-4887-b642-1d6309412ac1_3","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_12"],["pin-type-component_ac90f49f-b705-4887-b642-1d6309412ac1_0","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_14"],["pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_9","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_11"],["pin-type-component_ac90f49f-b705-4887-b642-1d6309412ac1_3","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_16"],["pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_11","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_12"]],"wires_removed_and_placed_in_order":[[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[["pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_0","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_24"]]],[[],[["pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_1","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_23"]]],[[],[["pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_2","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_27"]]],[[],[["pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_3","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_28"]]],[[],[["pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_4","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_10"]]],[[],[["pin-type-component_ac90f49f-b705-4887-b642-1d6309412ac1_1","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_22"]]],[[],[["pin-type-component_ac90f49f-b705-4887-b642-1d6309412ac1_1","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_15"]]],[[["pin-type-component_ac90f49f-b705-4887-b642-1d6309412ac1_1","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_22"]],[]],[[],[["pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_15","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_22"]]],[[],[["pin-type-component_ac90f49f-b705-4887-b642-1d6309412ac1_0","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_11"]]],[[],[["pin-type-component_ac90f49f-b705-4887-b642-1d6309412ac1_3","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_12"]]],[[["pin-type-component_ac90f49f-b705-4887-b642-1d6309412ac1_0","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_11"]],[]],[[],[["pin-type-component_ac90f49f-b705-4887-b642-1d6309412ac1_0","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_14"]]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[["pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_9","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_11"]]],[[["pin-type-component_ac90f49f-b705-4887-b642-1d6309412ac1_3","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_12"]],[]],[[],[["pin-type-component_ac90f49f-b705-4887-b642-1d6309412ac1_3","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_16"]]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[["pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_11","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_12"]]]],"arduino_state":"arduino_off","pin_to_uid":{"pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_0_0":"_","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_0":"0000000000000000","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_0_1":"_","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_1":"0000000000000001","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_0_2":"_","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_2":"0000000000000002","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_0_3":"_","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_3":"0000000000000003","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_0_4":"_","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_4":"0000000000000004","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_0_5":"_","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_5":"_","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_0_6":"_","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_6":"_","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_0_7":"_","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_7":"_","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_0_8":"_","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_8":"_","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_0_9":"_","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_9":"0000000000000008","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_0_10":"_","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_10":"_","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_0_11":"_","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_11":"0000000000000009","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_0_12":"_","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_12":"_","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_0_13":"_","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_13":"_","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_0_14":"_","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_14":"0000000000000006","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_0_15":"_","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_15":"0000000000000005","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_0_16":"_","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_16":"0000000000000007","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_0":"_","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_1":"_","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_2":"_","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_3":"_","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_4":"_","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_5":"_","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_6":"_","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_7":"_","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_8":"_","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_9":"_","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_10":"0000000000000004","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_11":"0000000000000008","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_12":"0000000000000009","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_13":"_","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_14":"_","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_15":"_","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_16":"_","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_17":"_","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_18":"_","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_19":"_","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_20":"_","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_21":"_","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_22":"0000000000000005","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_23":"0000000000000001","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_24":"0000000000000000","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_25":"_","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_26":"_","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_27":"0000000000000002","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_28":"0000000000000003","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_29":"_","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_30":"_","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_31":"_","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_32":"_","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_33":"_","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_34":"_","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_35":"_","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_36":"_","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_37":"_","pin-type-component_0767d6d7-c92e-4635-8656-1d8c21f3772f_0":"_","pin-type-component_0767d6d7-c92e-4635-8656-1d8c21f3772f_1":"_","pin-type-component_0767d6d7-c92e-4635-8656-1d8c21f3772f_2":"_","pin-type-component_0767d6d7-c92e-4635-8656-1d8c21f3772f_3":"_","pin-type-component_0767d6d7-c92e-4635-8656-1d8c21f3772f_4":"_","pin-type-component_ac90f49f-b705-4887-b642-1d6309412ac1_0":"0000000000000006","pin-type-component_ac90f49f-b705-4887-b642-1d6309412ac1_1":"0000000000000005","pin-type-component_ac90f49f-b705-4887-b642-1d6309412ac1_2":"_","pin-type-component_ac90f49f-b705-4887-b642-1d6309412ac1_3":"0000000000000007","pin-type-component_bf25649e-fc18-4b24-a9f2-ca8f731f26d1_0":"_","pin-type-component_bf25649e-fc18-4b24-a9f2-ca8f731f26d1_1":"_","pin-type-component_98bc3cb9-b170-4d4e-9899-7363cce84e7c_0":"_","pin-type-component_98bc3cb9-b170-4d4e-9899-7363cce84e7c_1":"_"},"component_id_to_pins":{"bc8378c5-ac3f-4da3-b662-1e1cdc615429":["0","1","2","3","4","5","6","7","8","9","10","11","12","13","14","15","16","17","18","19","20","21","22","23","24","25","26","27","28","29","30","31","32","33","34","35","36","37"],"0767d6d7-c92e-4635-8656-1d8c21f3772f":["0","1","2","3","4"],"b66c2a17-0752-4593-99ab-d606efa4d77d":[],"ac90f49f-b705-4887-b642-1d6309412ac1":["0","1","2","3"],"bf25649e-fc18-4b24-a9f2-ca8f731f26d1":["0","1"],"98bc3cb9-b170-4d4e-9899-7363cce84e7c":["0","1"]},"uid_to_net":{"_":[],"0000000000000000":["pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_0","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_24"],"0000000000000001":["pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_1","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_23"],"0000000000000002":["pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_2","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_27"],"0000000000000003":["pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_3","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_28"],"0000000000000004":["pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_4","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_10"],"0000000000000005":["pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_15","pin-type-component_ac90f49f-b705-4887-b642-1d6309412ac1_1","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_22"],"0000000000000006":["pin-type-component_ac90f49f-b705-4887-b642-1d6309412ac1_0","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_14"],"0000000000000008":["pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_9","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_11"],"0000000000000007":["pin-type-component_ac90f49f-b705-4887-b642-1d6309412ac1_3","pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_16"],"0000000000000009":["pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_11","pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_12"]},"uid_to_text_label":{"0000000000000000":"Net 0","0000000000000001":"Net 1","0000000000000002":"Net 2","0000000000000003":"Net 3","0000000000000004":"Net 4","0000000000000005":"Net 5","0000000000000006":"Net 6","0000000000000008":"Net 8","0000000000000007":"Net 7","0000000000000009":"Net 9"},"all_breadboard_info_list":["0eae91f8-3d4b-4e59-8923-87a6d2900cd0_17_2_False_1195_280_up"],"breadboard_info_list":["0eae91f8-3d4b-4e59-8923-87a6d2900cd0_17_2_False_1195_280_up"],"componentsData":[{"compProperties":{"mpn":{"version":2,"id":"mpn","label":"mpn","description":"","units":"","type":"string","value":"DEV-13850","displayFormat":"input","showOnComp":false,"isVisibleToUser":false},"manufacturer":{"version":2,"id":"manufacturer","label":"manufacturer","description":"","units":"","type":"string","value":"SparkFun","displayFormat":"input","showOnComp":false,"isVisibleToUser":false}},"position":[800.38168,417.0763505],"typeId":"11b06032-2d2c-49c8-bde9-6a809e00e513","componentVersion":1,"instanceId":"bc8378c5-ac3f-4da3-b662-1e1cdc615429","orientation":"up","circleData":[[992.5,560],[727.8524695000001,274.3795805],[742.8200995,274.41025849999994],[757.8853374999999,274.390736],[772.8585444999999,274.40816599999994],[787.9349379999999,274.3935245],[802.9240585,274.4018915],[817.9511184999999,274.40747],[833.0032510000001,274.41025849999994],[848.046214,274.40747],[863.098444,274.413047],[887.289655,274.398008],[902.318638,274.39422199999996],[917.3476209999999,274.3935245],[932.3259009999999,274.39910299999997],[947.3580549999999,274.40747],[962.3991894999999,274.41025849999994],[977.4525715,274.41025849999994],[992.5043304999999,274.40747],[782.1481239999998,559.9470125],[797.1743185,559.9609565],[812.200513,559.991633],[827.2294975,559.991633],[842.2110700000001,559.980479],[857.2484199999999,560.0055785],[872.2506145,560.0055785],[887.2450329999999,559.9409315],[917.3755105,559.9619135],[932.4044935,559.9776889999999],[947.376694,559.9470125],[962.42128,559.9330685],[977.4518665,560],[993.340342,394.067633],[1008.3944259999998,394.0425335],[993.3375535,409.091039],[1008.400003,409.085462],[993.340342,424.12839049999997],[1008.3721150000001,424.1702225]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[1387.9405150000002,322.5251404999999],"typeId":"69390a6c-c81c-fde0-536a-a1b73720f902","componentVersion":1,"instanceId":"0767d6d7-c92e-4635-8656-1d8c21f3772f","orientation":"right","circleData":[[1292.5,290],[1292.5000060000002,304.8744019999999],[1292.5000060000002,319.7488025],[1292.5,334.62322849999987],[1292.5,349.4976244999998]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[1545.1655875000001,498.05062399999974],"typeId":"81233acd-4774-4b8f-9021-fdc63c90f487","componentVersion":1,"instanceId":"ac90f49f-b705-4887-b642-1d6309412ac1","orientation":"right","circleData":[[1472.5,500],[1445.3065000000001,510.7414999999995],[1458.2334999999998,521.5429999999996],[1470.4074999999998,532.1914999999993]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"Resistance":{"version":2,"id":"Resistance","label":"Resistance","description":"","units":"Ω","type":"decimal","value":"330","displayFormat":"input","showOnComp":true,"isVisibleToUser":true,"name":"Resistance","unit":"Ω","required":true,"validRange":[0,70000]},"Tolerance":{"version":2,"id":"Tolerance","label":"Tolerance","description":"","units":"","type":"string","value":"5%","displayFormat":"dropdown","options":[{"label":"0.25%","value":"0.25%"},{"label":"0.1%","value":"0.1%"},{"label":"0.5%","value":"0.5%"},{"label":"1%","value":"1%"},{"label":"2%","value":"2%"},{"label":"5%","value":"5%"},{"label":"10%","value":"10%"}],"showOnComp":false,"isVisibleToUser":true,"name":"Tolerance","required":true},"Number Of Bands":{"version":2,"id":"Number Of Bands","label":"Number Of Bands","description":"","units":"","type":"string","value":"5","displayFormat":"dropdown","options":[{"label":"4","value":"4"},{"label":"5","value":"5"},{"label":"6","value":"6"}],"showOnComp":false,"isVisibleToUser":true,"name":"Number Of Bands","required":true}},"position":[1307.5,462.5],"typeId":"72c75556-baa3-04e7-55a5-e13f447c8c5a","componentVersion":1,"instanceId":"bf25649e-fc18-4b24-a9f2-ca8f731f26d1","orientation":"left","circleData":[[1307.5,500],[1307.5,425]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"Resistance":{"version":2,"id":"Resistance","label":"Resistance","description":"","units":"Ω","type":"decimal","value":"330","displayFormat":"input","showOnComp":true,"isVisibleToUser":true,"name":"Resistance","unit":"Ω","required":true,"validRange":[0,70000]},"Tolerance":{"version":2,"id":"Tolerance","label":"Tolerance","description":"","units":"","type":"string","value":"5%","displayFormat":"dropdown","options":[{"label":"0.25%","value":"0.25%"},{"label":"0.1%","value":"0.1%"},{"label":"0.5%","value":"0.5%"},{"label":"1%","value":"1%"},{"label":"2%","value":"2%"},{"label":"5%","value":"5%"},{"label":"10%","value":"10%"}],"showOnComp":false,"isVisibleToUser":true,"name":"Tolerance","required":true},"Number Of Bands":{"version":2,"id":"Number Of Bands","label":"Number Of Bands","description":"","units":"","type":"string","value":"5","displayFormat":"dropdown","options":[{"label":"4","value":"4"},{"label":"5","value":"5"},{"label":"6","value":"6"}],"showOnComp":false,"isVisibleToUser":true,"name":"Number Of Bands","required":true}},"position":[1262.5,492.5],"typeId":"72c75556-baa3-04e7-55a5-e13f447c8c5a","componentVersion":1,"instanceId":"98bc3cb9-b170-4d4e-9899-7363cce84e7c","orientation":"left","circleData":[[1262.5,530],[1262.5,455]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"Comment":{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"HW-504 2-Axis joystick:\n    GND - GND\n    5V+ - 5V\n    VRx - A0 (only analog pin)\n    VRy - A1 (only analog pin)\n    SW - digital pin 8\n   \nRGB LED:\n   Long leg to 3.3V\n   1st leg to digital pin 7 (RED)\n   3rs leg leave it alone; not used\n   4th lef to digital pin 6 (BLUE)","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"backgroundColor":{"version":2,"id":"backgroundColor","label":"Background Color","description":"","units":"","type":"string","value":"#d6d6d6","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"backgroundOpacity":{"version":2,"id":"backgroundOpacity","label":"Background Opacity","description":"","units":"","type":"decimal","value":"1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"textColor":{"version":2,"id":"textColor","label":"Text Color","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"fontSize":{"version":2,"id":"fontSize","label":"Font Size","description":"","units":"","type":"integer","value":"12","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"font":{"version":2,"id":"font","label":"Font","description":"","units":"","type":"string","value":"Arial","displayFormat":"input","showOnComp":false,"isVisibleToUser":true}},"position":[1465.495676540669,695.1842731137725],"typeId":"9a5a4baa-44d4-4aa0-8d82-488487322b20","componentVersion":1,"instanceId":"b66c2a17-0752-4593-99ab-d606efa4d77d","orientation":"up","circleData":[],"cirkitStudioVersion":"1.3.3"}],"bounds":{"top":"242.97084","left":"569.23593","width":"1130.49883","height":"548.61343","x":"569.23593","y":"242.97084"},"cachedBreadboardPrettyViewWires":["{\"color\":\"#010067\",\"startPinId\":\"pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_0\",\"endPinId\":\"pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_24\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_0_0\",\"rawEndPinId\":\"pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_24\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1262.5000000000_290.0000000000\\\",\\\"1262.5000000000_260.0000000000\\\",\\\"1097.5000000000_260.0000000000\\\",\\\"1097.5000000000_627.5000000000\\\",\\\"857.2484200000_627.5000000000\\\",\\\"857.2484200000_560.0055785000\\\"]}\"}","{\"color\":\"#ff2600\",\"startPinId\":\"pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_1\",\"endPinId\":\"pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_23\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_1_0\",\"rawEndPinId\":\"pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_23\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1262.5000000000_305.0000000000\\\",\\\"1255.0000000000_305.0000000000\\\",\\\"1255.0000000000_275.0000000000\\\",\\\"1112.5000000000_275.0000000000\\\",\\\"1112.5000000000_642.5000000000\\\",\\\"842.2110700000_642.5000000000\\\",\\\"842.2110700000_559.9804790000\\\"]}\"}","{\"color\":\"#0061ff\",\"startPinId\":\"pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_2\",\"endPinId\":\"pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_27\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_2_0\",\"rawEndPinId\":\"pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_27\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1262.5000000000_320.0000000000\\\",\\\"1240.0000000000_320.0000000000\\\",\\\"1240.0000000000_612.5000000000\\\",\\\"917.3755105000_612.5000000000\\\",\\\"917.3755105000_559.9619135000\\\"]}\"}","{\"color\":\"#77bb41\",\"startPinId\":\"pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_3\",\"endPinId\":\"pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_28\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_3_0\",\"rawEndPinId\":\"pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_28\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1262.5000000000_335.0000000000\\\",\\\"1255.0000000000_335.0000000000\\\",\\\"1255.0000000000_597.5000000000\\\",\\\"932.4044935000_597.5000000000\\\",\\\"932.4044935000_559.9776890000\\\"]}\"}","{\"color\":\"#a800ec\",\"startPinId\":\"pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_4\",\"endPinId\":\"pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_10\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_4_0\",\"rawEndPinId\":\"pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_10\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1262.5000000000_350.0000000000\\\",\\\"1270.0000000000_350.0000000000\\\",\\\"1270.0000000000_410.0000000000\\\",\\\"1517.5000000000_410.0000000000\\\",\\\"1517.5000000000_230.0000000000\\\",\\\"863.0984440000_230.0000000000\\\",\\\"863.0984440000_274.4130470000\\\"]}\"}","{\"color\":\"#95003A\",\"startPinId\":\"pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_15\",\"endPinId\":\"pin-type-component_ac90f49f-b705-4887-b642-1d6309412ac1_1\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_15_4\",\"rawEndPinId\":\"pin-type-component_ac90f49f-b705-4887-b642-1d6309412ac1_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1322.5000000000_515.0000000000\\\",\\\"1406.4032500000_515.0000000000\\\",\\\"1406.4032500000_510.7415000000\\\",\\\"1445.3065000000_510.7415000000\\\"]}\"}","{\"color\":\"#95003A\",\"startPinId\":\"pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_15\",\"endPinId\":\"pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_22\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_15_3\",\"rawEndPinId\":\"pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_22\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1307.5000000000_515.0000000000\\\",\\\"1300.0000000000_515.0000000000\\\",\\\"1300.0000000000_657.5000000000\\\",\\\"827.2294975000_657.5000000000\\\",\\\"827.2294975000_559.9916330000\\\"]}\"}","{\"color\":\"#91D0CB\",\"startPinId\":\"pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_14\",\"endPinId\":\"pin-type-component_ac90f49f-b705-4887-b642-1d6309412ac1_0\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_14_4\",\"rawEndPinId\":\"pin-type-component_ac90f49f-b705-4887-b642-1d6309412ac1_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1322.5000000000_500.0000000000\\\",\\\"1472.5000000000_500.0000000000\\\"]}\"}","{\"color\":\"#007DB5\",\"startPinId\":\"pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_9\",\"endPinId\":\"pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_11\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_9_4\",\"rawEndPinId\":\"pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_11\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1322.5000000000_425.0000000000\\\",\\\"1322.5000000000_432.5000000000\\\",\\\"1525.0000000000_432.5000000000\\\",\\\"1525.0000000000_207.5000000000\\\",\\\"887.2896550000_207.5000000000\\\",\\\"887.2896550000_274.3980080000\\\"]}\"}","{\"color\":\"#6A826C\",\"startPinId\":\"pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_16\",\"endPinId\":\"pin-type-component_ac90f49f-b705-4887-b642-1d6309412ac1_3\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_16_4\",\"rawEndPinId\":\"pin-type-component_ac90f49f-b705-4887-b642-1d6309412ac1_3\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1322.5000000000_530.0000000000\\\",\\\"1322.5000000000_537.5000000000\\\",\\\"1470.4075000000_537.5000000000\\\",\\\"1470.4075000000_532.1915000000\\\"]}\"}","{\"color\":\"#9aa60e\",\"startPinId\":\"pin-type-breadboard_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_11\",\"endPinId\":\"pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_12\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_0eae91f8-3d4b-4e59-8923-87a6d2900cd0_1_11_1\",\"rawEndPinId\":\"pin-type-component_bc8378c5-ac3f-4da3-b662-1e1cdc615429_12\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1277.5000000000_455.0000000000\\\",\\\"1270.0000000000_455.0000000000\\\",\\\"1270.0000000000_417.5000000000\\\",\\\"1408.7500000000_417.5000000000\\\",\\\"1408.7500000000_455.0000000000\\\",\\\"1540.0000000000_455.0000000000\\\",\\\"1540.0000000000_185.0000000000\\\",\\\"902.3186380000_185.0000000000\\\",\\\"902.3186380000_274.3942220000\\\"]}\"}"],"projectDescription":""}PK
     ^�[               jsons/PK
     ^�[B�@\�'  �'     jsons/user_defined.json{"type":"user_defined","version":"0.0.1","subtypes":[{"subtypeName":"Arduino 101","category":["User Defined"],"userDefined":true,"id":"11b06032-2d2c-49c8-bde9-6a809e00e513","subtypeDescription":"","subtypePic":"c7631ad6-ed21-46e6-964c-e953ba5165ac.png","pinInfo":{"numDisplayCols":"29.48610","numDisplayRows":"21.03642","pins":[{"uniquePinIdString":"0","positionMil":"2755.09380,98.99667","isAnchorPin":true,"label":"A5/SCL"},{"uniquePinIdString":"1","positionMil":"990.77693,2003.13280","isAnchorPin":false,"label":"A5/SCL"},{"uniquePinIdString":"2","positionMil":"1090.56113,2002.92828","isAnchorPin":false,"label":"A4/SDA"},{"uniquePinIdString":"3","positionMil":"1190.99605,2003.05843","isAnchorPin":false,"label":"AREF"},{"uniquePinIdString":"4","positionMil":"1290.81743,2002.94223","isAnchorPin":false,"label":"GND"},{"uniquePinIdString":"5","positionMil":"1391.32672,2003.03984","isAnchorPin":false,"label":"D13/SCK"},{"uniquePinIdString":"6","positionMil":"1491.25419,2002.98406","isAnchorPin":false,"label":"D12/MISO"},{"uniquePinIdString":"7","positionMil":"1591.43459,2002.94687","isAnchorPin":false,"label":"D11 PWM/MOSI"},{"uniquePinIdString":"8","positionMil":"1691.78214,2002.92828","isAnchorPin":false,"label":"D10 PWM/SS"},{"uniquePinIdString":"9","positionMil":"1792.06856,2002.94687","isAnchorPin":false,"label":"D9 PWM"},{"uniquePinIdString":"10","positionMil":"1892.41676,2002.90969","isAnchorPin":false,"label":"D8"},{"uniquePinIdString":"11","positionMil":"2053.69150,2003.00995","isAnchorPin":false,"label":"D7"},{"uniquePinIdString":"12","positionMil":"2153.88472,2003.03519","isAnchorPin":false,"label":"D6 PWM"},{"uniquePinIdString":"13","positionMil":"2254.07794,2003.03984","isAnchorPin":false,"label":"D5 PWM"},{"uniquePinIdString":"14","positionMil":"2353.93314,2003.00265","isAnchorPin":false,"label":"D4"},{"uniquePinIdString":"15","positionMil":"2454.14750,2002.94687","isAnchorPin":false,"label":"D3 PWM"},{"uniquePinIdString":"16","positionMil":"2554.42173,2002.92828","isAnchorPin":false,"label":"D2"},{"uniquePinIdString":"17","positionMil":"2654.77761,2002.92828","isAnchorPin":false,"label":"D1/TX"},{"uniquePinIdString":"18","positionMil":"2755.12267,2002.94687","isAnchorPin":false,"label":"D0/RX"},{"uniquePinIdString":"19","positionMil":"1352.74796,99.34992","isAnchorPin":false,"label":"AIN"},{"uniquePinIdString":"20","positionMil":"1452.92259,99.25696","isAnchorPin":false,"label":"ioref"},{"uniquePinIdString":"21","positionMil":"1553.09722,99.05245","isAnchorPin":false,"label":"RESET"},{"uniquePinIdString":"22","positionMil":"1653.29045,99.05245","isAnchorPin":false,"label":"3V3"},{"uniquePinIdString":"23","positionMil":"1753.16760,99.12681","isAnchorPin":false,"label":"5V"},{"uniquePinIdString":"24","positionMil":"1853.41660,98.95948","isAnchorPin":false,"label":"GND"},{"uniquePinIdString":"25","positionMil":"1953.43123,98.95948","isAnchorPin":false,"label":"GND"},{"uniquePinIdString":"26","positionMil":"2053.39402,99.39046","isAnchorPin":false,"label":"VIN"},{"uniquePinIdString":"27","positionMil":"2254.26387,99.25058","isAnchorPin":false,"label":"A0"},{"uniquePinIdString":"28","positionMil":"2354.45709,99.14541","isAnchorPin":false,"label":"A1"},{"uniquePinIdString":"29","positionMil":"2454.27176,99.34992","isAnchorPin":false,"label":"A2"},{"uniquePinIdString":"30","positionMil":"2554.56900,99.44288","isAnchorPin":false,"label":"A3"},{"uniquePinIdString":"31","positionMil":"2654.77291,98.99667","isAnchorPin":false,"label":"A4/SDA"},{"uniquePinIdString":"32","positionMil":"2760.69608,1205.21245","isAnchorPin":false,"label":"ICSP MISO"},{"uniquePinIdString":"33","positionMil":"2861.05664,1205.37978","isAnchorPin":false,"label":"5V"},{"uniquePinIdString":"34","positionMil":"2760.67749,1105.05641","isAnchorPin":false,"label":"ICSP SCK"},{"uniquePinIdString":"35","positionMil":"2861.09382,1105.09359","isAnchorPin":false,"label":"ICSP MOSI"},{"uniquePinIdString":"36","positionMil":"2760.69608,1004.80740","isAnchorPin":false,"label":"RESET"},{"uniquePinIdString":"37","positionMil":"2860.90790,1004.52852","isAnchorPin":false,"label":"GND"}],"pinType":"wired"},"properties":[{"type":"string","name":"mpn","value":"DEV-13850","unit":"","showOnComp":false,"userVisible":false,"required":true},{"type":"string","name":"manufacturer","value":"SparkFun","unit":"","showOnComp":false,"userVisible":false,"required":true}],"iconPic":"97fe1122-b934-4e82-b9ff-450ac31bc7af.png","componentVersion":1,"imageLocation":"local_cache","hasComponentImageSvg":false,"componentImageSvgUrl":""},{"subtypeName":"KY-023 Dual Axis Joystick Module","category":["Input"],"userDefined":true,"id":"69390a6c-c81c-fde0-536a-a1b73720f902","subtypeDescription":"","subtypePic":"d5d3b89f-59ab-4c38-95f7-2948dd30f8f5.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"10.60724","numDisplayRows":"15.77946","pins":[{"uniquePinIdString":"0","positionMil":"313.52773,152.70290","isAnchorPin":true,"label":"GND"},{"uniquePinIdString":"1","positionMil":"412.69041,152.70294","isAnchorPin":false,"label":"+5V"},{"uniquePinIdString":"2","positionMil":"511.85308,152.70294","isAnchorPin":false,"label":"VRx"},{"uniquePinIdString":"3","positionMil":"611.01592,152.70290","isAnchorPin":false,"label":"VRy"},{"uniquePinIdString":"4","positionMil":"710.17856,152.70290","isAnchorPin":false,"label":"SW"}],"pinType":"wired"},"properties":[],"iconPic":"60da03ea-f7cc-456a-983c-41a209708cd9.png","componentVersion":1,"hasComponentImageSvg":false,"componentImageSvgUrl":""},{"subtypeName":"RGB led light","category":["User Defined"],"id":"81233acd-4774-4b8f-9021-fdc63c90f487","componentVersion":1,"userDefined":true,"subtypeDescription":"","subtypePic":"ee130f24-d674-430f-bd58-6b2b8a983a65.png","iconPic":"193bec7f-e59d-4bcf-b15c-6ea8617b7acc.png","hasComponentImageSvg":false,"componentImageSvgUrl":"","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"8.19226","numDisplayRows":"19.27589","pins":[{"uniquePinIdString":"0","positionMil":"422.60884,479.35725","isAnchorPin":true,"label":"RED"},{"uniquePinIdString":"1","positionMil":"494.21884,298.06725","isAnchorPin":false,"label":"Ground"},{"uniquePinIdString":"2","positionMil":"566.22884,384.24725","isAnchorPin":false,"label":"Green"},{"uniquePinIdString":"3","positionMil":"637.21884,465.40725","isAnchorPin":false,"label":"Blue"}],"pinType":"wired"},"properties":[],"propertiesV2":[]},{"subtypeName":"Resistor","category":["Basic"],"id":"72c75556-baa3-04e7-55a5-e13f447c8c5a","subtypeDescription":"","subtypePic":"bbfae99c-8036-4c5e-89fd-a87441410720.png","userDefined":false,"pinInfo":{"pins":[{"uniquePinIdString":"0","startPositionMil":"-120.00000,50.00000","endPositionMil":"-250.00000,50.00000","isAnchorPin":true,"label":"pin1"},{"uniquePinIdString":"1","startPositionMil":"120.00000,50.00000","endPositionMil":"250.00000,50.00000","isAnchorPin":false,"label":"pin2"}],"numDisplayCols":"0","numDisplayRows":"1","pinType":"movable"},"properties":[{"type":"double","name":"Resistance","value":200,"unit":"Ω","showOnComp":true,"required":true,"validRange":[0,70000]},{"type":"dropdown","name":"Tolerance","value":"5%","options":["0.25%","0.1%","0.5%","1%","2%","5%","10%"],"showOnComp":false,"required":true},{"type":"dropdown","name":"Number Of Bands","value":5,"options":[4,5,6],"showOnComp":false,"required":true}],"iconPic":"a262aa33-74c4-460b-b0ad-c746896f6744.png","componentVersion":1,"imageLocation":"local_cache","hasComponentImageSvg":false,"componentImageSvgUrl":""},{"subtypeName":"Resistor","category":["Basic"],"id":"72c75556-baa3-04e7-55a5-e13f447c8c5a","subtypeDescription":"","subtypePic":"bbfae99c-8036-4c5e-89fd-a87441410720.png","userDefined":false,"pinInfo":{"pins":[{"uniquePinIdString":"0","startPositionMil":"-120.00000,50.00000","endPositionMil":"-250.00000,50.00000","isAnchorPin":true,"label":"pin1"},{"uniquePinIdString":"1","startPositionMil":"120.00000,50.00000","endPositionMil":"250.00000,50.00000","isAnchorPin":false,"label":"pin2"}],"numDisplayCols":"0","numDisplayRows":"1","pinType":"movable"},"properties":[{"type":"double","name":"Resistance","value":200,"unit":"Ω","showOnComp":true,"required":true,"validRange":[0,70000]},{"type":"dropdown","name":"Tolerance","value":"5%","options":["0.25%","0.1%","0.5%","1%","2%","5%","10%"],"showOnComp":false,"required":true},{"type":"dropdown","name":"Number Of Bands","value":5,"options":[4,5,6],"showOnComp":false,"required":true}],"iconPic":"a262aa33-74c4-460b-b0ad-c746896f6744.png","componentVersion":1,"imageLocation":"local_cache","hasComponentImageSvg":false,"componentImageSvgUrl":""},{"subtypeName":"Comment V2","category":["User Defined"],"componentClass":"textbox","userDefined":true,"id":"9a5a4baa-44d4-4aa0-8d82-488487322b20","subtypeDescription":"","subtypePic":"c88b2895-5e8b-4a57-9f9a-b80dd50058b1.png","pinInfo":{"numPins":"0","polarity":[],"pinType":"movable"},"properties":[{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"text box (click to edit)","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"backgroundColor","label":"Background Color","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"backgroundOpacity","label":"Background Opacity","description":"","units":"","type":"decimal","value":"1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"textColor","label":"Text Color","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"fontSize","label":"Font Size","description":"","units":"","type":"integer","value":"10","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"font","label":"Font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true}],"iconPic":"d3694a2e-5bba-40c3-8069-8db85c4c9209.png","componentVersion":1,"imageLocation":"local_cache","propertiesV2":[],"hasComponentImageSvg":false,"componentImageSvgUrl":""}]}PK
     ^�[               images/PK
     ^�[�:��� �� /   images/c7631ad6-ed21-46e6-964c-e953ba5165ac.png�PNG

   IHDR  �  .   ���   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  ��IDATx���[Օ��{Ouf4�t{�q�b��`L3�w 		ٰ!��dI�)N6�KB�&�,��lXj�	�L�c6.���i*�ьFS,��+z:�D�F�<������s]@Y��m�uM��$I���K
Aa[6��+���<����{�ߞ\�� � �0��-Q�b��YC�;�+W���*.�%�F�`����@AAAA����z��֕�^ +��"+Hp'K��-������ � �]�O/��AAA�����pۓ%7�zޞ�n�"cHp'���;�en���w�o2A����NAA��H��e�٪o��Y������ ������� [��� � �� � � F�tB�H�{�7��l�3�wb ��63���( � �����	� � �ztX�ϖ_{�Mw]�İ��N�#�Il'� �A�5AAA#G��4�\zí���vcCB�;�K���&�����CA�(R� � � ,�e�3��o[�r�-@
	�g����e�Q �� � �N�AAA��]Q�)����^fpHp'8��߁H%� �B�;AAAB� �U=�l�����9D?Hp' t�(�_AA8M�$�C4��AAaG�cq\�?U��g�[��N z!�� ]�_I:(@X���Z�e�nlV��c��)C�˧��W�U���Žo�t4���$� ���s)&IR$�{�5?$�n �7�%),�J�R�����ݭ�q��X��J�rIh��+A�͐I�&� � B,:,�G�{í����. 8$�8���648�л:v��v�P(ZW�Xе���Y����/$_�z����zHW㉧j �Z{[��C��	�fH���|mri�g��e�O�Q�����X�Q$�a�8^�KN{ǚ���;�l_AEO�������AAQH��!�����+����BG�\����ͭ*�$�sh�~�K-r)q3�!�UT���~�.����Kmon�����z���StM�&���ޑ|�.A��Kj�k@L)��>U�}M�؝z�� vAI�}:ƷC"ڞ���c������G{;�KK^��Ӧ�?
��9q\Շw��A&{� � � l[l��Ï��\y!�\���B撇\y�ʥ3��^ב`{�ᢅ3���+�����]��c��]%�px��i��%�>�K'���dN�~�[��������ݮ���뮮���弸O� � � � �rV0\�x�w^ w]�u�c'A�{S6�౺���DT-yD��8n�1G�G�k�h�㳝�v�ܽ����1��ڪ57���p�2@wwĭi��|��펻�.5�ڊ�h^�Ǵ�~�OS\�.ĥ(zIQQ�
ĬY��P�1�'�$�
� L��=�k�OAA��pFȫ�ײr奰r�)�'�	���j�%)�s�FT-����)�1u�L� �X;(������Z��q+2�//��� ����s���rA[w�=�����Z����k!�$�N�5AAA&�K������\��B�Ip/`$I:�x\���bo���N�mHm�N�:N�2M��q�p��a����6l�����?��~H^m�!qH)�AAA������h�%}	�\�iw$�6c!ω��i)TgS�no��L����¹s'����#�Fy���X�ן�"q^�t'������ۡ+V��v�@�w� � � �D��/�����\y%�\YP�	��R@��^�wFՂj��q�-�w a)�$�(���·�fN ���.�<b�G�p�{�U��ޖv ��kz~�#� � "���K�p9��_/$ѝ�F��9lN{��v�11XD�F,���f��0��J�������ų��5���Ͻ���B8�3��3''� � ��ղpE���
#�%	����ռ=��=B�~ә1�n��DX2i�%��Q��#������W���A8]�S�Z�h�'� � �<G��B7�%�ܢ�S!��$�yMgL��(}�T�=t`��ࡧ�Z� ��bO�b5�^7����������� ���py�b'� � "Ϲ*t�]�-���;]t'���k±8	�w%�0&T�}�p��Q`7�ה���^�x�m�㕵@�LN��2AAA�#�u�����V^���$�yM{D�:L�%K�d	TM�í̲�up�e+���vŭ�<����*����;� � � � rG�겶r�y�ʫ�*��XY�����<��� ��.��=��&�xpɑ��?>*���O��A�ܟ����.aוu=:y�+� �5���t)?����O7EF���
yƦ�����yw߅���ARi�aA��Җܖ�tťk�˒s4م���y��V�L]Q�v�v��ӝx�<�'�qf�|����y����p���Icm�a%��Q �(d$�ƕ�R���*�tx�AVc��<l��h*�G>$�1I���5d�]}Қ�xؘ���l���>|�?U6nD|b���|=.w�\��U���w�	��y������L��w�|���A���m�-@"�nɌ�qM��fk9V��"�Ӌ<�*)��]����^Eq�e�_4�[��.Ev�k�h>�^�lqeG���y��󖂜g�.���'�� ���Ǡ^���t�w�,�0��m`'�'A ��OtI�w�f�e�_n�P�^ � �Ŀ~�y���|%8u��/�ʕ��ZN�{!#Ys��GV�E�#E\˧�j{+�ΛYp�\��z�1�ś����ų�W� y���2sT<q�p��Ǝ�Ewo������A�tt����s AA�5[���"���P�����;/�����C ���k$9_%<�bj��nQ$������RQt��/���q������E�h�KA����{wA�H|��P���s�^��֕�^+��@����̗H,�����+�y./�a�*���)~��&���.>����9]���N	P	� �0�p'� D���K�~fY8�x��^����f$�2�*	�H�$����R�`1T�����<|ng3�=^߶X3�Al�K�AA����Ys�tA�Ÿb��� +�e���y��8K	!�aB�,Q�;!M�D��<�S�å�aLH���v�ѿ�e�km�߻#�n � ��X���HA� �(\���i�u���BƢCSE�k:	�0t�|"�#Y���j�8�8e�xp*A���d���'G���R�� � ��s̹sA������4;,8B�#��0��$�"�(�=Gj�%�s��s��ܩ�Ҧ�Y�����w�MvR�ti|�3�'7e��K2!,O��ޟ�>���C�}.�}ݾd��R�c0�4Mg��z����XlS&e�v x�鷛^���g8[���J�<�_�+'��I��pm<Y.H�z6�ږZ������P����֖�^�2����3��l�}���J�����Pm��LD��-�p�s?2f��M�zD�������|�U���j���Dz�������2���|�ӹ]���$��SΖ�s�$Ґea[���Sǵ�����F�Õ��,;����_��d�yS�����k�s�\�E�w�d@�;�װ�"�c�	[���T�l�`l?>s	|(~r�x��]���uC���3y_WW'�����N�[����`�Lؤ2�A8�v���?u]l��.�&'��`E̜-�CGG;��'�M�gҮR6�6����3uC[��Z{ʡ��E��(�>A�^�����\m	�[{�U�a$h������\�mhmmU��A����C��SLЖp��wA�l3F��T�<JKC��������6��{�b�(;Rی���bq)�Plliifu,!:i�X�'��6�uM$I[�"�mɸ��֝7%k��އ�Z4�i��.��@��~���#��߸ �>QT�c޿���Vq�ݍi��ۂY6h����u\�H��M{oK��F�1����/�D"ݼ�!f�kɶ��PH�#�� b���
ڀ���ChK{{��u�J2>'���hOYYEf"����w��6��䄄0�0��~�1"揭�������+�ܹ����f�w�Lއ�P\4�"1c��4��"�P\.7[�yق>F���&����v;�8Hu�Ij$.|E��^������FӷHH��n�O�؎�->_���	£���`���f��YR�Q���uQ,6�����H�I��%\t7�/N����>�X�eYa�]j�-�k'�}�^�հ677�R.~���:fJ��`���4�"�v�?����7�>'�Xű~�n�8����⛙��@�؎`{A[P�6��1�aY'l1'eS�oC[D�9pN�e�t �:�E��^뮙�`?��+�&lq3[:�,��Ҍ׀�N�@�;a:��CSY'g��p4�$�7�9��X�C!qՒ�Y�lF�Q�N�Q��M�lOD�����]��0s�`�u\P����gf���^� (v���эfaD�Y�~nVC!vF����at�`0j���u����rA[�r�%�AC���m��؏a
�@�;�`u̲���f�LJ�CG_�Ab4X'Pt]'Ѧ!�1�#�wr^��b�3$Y.F��miQMs �ڈ>��}���W.��5��� �� 3H8,�9�
�'3m���([����T[Й�)�F�{&��Nd���㠮"���	D��L`�R��		��"ӎ�2sT�:c�M�m�x�1��K���~d�����!��D��:	N��q�QAF���0A�����u6�l��*�1ށ�u�(11����dL�E	�mID��M�Nr1ot{A[���`��-F�KR �ht�H��IYa�r1FlO��h���Dj��"%���YD �|S<47��O��2��v�)Pt7#`�W�lI��3�\#�%Y�r1VK�9���P����ѻkp���s�D�{�T�:p>+2��`�i����MSS���Cl+ٗ���܉��.-��\x"\t�L��OO@[�9޶�P��I��¥(�VЅ����	�A*8�\�h|����W��Y	�
o("��6~���$�02Z#�0��⤵m1��kT��t0�FU�u �F����0�Ō+\d�J����kdj���มр(J�L!5f�1��0��$�4��8��0���X����<�9A��b塩�n�O���F��8�0�N�·dt�Ѷ�-g�Kb��MbgC��)��;x�&��	��m1bWK:I�(��Qk'��fؒ���8[FX�$���Ip'
�xO#�[W�?w)|���j�x`�P{��]��a���v��B�r!���O��v�	�<�4X8�BQ���=B�
�K.��Pt1Ö�$����*������(P���E����QAmf}���x� ���h��F�^I��c�2j�z:}�F�K��\�I[��LԱ<;~�ژ�� q���W��t7J�E[���M�,<�	�� yX�hPp5����\���5�ɬ�9:y�$��]I,jT��t�bT�1#SpF2͓m?�r��_���/�`Hp'2ƛ��>��ϗ�����;dְE���#
��S�1ڹq��IP�5G�#5�Űh�hx�}��>�s'�<�'[f�;��K���7)%Yf�RfH�ۤ��,RQ���u�ۓ$��dvKFb{.�E�5�C�EG�b;yo&$�	���Ybd�D�^Hx�f�\̵%)�N%�}�Y�)���n�.���+��f	U���ٶ`�8����o�y8f��Jb��>�/�9F#�1H�#9�7cZ*F��6hƮ�T��xD:vr-�`=\��2D��s�UE���yS��n%���<*�:t��l��]�u� t��C���}ے"�' Oi)����x�h(�����i�.1'���ȒL_��p~�F�'9yڸ�wE�F�0�BI��#�I=F~y<n>�3s����(��^��$4M����r�"�}{s��H���GMYU.{��""�\�iQf?�����g��D=N��z=���n̮c����67������h��G���=�l��UUՀ$�C/45��������l�-(P��V���"H�b|j/#ȥ����GQm�P3Ό���+��ZmKWW���v�vr>��$Y67�"I�p�4PEE	�݊�(����2�V͟P���%�\p^i�YDÁ�`uVIii�%�A�ֱ�c���~,++ϭ\$��($��E����u��90���?o�DA&�$�j�~�Ax|�&h�~����D�����Z�U�h[+4|�?�����"P�89ۻ`�ƾq���P5o>T�_ �f���;x���G^WvEw'�HJ<�w:B�Jԫ(��r�$�#������c����S3A�G�{�Qq"�B�Ν� W���أ²	=
���rX'�0y�DKD��ݻ�I�2jT��[�8A�
뗈(���JfO5X.��o�!�Zc�Բ�u)%"l�%��#�G�b��i)X����f.~ǎ���Fc�l��Vڂ�([P,�ҖX,n�r�uwO����*��0a[��`�e��ɓ���ZfKwwD�-S�Nf�ǲ�Sss�0�شiSz�f����FaN�ɓ'��`XA&n�����ءC��\˥bᴶ������\+�h���'2O,R^�*��T#&]p�	���d����q�=�j���`�b���j�k���J�b18�f�{�5hX�]�b.��бo�x�i�����`̉'B���%����23�iy���Z揭�����u5�Vd�\i��.�Pp]��`6�`��eK�:y�_w����n�0���ň��Nj/V!�\�<@�аS�Hv�z�-��q���Ŋ�NID.:ڭ�Et�7�c�E�cԇ�D��U7�ϸ�a��3Ip'2��k��Y�[q|V��a׋/����������y�w<�T̞�>��t:���VDV;q4xƅ*�����[�e}�{��9�DO��Ωh���-ܝ#����rqV��X1Q_� J��A����^8i\s�-����S݇[i�H�ۜ4N��'��I2a9� 6h܉� �ۍ"�b?/� tU�]�?�{��c7�thܰ�?�g΄�����{w*��x�A�{�L�)"����
� zq��6��S����_�/q;L�����C\�X���hsJ{�]'�0tXlA�Z��Hj�DjѶȲ3l��be�8)���{B咿�u��=���l�Șh��sigC+��u7�U:���m��g�Q^E�&ɭ�4~�1l��C�{t1M7�;?Y	��ӿx9?x�i4v���]@� �������[i0�#ݓ�;qG�r�MdJE���	��c�P	���8i!o�nZ���na���:`�A�>'�b��@lJ	Hp�N�-�S��q'��7�9g� �`[G���»<'��xźS8 �o~�~��ܳ}y���}�WC��_�
j�YN��+:��څ̸r�9_FJEq�Q����+2��� 5��Hj���(sR���u�w{�Sz[b��R��Cͱ���
w��b�-"�/e�-�۪S�i]��2N�|��ߋ��y��#��Ș-�N�n��3뷂հy�c"����uw��{v���������D���+A�8#�OKW����	��s&Tt��MnF���>4MLUM�qK}h���] �������+��Iq�贐&�!�_�p�H�sEp
����V�m4Fc�:fB[S�]�Non��({=���M�Y,��:���G��wX��}��}u���n�	��U��4vGI�ʒ"��Jd�$�XՈK)#9**�))el4�Α���9u�Iy�D	"*c�,ll�D�F������]6�! �v�����i-֙�B�#�J���1xl�&������;�=���a��������o�w�w~�#X���C�����(��Y�V�#�� �9���@QY�W�a�&��hP��^�~�*�tK�bY:��.]'�z0tJ!��u�;����ܽ�h�4��Ael.>����C�H`"��7O�	~��h;��y]�w��l���o7�HK���?��7��'C���9#7��t�(�}*�|���)[8�5��E�S&�(ZmE��3� �X�,ѶX�D��A�҇9�bY�J9޻�~��qZ�-�i����)��w]'�4a,�����KZ�G��XI䈞�*�3��?��f���?��� �b�������� 0n�#�x��%���*h���-ґ���þG��;�.�A����G��I��s���r��B ��r��bm��:��H�$�;�\r�^%ꌱ ��}�H��s�m����j'�;2�m��^�b���Z��$�2]G0(iÌd؟�<��Hڰn|r�=�ۓ$E�E?�	���!߈�5���o�;J��P��u�7)���,���	��}P�{��D���:�j,��}�Ha��!�".�%�}+�Ly[B�b��G�z��#�9�C�=V��O"���-4��@r��F��/ZT�{}&� r ���� ̨���c��>������O����NeE>wG�0�ɞC �C4�$�k���������2���X�����!���Z^:o�Ef�loh=�{TY���%�Y-����`�X=�������mE�(am�h�kK����K)v�9;k�8�+w<�ۜ4N�-��hl3nE� �X$��d�x��s������ӻ{��*P�]ql��_P��IG��)c������q���:pUʣNT��u���:��={`��G����J��SIp�:`JU
�K~z��g[�+G�]l���&�V��"�5E�K���eu{���zE�N�0�6�n���[ם#R;'���2�{+�<��Md�=q�8�	�K�AX	��S� ��ՓB�������3�KR�L#�y� 8��>��>�8򅸦�}�n�l��'��BgWs��s84I��*{���頪b"���88e�k�CSE���շ l1������a��"YXǜ�<�I��bR��*��8ř����0�a�d'壷��[b'[�_�1�R�y�.f#�"K�b�T����$�#�m�l��Iy҉��M���j(�<� TΝ%c��\>�� �[�����ťx$������A�HjkED'Ei���I�����rqʶ{��I��D��9[b'[,��c;�V�>��P�;�c��N~r&�N;��Asc0Cp�%�}!$�2�D��4��Ue,���e�~���՞���H���`�]]��}�BB����?�����y�Z�Ȏ�v:�F&��=s�]�����Hpǎ;�8RmM-
�!�nBpw�#�]��w�Ejт;m�9퉭�E��18刓��vځ��g8��;X���8VC�=��-&�Ut%����w"g��"�T����p�w�G=6A��À����!���F�¾�_�ڥK�p&�~(�	Ձ"(T4��=�qG��Cd��%�R��'���]�1"�f������ G��>_���(@��$���#zp��T�Q��۬��vR��H�:�Bc�$�m��vHf���w"g&WW���:X�+�kOF���y3�j���/� ���G�Q����Ɖ`e�.���P���y��1��r'I2L�4���ϛ��:��:�:��׊�Gh/�Q55P2�=����o$m@+���*[�'���>������J��_ds|����������B$2�_��N�1�),�����KKK{�k��5�tM��])��W�"���Z�]�Ux�^������Nڑ�Mɴx<n(.��I���a��Q��ˊJڹX�Kᯥ����(a��.���c�H�2����-y�-�>m��Ta^�u��z=#�%�\<^k�c��ϖ���
����m�3[T�3�V��\�5}<��}u�dߢ���_�Jʘ=X���|�E[��v�X �1��}��_d����w�����$^��m)*�[Z.�@ ���z�@>�ݦڃ������l��\B�`���������^���/�l�؜���w�B!�&lL��DpH���9�_�������PΝ丆���b�ے��,�%����>y���7�!��abl��ڒk3�U�{o	)`�L9���������R����u���;M�=�h��|c]���UPwʩ`gIr��P�y��-�?�nKv �Q�v�1�GC�M�D�}yCsD��?�U4��";o��k�wvAK[�&(�%�-�z�Śr	�0��3�tvvBkk+�My0 ��p��롐X��ј�絏������ֱ��fV�̵��ƌ���ŝ�Q�-�v莘�^�-�bm��pK{tvu���-cGUä:q���h�f�t�xS׈@[ƌ���u�����KGWW���yh*.��T�ı��D4g}h��)LPL�cmu�8��4�\�:6&�v:eB��k�8���jz�1t9g�P�?aK��um�7k�P[:�8�c����q3[�g�5�Y������L��:�m�BKkx�@'�@���`���®�%�eD�ZSR��$��I����狠�����߾|�p��i�s�a��
0��)�6�fX0�}��נ����ؓN��[�\.�p�"9�j��M+��\�ݔ�߰isl$���)�#8�,ASktu�'���\�MI��/F[�w��x�S #�+�ˠ�����ybUQQq]<�ML�VZ�l�DB�˃����\fQ,�(R1��U��Cc3�c��:A܂w��\
�ǂ����Yp[�bmQ*�u}���Z�s���dٛ.E�����]���fQ��I#l�v��z�x��V|KM�A�`s��#
y�ll�oj6M���V�.�ZhKMejl1Ux�6���Hp|�r9��l�񴲬Txt=�RS����ڂsѶ��%�9�M�<��pn�uL�-|� ��[Q�;f9�q=Pn�-^�Uy�Z�,G���1�u����R���0Z����%�)����ph*:��	�If�V�t�U��̲`��/��C�FJ��иaTΛv�#�TP#$�&�����|�1Ph`tkWvb�r,��CB��������DU��,0��~���o�-m��X�ș�A����IpttfU�-��7h�-�����r.�].(�K��m��<Q�̈��7:�� �X��6���l�]-~�q۱����nn���*2�,w�;����Q��g���#��p[�����c����GiglK�%.J��d�p��(碻Ѯ�L�L�s��DͰ�|Fق�mAǢˠCF�h:�>���	؜ӨT6�w�-�o�����Q�p���fF0I9�E1�\�k'�ot��Ta`� e�^�q'W���J�e�"�	"[�l���#$�0���uM����
D�=��dk��%I$�����\�r�B���I$�h���Y��.+1Ȣ��d��-N�αY�=o���r9c4(������(��F�`��Q`H���`P����Hw�:,7��a=��ڳ��l/e:A�`�..���c��r�()T7��rbDX���]���������:*��(t�T�~��@[P���˿�#��2�c�d����/���0�|.Tc�;����--6��$l	A}K+?��(pזi��r1nYbc���s���똱���A�JjIQ�hG��Ω$���Ƶ�E�Pi�x[X����D���q�g¹(��N�炒	��P�;����=*�|����J�����1ϭi��C���}��ԯ[��Np�3�K�)�{Էw�=on�o�0
���~
���t)��E|![0(&�c��`�}���7����f΅�S1zW4|+4+٤Ԃ�@�GU��m��s������F�t�:��R�&7�8ec���$��>d�-!�c���Ŋ&���,x���,�#��� ڂ�̈�,ܙ���9�y�0$Uֱ�PȴrI8�1���s +s��Y
">�Ǵ�����<�h��c������M-��b䮭t��� jD�,�!d���lL�����ؙ!T���,0h�FD���L[�X��g9Q.E&��<$6#ǎ	íK��D�޶=���V�����/H�<Ҷ����k��C�Š���0���`G<
E���-/��=�~kOp7��������j�+㺆9TE�;>�=k��hW��@mn�F��$X�P-�H#s� ����Ao���WQQ��3���8�oo'"&�%dzÅ�|"���
����"��$�]���J��N9�����������nK��������n/(~�m�cAL�6|�law�Q��{��ߵ�
��������]�l5c7]*8%�]�9�ѹSn�-r�y�Q��`ښ
S
Oc��S�%"���3Ԍ�A�$�#@[�
ո�(3�\)�Xkjz&��bv� �]�݂˥<d�.�T�W����w ��+��N�l�;�Rl���ͮ֭�?���XpW(�=G�:��Ͻ�:�p:�}�=��<2QJ�3�1�N���Ol$��: ���?Y��k:?�S�D�"K�89�v,����Q6���ك[}1�zDЄ'�n���?�����s�ʆ��e�-�KL��2ء��+��ae�v�!&h\a��x���{O�色��Q���PQ�F�>�u��
ݿ�$������~���Q����gڥ���Ol��E=y�_jK�3�;�p<����6v���i�bs����a{��Q�(��g�J��f��>@���H[D�e(�s�����z��}��3Nkܩ����o�$v��u%��0��2q��gJ{���M-bw?D9��灒����>��Z��2"����˱����C�A��)�2H��=�s�ّjK��1��&�@�Z@2���/����`�Ĳ9cH��@�w:���B�M�8�#*�\N/�[k��m�����ظ6\�7Ep�(�;AX
��]-�������d/�h�hCb%)ٯ�tS�����pтip��Q�T>�����#����d4���2�3��6�/}�e4�I��O�5�	~r�`&��?\��]�ђCJ6,���_�Bc$��:���Uv ���!+�@��#)|;.SE8+�Mk{'������-��bU]ôa���_6�L,+�+��X����>l����V�<�s���`��IVق~fbK6�@��T��%۹��c������Э�����lɴ�XU6����X���NGtیm���2蓇b�9�PL�U�Sw��I1/qZ�n��@"���y� ����)��p�r�/�+������Dw,_��Y��p���x�΀��D��@|M>���9����z��r��ƝT.���?�m����LJFC;�A�'��|�Aw��5���L�9j_f�QN�|g�D�D��e�28��'O�����
o|�b�1MR0��,	����~�͖��[��6�ZƖ�f�����.[N���_�Mr۽���y?y � "$���A���c�g�q�p'
�1}���p݉G�/�{~��~��t�X��ajUY�k[5Ê�=͝��oH�O�Ȁ�@Nx�.��8�����6����pͲ�~��:��;�|���Pu#� �@�.�bn[n&� �M1^p�"܉�����ӎ�����~<w�d��I;oju����p�=O	�	$s�nΐ��F ���!�#.Eɯ=ry�����	��yS �yr�6f��B���<y�'� ��H���CSU��j�C]	� ��Du��:V�Hp'
���p�){O܏���?}q�؞dŬ	�h�hxg�~ѷ�g�0�f��I��<W918�6�e�Ip�s������v�> _yj�6��gA��T���R� � �B���e�WEx$� ��.�wP�@)e��ٓ�	���	�������3�;����9ue���ӌ���]�C`b����(�d(�m�tFȲD����_�����W���gO�|��5�_~Y�9��&�� � ÉxIp'� ���!th*QH�]��ŧ��nPd	�l����O���b�t������sP�$˝����u����X{;ؑ�w�ژ���W������p�I!���~�]���������gG���e�S���.�Q��QUK$]g�׊$M3!y �Hd�$)��>�3��i��˒�zX�j�ʪZ
6ۇ$ɝ:޿��J���g��X{q��b�C�	�Td��-"�qP\]ɗ�x�i^�ڊ�ݾ܏��A������ZZ�x�@j�?W4�x��wE8ǋp�H4�4Yf�d7.��=�����D��N$��t�\.v�.P����~J�Ȁ���O2�������>1`�ras���<䞟�#�+V&�(��,�����-��+���<��w,'f���>K��q��["���C�x$�~��C��\_�`��՛�v��a6�������ǵS�ޙx�
�"�X��Ñ�"܉¤��������a�Ժ�~ϛ����o/<���1!c�7��bYUU �5b��7�"�gv�@0�O��&l�o�__�����+�Z��^�U[vr�nieGQh��ob�����{�&�:�� �q�M:�]Q��&G.5�J�(責+�eQ���n��&�^P\Ŭ3/c`�@.�(�y��;Aךe]C<ީG#Q)ՠ�]�;�\P%��6�T=.��.K�������&�9_[s�u]�� ^�M���:�N�d˃Ƈ�������1ţxb�8Q��.M��ĺQϑp���QY�x�rit�ף�]If+E.ao	�w��\6+A�}@+�ԍW�Y���c�������:�Z�$I�cJ_���s]XN���RO�I�{��%�^b���I�!��"�n�\n?k?Iq{v�yRH93Eof�ڢkZX��:!�q[�a:�3Z=�W��$lq�G3�5.�/)���Ud����+��=K��t<j�BYV�(�C���ڊ���"p�J$I��_�q���8*��̎f��ì�v��%.G�l�a�M$�V%��{6wd����-"��e�H�pt�-�$E�%^�Ou`�������&�p�8��߹h��?�w|��U�M�GI<�"�p��<�8���H:k\�ˍ�Y�U�%t�}�	�K��������d}*�F��B����uHά�{�
yd~�4L�d;h���^��3v���ј2+Q �;C�QJ�pX���tEq��'�Q$��l�+�=b���"6]L���63[��G��[T"����?���zH3�w���I"�v_��B���;+�b��1�2�r���2��Ⱥ�
�ݷGu�R���(\��O|X;��g����[�rA[JV��˹�zR?�3+��H�����^g�,{D�'�sl{*+?I�z�S���{��sA�~!�~{�O��\�Y�y�xO�|t��:��X���=/iq�&T9!���y��}�p1Q�E�D}J���������'5�}kv��=�Вƕ�|�,K�
��T��wH�����H��_���c}][	v���M[͝�u+�ޒ�-3O�l�m��)Z�G6�i]�>=+Z-{�l�J���P%��z���
��Sc��1@��h�ҷ'T��<cϞ�V�z�7�M�3��~�}ztSH�j��QͭiAI�GR�z�'� �\��1�����Rj����J-[�5��]��H�q/["��u}��xq]��T�+�g�.8��*mrѴX�l�6D�0Ķ���}Ek�I�"�^���F�Z`9��t����]���}�Vf�5҈�+���G6�`�3��݂�m����
4K�ЊQ�Ey��#�*�c�����8��#Z�Y��5h��A9�EE��0[Bܖ..��JR��p�J�-n?�E7A{t�r� /�ܜ_�+�q�I�l|8�C�\mJ�4�O)�w@P���s .)e���J<X�g5_G�Skc����0����m�­�{��?��s��:"��K�B���g[D�p'
�ww��_]Z��rH�Gڻ��y���@&U�ezi�6&��u�Q�v���pQ��Ƨ���;�^:n>�(�A���Mm�ӧ߂G�m�x����.y�+����Dr�b�}z��M,U6mUp�'`�б��$G5���d�F"��D$w�<t	���L�y�RV4�_�.�3�=/��]��}��x�O�Ep��^S0����&}��)�����2D$���1�=Qy"{�D0v���J��枠|�T�>>cm���n��in��%�wD��O�1ܙ��Z\�c�%Ee�'�{ʺde[� �p ���r@	��
�6�l���f���PU�7Tt��MMO�/Z��
llQ�����ʈ��cm�(0:%/t��E??�FX�	^{����]�L0���ĈN�y�"�K��]7t�\���K�J���R��"V�\(,�Z�?��a7�C�y*��
�=��*�S�T�{M�z�磇�-��-l�EZ4a�؂w�Y��F"��5&���=�p;z~W%s�K��`���k�0[$<��LD����z�jOw�Gt���Gˎ���km��&W�?��*R#�c�ڡ'�l9%�^�?��=.ɽ":
�	q�q�n��a���2�Y+��H��j��!��,K���\����#�9�2��!]˓܉�ye�nh���"TWaʈ��{��c@�l;��/����6C�K���v"�cQ<^{:%$�w�s �\�><��f���G�����}���g��o^|�Gދ<��6�&�cڨ%����W�l!X�	�Y��)"��[�*l�4)�I<3F��L�N#AɫJ��ݺ�l8��3(ʠH��0
F[%?�;QpATvA�?(���E}��q���X�C��I��T(�K%�k]܉����O��=mр�|��yl�������'���c?�,K��C�$J82\E6�t�!� t7���㕵�����e�̂��؅:�q����m�����mA��� AA�?��Nd�m/���gM��c�{_�o{��>N�=�e<JB�~ՠ]�b��T���٬�A���	���5[U��S�����gϾg1	Ν;N�9A�᪸���G�����`{c+�H�  � � �BA�4�y	�F�fӋ�iw='N3kʡ���ڰ����D�*���+�cg����}�@�$[)���+/���z ⯪;��F{[���G�Cf֨
XPW��anm�����y����`ws�?6쫇���w�n{e�""34 �p'� � �BA��D�y�_ظ�?�}�m�#�m�{�_YE��UW�a�:�;t��}͇{����{]�$�
AU����[Lk��zkW�;�� �yˁ � � �B!�nHp'�;�BM��O�H`��#���C������ � �$;�AAA�.�}@$	�D�����J˦N���^b �	������:A}�Nt����QAAD!���N�5�S�{�0����1&W�P�1�-4m:qC`��#��N�� �8c<�m�&����`z��������aNm%\���=_�CsW7��}7l:� ;�[��R �����JX2~ԅJ�|�$��NA� 0�d{$]y>�EYѩ1"�>�2}<<���g&Ua���?�|�i�P��܉����3�kK������a_|����u��
�^~:�a��
��Ν7�|��O�7�7�^�}�6T܋G�O  �p�>�g�
�~�h�:z� ����D�j���'agc+�Ձ"8yz��1�M�� �&����|�R���- ���p.����YC�nj'�ʶ���W߂�����,�.8e���)��҉�r�<	���UÁ�N���>��ƄJ����l��;���5��\�(�3:�ǎ{=p�����o���v ;1kt,�Xs�T�C��1@w�ԇ;� {|���o}��ϩ#q�ױrVo&U������v��M������s&C�����~H�k4k�G�r��5X�ytD�y����c���[a3�� �OU]�`[=j�(���+ۺ#���I�-a󞫖΃G�l�=͇_w�H�>/�!�Z�!��9��W_��_��ęO6ĥ�p�:xc��A�ǥ�헟�U�?����i�q,�n<�������.��5{2|�ԣ�Y6g�[ZӱlM�l�X8��f�*�����z16om��!6��x��^ۺ��y�С�D^��:6�c�6b| o���Y��?���'������D{Re�M�y����\�Sp�PǅGQZ�4*����u��#�0�"��D�W�/����z�.���0�G�/�1�]1�=�ق�޷�=Cc��J��g�����ކ;^x�����b��y'������|�lgP ���'��u�d���l�����9�^v#ݤK�����<�?x�u��O�-��#/�7n:�h.�"-lqr�C/�S���_^
'N��Ж�fX��-�,�6��|�l9Ԝ��{m�~vች����ǶܧՔ�]������C��9k�$�Ŀz��}vcrM\�p&�0mL�.�=؆�l��X_����݆;��am�'-�����ᣯ@G�}�Hq�����z��F�~��'^��3(tn8�(�ފE\�yp�&x�����a'K:����;.f���??�����O��/>�ב���[_Zw���-"��Y������ˎ�+��;��m��WW?;9~T�k��xq�s����OM���k���}��˯_x�V�+J��/�G���w?�?|�%8���O���MK'���՟�۟}��̱���糹���J��`Ֆ�����ö��N:�8l�o�|�9��wp屳�Xm�~~���X�"�qB�RiŬ	�gw\��z�C��3o�?�D��~�	�L�)e��!1�DOF�#(����$�θ�+���A �;{Q����|�^���$6Tuؕ����N%=�;2gl5�U	�4��Pd	�f���N���N�Q��þ�Ͽgy�h���.6c�����������������HlO���~�?���S�`��}_9�G."w}������aOK�L����u�"J !�����_��'�o;��/�[
�3�_����5����"n:��#)��y�#?��A���o]̣˲�[/:	���ӧ��pղ�p��E�}V�i�*�泏��-�?j5��}D��/:�WlGN�5���������p��)�g.�Y*���?�n��YX�q'2%1U�`*|��}_���~s��� �_>v6\��M��gܗM��?~�A,l�?auf7=�
���S&�����q��ˀ9�rV����3��!��Ue���O�Y���K�98��tጌ�{+�)U}�~7�vwr~���"�݊�]v:ۑc&��G��<����lN��W��E�T�N��k�?����8e�8��/��wp&��������ހg?�>�op^����{�38>/�:�9�;8���7/�9�UY���ջkO<�;��p��A�)s����^�d��4��+/=�d������'V����Ta��qMs��S?Э��-R�Y�1}�7�Hk��i0���s�S*(���Ip'
L�ʒ�cm#���iupp��	PV�L�t��G�YMzP���n[�������ߪ�/�Qt�p�t8nBd�bϛAA3=b�o~��<e�q��>g�?I��LSg7X�.]�S���B<B\�`|��������:�x����v����<k�=��O:
^ټ{Ш[�Y2e,��i��өí_8�x���յ`5c�K�ۧ/��x�n��?] [5��1�C�=������rD��H-�-E0���.�r�>����`3O3dg��ط����<恶��h�/�]:d�h���>�խ������zJ
���`	�4c<<���B���/_1@lO�['�v�g>�� |֒���s��o��p����ڔ9�,?�9�ll��%�3&��Y;X��}�q|��묝ע�{ߕgZ������z6ܿf#���U��-a��d�:�qn���DK��<@�k[��Q��ccs�b{*�͜ _?n.��u{8u��=�J�����s��h��?ض��2�?�*)��6�f�Ԧx3��I6=�#��,;>{�	  �N�Gt�PD5J)C���bUE����y��6�=m�8(Isd��g޲E�n�7�p�T$��Y�:cI�ƍ���̄#j���ok^ܲ��ɀ��o��.���h��3&�o(�'��o��.9r����LlO��Q�?vb-��ث�eҞ��Z���F�c�d*�TPdx{��3��}�n�ue�0kLSv�b=���m!�_���M0�#�x���8�O�w���O��7-��'^���^|=]l�42;Z`��J�#��ק͞_g�S�
dy���F�Uw
�<k	O��_o�t��H�i���d*�œj{S�%������~����,����)c��;��[>w
:S���y�m����������sfi�k�/�O���ϭ����{��'�{0N�3�������X.�����u� _8j&�c��M�=	�{*(���~Ĥ~��e㶕�;���d�H���<�&���9����������ݥ�w)���z��%�R����R�����#���+��$dBy�ʀ��9����3��n[�b�g��g�-����(|�Pu�`g�q�ڙA�Lz���c����/.瑄������Eo[W7LU9@<yc�>x�{n�O�%)�B�_���0"��K΁sfM��+΅��X���QX�g_�뫶��g��J��SǤ~�z�C���?[���?�߼�����:�������`N�2�0��EG���r�����]��O�3	~~��Y��g�ft��ъ�: ���4|V�<��`ځs�O�_]��W[>s<�Z,<ج�����	ѱxza5|�m'w)Μ4.8i	�8�l�%~�ܓ���ӎ�7�>V�畜2k"�k��{�AsS3x�^�:u2�I啍;��ǝ�<m��g&�9x�j�
�n;1�(�n~l����a�F��[�����Y���ys�ҽ����_�ѻF��/�ɣz�V��0�6g�^��,��9�0-��R_cc�6vϩ�;�����۴ߺ�jgFyg���6�ϐ8����GG}��]0#EIs����\�Ǿ�-+�j�j�&ZwM,"
?L���5�E���mi��N�7<�sGN�ߢs<�Z�S�?yLoj@d����C/�G��ީ��޿�x6|g�Q����yc��*%X�a���K�t�Rx������@��[lPpǃ%RN�Y�ɒ}�=�A��8���*(dƟ~���݈���]�0�ⴈ�6��X���ހC=ۃg���ˎ�s�?���x��2���l�cfÁ���`z��`��QC�BY��ꋰ�w����ġ_������Y�*�g��mu�+���*7�2��"���j��k����	��Ϋ���m�x��w]�s�c>��R��&��篽�G��G�� �N)��΃9�_�G��S����w������P�T]����vN�0eZ�X�i:�bJM����{�G[w��8�G�]�4�R��/��G�ON9Xu��jfKlo�F��ZS�+|577��W_��77{}��	��wD��c֎�养��ȋ�ܷ/�����hP�M��Ir��}͗�O�A����3��������s������oW��9)�/Mq���{{�vdӁ&.�?���{_þ�J�ݝ���>*��P(�ޙ�(���êM;M�w4'��;��u���o�?����iu���7^�t���/q粕�������������<�L:x���}��|���b�e��0oL���yܡ�iUN�>�;�S�!���o^���q6��?s��](F���c�\��VFMO���'V+�#��y/��'�>�wGɄ�R��wbD̬�]r1<����+/��o�@�A��b�5[+�Ͽ ���F�F�{��`ܩ��E�EIZJ�pľ}��)�8�����жv׃m��O)�>hI6��΂�Ȫ�;�؞M��'�%���l���kC](K�Jឺ@�:���	?{�->o� m��"KRl��I]8��+���,(T`^��7��<�����L�?\���~(�09��w����-0��z'�RJ�}������'���a5���6wڎ�-��xρ4}�}|��ז���x��Z������--J4���`osZ���������Mm�<B�Jp�:WO�F��m/���x_��=�~����~c�_�<���AR�a�w�z��I^ݲ{��v5�W>����߉$���-+�)�~v��;�l��_|�?�d�7!M�3��}��������9�� ܁���x@/������E�����y �x����/���6�����i�<��~����}�zRlG�J�;Cdɺq�4�~��gնD���0%�䅽�q���5������Y\���g�wD��V�=i6���ѱa_���Z����%�g� ��Ș����#�t�ֲ|����;V���v�WW��3΄���}�y��v2�	qM/�U��`�ѕ0F��~�s�;�`	�}<�R�"D�����;1PPOO)yCw<�o����ç`I��S���������5{�] }oM��	�|���, G�D�aʕ�);&�Y}K�f�Z �g������̝|��/�_���l���ň��<� �[;Ep�z����4���͙��_�_�:�u}�csƄ:�{�����}y��l�|�������o0�B!���olKy�L�YV޿�M�*�Z��k��6:T�z�t���d+�~&��IP|��������p����|��c��bj���(�Z�dǨt�jO����m{���x��#i��������	WZNf��?�8}��ｅ͕�}>����cL��mt�,��~�锣�_N>������惉s�{hͮ0*�_(�]ivۑ�ÑD?�j������)N�_=�z�؎T��P��:R�Od��*.\'A;1�ރk7��/X�w�!(���oGQ��Ow�GL��ZV����?S�|��L����?�fϳ6�	d�s���G�i����n{�E�}�_�H��g�,ࣸ�6��n6�F��$X�ݥ-P(������ʽ��:mo�)JE��[p����7�Iv���Mv6�Svd73;�3�<�}��r)���%$��������2��U���f�Y>�R��
��3 ׳�����<-�P��Gw�c+v�N��S���qt��a�ՙ�c���6���*�Z05Z]�%�pOOu��\p��V&�D&3[[�l����^�wV��8��Mرh6���f�Y�3LK,���e	Ƨ� %%���N$f`�����=�11R��)�}��DܫV�+������Z�:�¼Tk����=��Њ�pB*�wG{���,��?b.`��D��q�½lPxEcLd�@F�\�,�F\��c"���`L�^p�����q���Ȱ��[���i�� ��$Ꮎ]T�<-'��  ��P$���;�N����R�����A3����o���R2���O�&Lγ���H���Rp׶e!�~�뱋Xs#�k��a��h�=�\+�}48���Q�� w,���A�!���8�lg������9�hY+m����UgY�p?�t>Nc=7�l��ٖ��(���ێb�٫�|�h��g���7Rm�'������w���5`Y�&\�����/,��MJ�>�d��VlA?�3��\�vO=E�	�7�؊�,{䓻F�)#������#����	τ��j��V��ya#��V��������7�j���5�oks#]c��!�Y�ͩ�,�I��0!���1�s{,�;�k�K��ﾭ���E�����Ÿ[���6���\�N�	n�RD=��%�Dq8-��v{��S��bJ�0���$�{:;�}��N���waڷ둘WK��N��>.�0��йr�ן	doc٦ZEu�uA����lCDg�L�E磠�t��ƌw/$����Y�1S+:����ހO܉��X�A��׹T��Q1�7�f��Dq#Y������Մm�����#q�µQ��b�r����F�C��o�9�����sqx���ﶡ�3�[8����bTT�r�=��V�=��4��X�7���{�]3t_ҫ��q4��rf�뚂���2[�Jʰ��uL�/�����&C�Ĳ'��S�Nqn�Y��I�/RE��O3|�.E��D�$dS1Ry�8\+#�%G/`��O#;�����^g;�3�����M�t)7-��Y#���u�dS=��&,�ڼ��-y�O�j5��ܨ�x{�fsG��Y��)���f��,�6�������;�r�,|�K3C�E��IX2��F�;V�6��fcPV	�+���/���&�H����u����d�M΄4��U��V��W�n����v���.MY�4ҫ~ �
Ծ4�!j�7���:���
���sn.�s��Jfk�4��)��1��PQ��i��h���={p;>c&\;��Z�5���T� ��:��8�&jO��Ԩ0��Ԥ�"Y����tL�f=Ro�� �Y6��\Mp'�$߀h����}
+L�f�5�*�wo�Hd�I������V�Xy�k�n$�X�1�t�I�<a �/i�u�_X�q��xw�0U�Z�:�����S��k���A����;�C�lR�X�(�Ż��	���¨MA�����^��&u���Z��>��|�+���q)v�>Gn>��!�:��-�S����\p'v��$��&>���G�ocv��|�kD�N����lƒ�'�������}�46F�HL_s��r�̨�1��=����'.cߵx:ٳ�3ch�]�g���~>��&cH��N~�fۉl���v-ҵl\�4����<6�iI��tC����j���۲�|CЀ��`�c3T�d�"�"joP=����TYr4iRG���J8�2E-j$R�A�|�-*��>�jXz��xKx��~t�N�(��V�P���}��(��QH�B�k.�s��*��J_�Z���;�{?�/]FI���Gs��5w��c=x6!��6��[�e6�6��3{��TPW��d���1���z(���V���k-EQ��R�-����-G�5�Y�_X�7X���f�YX�C"�>�s�����5���2K���q,
��Z~�_�2>*̧׸�1���v!3��@k���ps��z6�D�e�����,ۂo�j0�x�A�: e��x,>�;��yz/�����"q�߶��������XǄ�y�D���&<W�����)Do��?c.���ۙSIu�)T849�4�������W�Ok�İ$T�c����ͳ������@�T�[�G���%8����-e����S}Qo�&p�Ϡ���=Q���������� ��+����'.�'�'����<w���[�!]�h��)���D�Wk@Y}O������=}�|F��������g����gi~8tV���d����2�3$�� =������1Q�=W�D���s5
ϵo��Ҝ{�'��R0-�8���pn��*d-���#���QU"�(s`��1KkB���9�����5�g]�W:�:���5��(�fHX &F�bB��LdWghx ���e1�a)(��ZQ�[��M��ܛ�n�G<�>�~��:��r >_�=��?�AC�A"��%���黚�pWg��k�t��SD�N�~,�i��o"��7����Tt��bޥi��8#�вz�?:�'+f�T�A���m;�m�}NL�N���/W��	1�k��Ϝ��i��a�I�t]�}o�����ܒ
���3n������=S�'g�P�v�ӿmA��f���]����������G��v��f��<pB�Z$��W%t?����G/`R�06��-���*k(�]����c7����x��-�ޙ�̺"�98(��/v�E=c��+N�����R��~��}B�j�W�{�+�vbh��l�u�8�ug�pQطE�� �ݸ�%�C2��LtO-��A�)�a�٥���]'�ӽ�MY�J�~t*i^�8�e}�!�g�?
����9(��n��w�U#�$$
+�S8��s�����Em�8:�����}^xv��6��Ҷu28��B��c�h���)�}5�M/�"�=1�kFwF�P?&l=<(ʢ�;	T�|�mJo�ݣ�AGo���$d�p*��Bw$0��V�MLP�؄/W�x�6���i���*��X����ט����I��pNE�R�N��;ݝ�����h���������\�=!V��
���ۘ缿����0��Ƭ�
��$&�Gygl��ˍ�|���8��e�ޫI�r1m�����e6�.����F(Sm�����BT�7��X��tcdo'��M���Il\���3�2�=�58Ux��ի��wϲZ0����5����.�����<�r'��v�(�@7g��ۢ���~P�7��8y�_�ʇ�DH$
����wN�����~���Y��bJ6�d���z9;`l�06һN��ܭ �X���g׮���c����PԊ#R�V��ڢ�?��KH���'��X)��yl�l�i&l�Ǩ���^�O�F_�9�N��}Z����=+M���戵q�7�$&�k�^�/�"�AS!���,�D�rZ�������i�p,	X�๱�8��2�9pb�2[���4�Y��%��[�oB9��\p����}�HL���.G�i���ߧ��JF��Dv���p�n��
�<��F��S��:;gÆAjc�s_i��������<#��Zq����C����Il�mG�p8kg�ն�|��P1Y�p8�@~���=���|jΧY߾����1�'�+��.��?(�M��E�ssf"���Y�i���ZXmo�o� �w�믠���<u�NN�Fƽ��R�L�Yn�w��C�e��ɶ�*����ʤ�8��6z��c�
��Ԩ0���(8��������]�a�P�fj;]o��;�erwaY�$���Q��0w��O��0�[|1gf��Kk����`�v���4�g����"XWmN����N�)*ĕ��N~����p
0�3^���R�c�Pu�/��i��t�	�޳��;p ����e����na�5}��!X�8*&=%t��:u��]��5p����J��1�4�;v���]R�����W��g�N��v�jn>ʅ�/�S`3��\c^.���V���\��X?\�l���*T�N&��I�*D\�pz�p|;o<{��U�}���(tŃS���]Xef�ֆjFl_4�3�����J��N����Оg�FR^!��� +|ɱ<4@���ss�=?o����#>�k+.�d�].z��;�v�
%{i
��e(*�@�w�E2?�~W3r[d�m��E���~�/F����lׯ?��Jm�8ډ�g��4��T��L��.!�,2�#Q&4�^�8�	'3�]�l�Ч};���4fMf*v4�k(�^�T�'�mé$qxy��������8t5Yc���������\\�~n��B�����ƣ��"&>�%��HX�"V�M�XP�����t�89�,�K,s��eR�{���:0;/��cK��Z���|�:��±P��G�a�P��K�=�
�R��ߎ]d�Ь�o�apq�������u�����v�ߓaӅ��Q��6��i����捇��-~:|��ɤLVX���'�xx:ϭ���ki�d�go{OW,�o2��ˏ_�rP����f�sB��`
�
���ker�0�sub��Upop��c4](U��R��?Vnǥ�|}�dD���}�Bh�-�S
o���/���7��&��Z��6"�آ⨝���Ж�r�����΃����N���Q_d�{��б�9?m��,tW?q�I�Cj ��.���F�A��HL��<4�7�1y{���9�H�S����5��y;0"��-��L{OX�]±�y�0�=��?��lYƅ	��q�������#�sB�5_G6���Ú����8��q�	�@�������ݬ3O7Ϗ�Ƣ?w�ñvh��ZV:��ćw�`6}�O_�5B�Ս�������Fb���Ξ�]�|�:�֓=�ޟ9�͋)��v��6�zd:��+��?���߬���X#���l��k)�7�1o�H÷�>��I���[��a��9��i���=u�o>Ԣ5�
Xw�W�\�Ns��7:��ũ����C������mO{9�r�j�?7�o�ޛ^/�㺆b@�?�Y8����Y���AQ��̟���GJ~,��c�ٮA������Ι�T������8_YY	��
�T��H����Q8���%�co�s��ۿG0�}
����x�,��[٩?�$R��͆�\ԑJ��X��y0	ؒ���;Y��̞���}(���p8����iL|�{��G��ߵ�����1����Ij��Kǲ�>}�	�-�tno�;���V>4��$ц�I����_V���
�V�&#�e��h��U�=t�4<�r�+��FA��'.�����j�����Gt���>@��]�_�����ɻ����{��mw;��W�8�[$���nΪy�@J3VgJT������R%�ո�S�J�:"B�⌠���F�-G &�#�;�y�پ�VEf�)z�kWUe]y	�r��$8�r��8��\OF��"��Ҫ*쿑���B���R&G��LE"q[��b��.	�J��Xܵ2G$�>/�j��\K�'f`��k��o&E�y�Tr&8k���4,� �0�Һ��F�X(j_8ן�~r
����u��{+C�:K�a���subV3$�g�*Y��m$n)c9���1�z���V!t�l0Pw�	��b���۽�0&��r�~!��m��ۊZ�u�� ���~�x��m[��c;*��[u���>����##���N�����)κ;��X����YƲD�i=u-GN���{�a��T��@7G<3$ue��J&t�`q�]�R�A`��**.�j6ł|�5櫫�wy�e�:w��d�64 ���#H/.�>H��h�p<ѯG����5f��n��gh��2�L~+݃Ll��P�--�w��b�J�EtmH���O���롱N͔��cHǠf��ө!��
�vv��1X5���wN� �]�9MEG�S4v�(��jO��,-{^L�5�����L`��(��Ve�ѳ���N�z�U�����5�]!���P�p��c4v�7�A��Mg}ay�*v|T��#�pc*&�A-=t��%ÜH�6����#l�Lt�:��c��s'�\���<ީ����=��p�`#���ɤ5��+����r2��1E<��]i)zj	�_��n>�z�I-(ſ6���t��wl�-�(�:�%����til]�5o12-K���5�k�{=m!�/�*��'���v���� 2��G��8c鬉1@b��Qͳ`RG�n�v^Xd�c���n/t���B{/W<m��b!�CÃT�8��Ĝ>�5�%�������aWU��z��Mpg��̒6�&6>�c$�BS�WZ�]�1�����B��(�)8����a��k��:M�dgc��KQ�t���ok���i�؂���NIi��������z7uTnv�&y�T���˪����k۸஄"��bSEArΜF��Sȋ�EUɭ�89���3��EG��K�6D�l�v���í|�p͗�e���jӽ8I��U��ߋ5��)��,��$WK��a�E�]L��b�ԝ(���=����^l�DWg�e�nF�:��.�Q�nZ���jN�)Fv��3k��	qp&=�6���D�"��/�/�7{�a���9���c�e��KK���,$�"����D��<�����#urK,��pn�nW����F�lO�*S��^����E�֘�}^r�yi-^��R��Wb��1�cC��L*œ+��Z1��R�?,�o�/٨7�5�L�NE��;�+���'3�u�u�
��Rb����ā/g��y1-w	�E5����9F�p�)h[��3A���>��㓽a��,*:��;77��&�,'E7Q�����BT�R��J����EUi	�\�������>�p���s@ \��a�µab�=#�m�@��\*����Vxl�C?�U5�����Ns.5�5�(e���u���3��@F�Ƈi�d�ϲ4ʴg0xa�q��<�:r/�ꡊr�quU�� W��j��.��C�u
rJ%R&�UJ,?�WV��<��O����p&���=�h�Ӳai.
��l��$4�Aؽ�i��[��M���^��9R̵L���Ԉ��K��{4Dҽ�bz8kgX��%ԁ�XkP8E��H�Nlz.8���-������Kk0/�+^�0P5Os����w[����n��M�����P�7c8^\�����e�]��Sg�G_I|s�a�m�}B�TO�h��>l�A	Ygݻds���.���HL���E�}���h	�
˫��ۇM����4��*�K%��>�p���TdIY܋��q�ݧK�<z=7�
�vd].4����'�������$�^�F��x:-7�*`,B�tj.�����6�Z�%���h�ɱ�xu�n�su�X��V7�Y#�b�̱��E�U@��r�DQ3?���WwBN�n+E�SD���z�����iF���N)���C�vj��R�{|v>�PZ������Rr��Wַ�2ˆsq:�{VQ)J+΍����7������Yu�.75��²
U�:�ʤM�i��S�I�S�C8���cS��X#]�4k��|�
E�ɦ����,p,K{O�vj�﹚N�2�S0>�=Z��l��܀k�:
��2y}��C��i+���{tH$�ዽ�`	(�l�c��Y��+���,�h��K��
��Q2�h��Q�xc�`�|��"���z��^����J�;��;�hV9���Y�*u�_m+���J(��yYe5�Kʅx)=�h��CMm�m/�s�CEe������X��9���]a__&�pbd6$*R������o�t�97aI�S���� ��{P)tB�J+�+L���`yuJ�gL�p\eUu�՟Kr�e�Z�Ϟާ.�d�W�h3;�J.�3�C�����$)Jm�Qlc��qS���c~Y������rwTg�5f��\�kL��J*�^YS[Yݵr�F:��zM����m��U͋@�fHIy������3K0��nO��Q����	�VlTQ��3XgeǑ:|�?Z�<U��q+�������le��E�F��ޚ4X��W�?k��l�h�G�z$ �TV�c-{4�[�`3�:[+$쪳�\�Ŭ08�_c��+I�:�aB[���&�����R��o[Z�����<�w�f|5w,f���}$��rfv�'K@V|w~��������������W_/��8%ꭣ�B������?jk����H/д)�q��8�"^�@ě��R�P��GTSS�R�Y����uY������n=���ѻ�x�HDm(��?����V?6��zC����h�+3������1�w���C��n���PXQ�Wl'(3b��+lj;[v~:i�	KABCj~�J�6V�U��$�"v�e�5K�R��g�G��o��9����HM�����xdH6��p?kJl'�ӥ	�Iڂ{�{��7������H�
����tm��-�~*9�y�[+����݁��X��������̲��������vK�^h�*�V�Q�ƣ˷1�)�I��q���ߟB[�2�dC4��X��L� �/�M��/V!.��F���>���)PA�H�	�ل����g�u��α~$
�Td�X5U����p�Jk���Q�H�Z��.�5ձ���I"���0$��nP�[���C\��7©9�t�ғ���"��B��3����>�>���}"q��]'���ql^"�c�P/�S��:��PP�9"�Cav?�P�QSP�¢�w�W�#L�L���M�I����5SV�0v!ͺ���]Hϱx&#��b�A|z&��N�@�o�e��K��c��X�g��G,=v��c�9};c��S0��,�<�����mŲSX`�|x��$U��#K�t\��t��Y[� ���u~��$\p��!�*�tN$f�pWX֬�Ӗ���jy~�f1�҄Z� ��E��w;aoc��t�����޲I\��=�a*�N~o�a�9u�uJJ**aEj�c�2�}-�oG/�Jf.|�5,���P\
K_�:cR��ԇR���2?[cPF���!�WS�/1���e$� ���.F[8�t�Y���!zKu�m�kǚ��#wֿ�n�kF�g7/�
�	�-N�C�EY��DP�8C�K[�"���z�Q�*�j��Ƃ������l�ڒ���{��羾{S�½ݱ���,*UmC���;��}������ڃ-��Ӳp��vFb�����g.�r̃�iw�c�P��='Y���{aJT�������eu5ʘ�Ei�)*Ѭ�R�6~�'����LzOEU�^��l�F��Sp�t0=!�<�����l6�E(w���(����-E�'j�5�����"������k��䗜YX�����|T�#9-MVa	6��k�{�:���L��b��}�Y�5�=�s������78%�>��ā�5�ST�ڐϳ�I�)`��=]Y����`l��e�A��ə��������ٍ�h'*�2�J�lSc��<q�ݫޙ6��	d�Jf��������=�R�4��	�9VOmm-I9fA���*!��YV��pnJ~a�^6��8���+(y�$E�xo��2��%�ESI�p���B6��������)�ˍ�\P�rq�f$]���e2�"q�.��-�zEjJ'���
��U$�G������������ o칚��9�����Q��ـ�� �`�|��>�=���c₻8�t�IfGB���2^��g��i�X��w�Nxvt_6�0�.�����9p�ց��F�*��{�s̆Տ�r8�d���Ϛ��iY��>;�����T,&�N+�g��A������ .�s�/�ߏ�g����"��Zp_~<s��`P� ���q��b��ԭ���cyʪ�wq)�-���d��tӻ��ێ���'�i=���iu�4(��]r̂D®'p8GH�R>��j��ߪ]���E��78��o���Z,��G��!��y?od�2�c0�w��S���"���Y]�|�ؓܮ�4|�9Vj�F�����������ю��.\p�X;��w�Y�Ie�C�w�cV��G�7K����EM��An�Eak�u��*�
���z�I�X<e8���ښ=xdpp8m��i���r)j/<��^ȸ1����������傻X�kj�w��Ȑ���Tp,GFa���u+θ�A�ǖo�����"�B浍��i}��αn
�~��T¯'��"�J����1���0��vϏ�Ǌ��� 9�ol:��g�Altj�y}�ࣝ���(ұ<7&�";��͙��φ�,EWL��K���ѐ�JCPgwٱXV�V��y�?4(
�F�a��r,���=�q$1�{Dg��o~á�-%��3ƛ�w�^R��3$��p�8��Ql+�6P\jEo3�(��΂��Yu��F�u[\�M�K7cÓw���4��� ��Ta�Y�\p�:
��l��'ȫ�q̆�F�K�s��ߝ>!��x�-XwV��`�@�xp*ݝU����t�D������O뉷�e��;bt���e�ֱ�y�aق)xa�^�,�cy}��ߨ>:�)���)�������ˬ�Q���dpw,ه((�K�܆���IV�����mj�h�MHl�������p�2
n��*PpE��#�����)x�Z�~I�2U�vǡ�T���)�3�]+�#�e��&뙸웸�����;Ǫ�E��N��Nn[�ʘ��=0E�rS3�=��k�	OG{���{ޟ9�3p.5�fjT8ޛ1����E��ӡ�X<�±������D������ƾ�6恁�XØ<�i���$����C�U�A[�L�v�����9(����\n�ߗH����p8�ù5�/f���x�q�l`j��{�A��#�}\�P�8a �l���o��N�TӁ�:�x ��i��αj$�p��c6l�r_��*(R��;Fh����	�v62,_0E��Nޑ$��H�xm� ���oX:�7�V�S:�z�4	�K��Wl/�š�X(���`i֓�c���>�����	!�����yE߱>j��'�˫�y��Τ�/���p8�����R���hļ|?����w��ké���$п0�:��d�>�vb�.�>}���>��E�＜ؤ��� �6y0����e1�V]�B�p��c	��V[[���QTYUU�%�e6R8H$R��N���Dg�pq;��i%���#أ��%���j�/O�H/��Q��q�X00�͏�ܞY���4��li��0�%ڍ��G�FT����� �����z�_�:��+�y�$�O������9?n��� <2����!ʫk��`i��h~��F%ߛ8
7�o�fy��/��`�5�y7U��7�Lܛ�>�c8�v!�����p8�a^�p��������}�aݙk�p{�������!̖SIVQ)�;pb�Y$��%�^�C2��$��}����f]����xu� ��|JJ*���֣�\p�:7�+�;/^c�Ϻ�{P��Q��ᘃ���%䗄�᣺��i��t��PF����҄D��VlS��EI�ի���,E7M1]]p'[����y��˶bz���{w�;l@��:���V5O6?��3������v�xa���?�f,݂�I��4՚��c�w�w����S	�ͱ�i��N�k��ù]Xs�^���1Llz��O��òg���=;���X����צƠ�@��1˙���XX.��~�?;���.!l:���Ow�`��/O�l;��"���F�X�Q+�z�.�s�G��es�9m���2�B/9�l�針Z��(,�z�8��&�a����Wc�z�%p��<�r5������o�y�1��~��n˻��oM�#���2�&�����~'�y�fk�u<���,GMp_g'���Z��Y�%���i�|y��IiR)7q�p8��ᘇw6At�t`�d��`pw�;��A������3W!6(Hg�7k�hD�2q 䲺���v��4E��t�<8-�9V�����G�8�@��n�Uպ�ñ"�K�5�S�ؿ��9>�����i�l�	��]�3���,IqE�Ƽ2�}N��,RC���|�I���Q�XB=-{,�Ʈ�4-H���ضp�jYM��<�w�hx�[�^��eUU,�G҄N����ENI�j�����_"1]oW����p8G<��o[�빹�uih���i[迲`pSP�3�Ot�F:��?A�.��6�g{N��-�J�5��;Ǫ��Iy��c*kj����α*b34�Z�
J���A���jD~ڏ���e���ய�jk��N��n����a:�R��S+w����^�Xl-ۼ��)�D��QLi�40B����j2�����
߯��<��Z��̞��+�m�[�7b��4���^�B*����p8��1�ť����!�����{�"&� յ��^c�;ه���8��9V����9桰�� ��q&%Kh0���ف�����`A�gW�f1%.v��,�Ix659±x�I��L����ζ��?�k���y7���L�j�dw��ģCz����lmd,Z�m/���	YAU���:�%�8�ޫ�,"�R8�m���>�`oC�|텫��%���c"B����1!�&�^��-W�Y��:����o��oN�{c�~�TV�(&�߀5SP^��Һl��c����e�8�'48Wc ����V'���=+��A�0�II���
S���Z&ͅ�w�>.����[ӆaHx`�۽9m(��
q0.b����=>���'��ĥ�\�q�2D����k�Zɱj�2poW�Y�-�,�ceP���#��������%G/`��8�eNZQ��r`I�X~����u�b�S~��k�x�Ѷ�9a�b���e��:PB��!~z�E��#���$����gc���0.I�ڷGO���w��,A�����_�=���XF���j ��2k���1�c(��j������b�鋍nCY�	{}�����{��[��%X~�"6^����Y�+սF������09⮨�x}�f��ck�`��+���Xƿ��ǿ��m0����瓍nSQ]�w��R�鼹�ٲ�G��`�1F�-��������]±b��Ϩ��Tj���ẗ́z�!����|1�S8F��7����ُH)(T���8#���?�~Z��)��:����磪�&3�lڅ>�~�}�tt��4�3\O��k	������v͝z�AX�%�p8c�)�����JhO(�j��A}�����߭c֜b$��k��Wl'�Q�,f��f�8�����%pZ.�s����.9f!�����X%��=�y��L<������Y�U�t�
}���6|,�����:��#�)��*�6����r��JHL��;1���(�4=�"��3vH���DҼ�����+�Y�Y!_�O-(�ѤT�<S�F<�c(^3�:�7�9�Fd��7^����²�Kt�!|��X��D䌢b6M��������@7u(#�V?SI�f���QXQ���VUi�8�����bt�����l�y�,���i˕|��(�<=���Q��Cw`����3�T�n&
��s�Z��N��g�� A�K�������5qײ��V��z�����p8⇂?>�k�F��K����;�����#���a=Y����:K��	���sĕOY�K�?W'�2���|>�u�Yv.���V	�t���jL�&>;K�R�����αj������(�c��TT��6`��w��X�PCj��UH�PC�ѶAp�|1��$��WTbΏ��D��,�߯�5)��E-��cp����R3ڠT�X^p'�fǣ�0����*6޲���+��D��q��ژ�R���v��n�����Q�ӆ�[E����7w�Zl�S���o�����!_��`̵�.�p�>u�7]�ǽ���#n��1g���:L��.��{�O4�D׮1�����
�hՑP���;��U�Y� �<�����i���}���p8�3�o�x����,�p.�l>��B����7�O����ذ^Lp�(��ǔ/W���d.���uY��L[}�*>�sW�jc}w�,~���cCz��Q}ر����s�b�Gˍ
��R�ñ,Rp�D�y�-���ñRb�s1t��xy� L��,J�Ǉ~ۊ�b��I%���J������X _�a±<?&��c�r�Gb^!X����ڸ�YtPd�K����x8��;�R$�;1�} �?��߸����*Z������w'�Dd���X!Q"�������/�����{c"�mj��N�;fܵv׼�{�̬�����6�
�[�ˊ����1U�5����׮���v����=#U��==t>�g]��5�
���Kx�U�ݧ�5rk�����2���F�|��A���j|r �ñN�ދ=/�>���E\V����ۛc������јۯ+�C�0'�V�����7�/ˆ]�
�R�Id��ٞ����y<>�'��� 7g�6y0^X��������Ϋ�q�*Jv+�,W�!Ѡ��g�
�P����Ϧ���o�e��17�!��������Q'Gl����	�͝�7��g/���$V,�</۹8���/&w������*J�<K�?�	o}o�H<5��

����`��=�:o�:���"�K���un*jj��_�c�A~�Ay��I_/�sͅ+����F@��;�ͅ⽖���������;��~nOw�l�@�J��^T�z�:!n,�Y8�ri]���\�+A�}d�l'��1�G[�}R�_ɬ����TP�&G;v����8�����Ƴ-�^��2�lS74�!��������wV��w�pJL�#k��rv�����د)�{y�lC6Bڂ�v��;�G��dG����5(*k�o�����Z���¾�z�<��Cgݏ1g�V�;���p8���L���p�N�Mɂ1$�ᅿ��������^x|XO�y�(����bYL,��w�������<��N��G��`���g���
�RM����n��;綁�/7�*� q�����jW�2,]败!���=-�T*S����<("��({D���z�ek�'!Qg[�
��`>�6^c�_�����A�~�<�����g�}Ԩ}��e�^�����ofNdQ��P�A|n>��N+,�+88i��Ϝ��Jl�zCg�ѧ������:}l�f$��
�	/>���ư��n�	|�E%t��^M`Ec9�v�c'�u��cOޏ?���tMу��k�Ա��)WՆ���5��OĻ�aN�����%Ȫ4�Y��ͯ�;��ߗm������%(��c��|`���p�ORn!f}��Y��E�����,A?�pB��e�Q������X����{�s8�PRRZRPXXP\\Z^RZ���;9:������f���:I$�}uj���U�{�յ5�EEL��$7WW��L&���8;ɤ2����+�7+���1q8뇄`S��%�����7��1�]6R�G)E�oZ0�Z���:�/=y�O�!ȵ[���Jv��r/G�<k�^1��0:�x��T�o����[�N��]���?�8��|m�U.��"ڙ%v2���Zu�Lt��'묋�9���n�{Q����殃�߯���C�F ����m�Z����fT��w�Ⱦ>r
��Z�D��'�[�X�����X�,��p8-�9lIxoKPfcR�H��wǲXk�29%5y��݉{�DZz�GiY��B����Z/4�D")������]\�J���B��l;m�$7G�a��<�[�fE�����������Ds8� ��㺄bbd\H��;[��vE"m�z�2���5����5���Ug�Ͳr����:����:��+t���&�R��!+��jr5�7u>#�EA�3 8c"Bu��c���w�~�>v6��^��W$��),ohw�;س�%�WW�W���/!�M��W0b� �:�@��n������{�� [~YC4�{{����=�� z�/̫3�S�]M�1�M��ث���vv����]�ѭ��eչ�Xq��Ȥ�p8N��n� Ϻn���\$�p�]p��o��6 oyrLBh�V��'��cg�.�6DV�J%����ń�I�u&UͪeA�
���+�k gX��%E?/]q���������(,
��"�n�{UuM()-EFF6N�>�V~-�<�����]j��KF7���R/[{g����\�a#�� �Xl\�˪kTҢ�}X�I[���?vb���p8��"��S��c�0�j�P^�yE2�
�V2k���O�A��_�6GSZEpߗ��w��Ȏ-��G��̹P4#�i��k:�F���¾�P1���I��9��#��aSѱ�ib�cF׎:��v"YXi�j�2���-.EmW_A��/.6RvGQ.U���%煶��z��{���b��X$��Tm;�ow
�Ф�N64O�ߊc��{q�nV�x~�(<>�7T��=X�~�\I�[ㆃ��p8�����70���j�q|�F�Z�=\����!�i7r�?.���!�f����"�X�T��y����\p�� ���rL�Glml#������-vJ������l������n�W�j���mk҂�J��`EU��յ�f�����J
*�����LϨ,-�����R�PZrDQZZ�(+��-+U(*ʥ��	*�m�P[YaGA䨮���o�ښ�?_QK&V���	=�j� թ�E��nH/��iWb���ld�^���v2i��ܦ�A���FR�bk[e+���P(���WU�0e�R8g%¹S��/�T��eU��U�
��[���r���^&�t��X�M��w�Ihq\C
1Ef�:q �9�����������O7�Ě]Wq;#�5/½N�3�]a�HdR�p��{lv6Z���Wh�l%z�����l)�ِxݜ�u����Q�!�tG;g'dk�Z{�J�����\�]O²S�����oMK�TfAw=Q��^������S����q�oWg߅X�ׇ��j]\���ښ(��l�R�p��&�g,]�Z�Ɂ<>����n+�]�#5��{�nܡWlW���W��Ż{aAt<38ZU��>�w��9Ȋ��箨.�p8N�)�j�uu0)FT�P���'�D�g�CnG_�����ELb:�<u�/$`l�&�Gx����t�E"�2�ۋ�G&�����H���2����������ǳ��`8�A��᎖è�}�*O),k��j�����^:�j��V��p� 	:�!~u"{TB�&��m�+�TZ�^���p9�^����(��YT�wy������[�`�;��h�I��XF��2�}@� f#��:a���Z�;km.ef�ǣ'��nh�X�F~[7�syZ�\���/�_cE�����ܥs����I����
��5���W���V��1=2CB�p�F
�'��I?��QC��@���&�4���s�����rPq_��ᜒ-ҝݺ��#'� �dr�p��p8��c/o�psK������~b�:�L�ϦO����rfĊ����k�~~�_�n2E��T�]9�P(B*++��r����55�b��q��9��mu1=��H`�D�)Qah�j\i��b���nw��nb��$;OVŕ-_d*�L��� 7��~5;��bx��j8�K�����ֈ�Ӡ��H,eH<�~���Hj�r��sJJq�F2F�Y^�6�~e!��� q�25b�rX1���\�����ͤ��v��=��s{t����5�U��o��ݍ�5���_a2*��_�����ǡߗKT���b���������5&�S�������)�����x��l@���g��0QqVuhww^��&u��^<u�ڲ48�8�5�Pd��C��t�X�YX�Ҫjt�j� f���F��5����z8�Π��vZ�����B;�2���u�1/���><MC˾�#L9�i�eR��I";>�01����g����-A-z�)��X�zGu<[!2��@Q��
��V���W���Y���B�鏀RG*m�wS×�_�c'�&���>�M����T�������N~�]0Ζ�|̿�>^g9YʨC�u��{�tz�8tBc��g0g���?�zO��ߴ��������a��Ѿc:�^�<���zt��`	�3�1($O�Yݻh�}}�0�:z�.��kt��^�d�4t�����pn5��[�ޝ5Jg�Ҋ*�^�_��v>g�2!z�­������[c��)���&�~�>ŧ")����[�p��"�;:(D�﨩�m���p.5C�����ƨ��ؾx�	p8��t��Ċ�\O�'3rY25���q��Y��%� �fF��*�W���˽�w���#Z7{�����N��TK��
�r#�˖j��\S"��+p���C��3�
�����I%:�.�ᳩc���Z��ct��{K�G��;����3a�:�"��f�r����S�"��+�ƪ�o:��ǎ�'�ߵ��3�(�櫪��2zw�ILcYJ���s��k�1$��䢇�'����R�ӝQ�ٔ"\��O_��ث8����κ�x�������pnu�vW'UUcI�-���-��j싽�Ub;��B����c,���G;��{O���n)ù��ADFmm�9f'��on>�&�c}�	�'����n��I�����ŻO�Z�M����`{>�u\Y9�S{�|x�>���G�oCa����ۍ�f��*��4���w]��>��4sA�r9�xV��d�u��"��r#��z��@��t9^oT��;����řy��w��=$��dQ����6�&��k�T�?�N���.oj߽������g��םl��q��*j��;���������l�Jirs����P&�8��CT8�L��*�X�t?���l<�jV���VΛ{[vC�C4d)C�}G�/S����FbSvI).e�=����p8��V�JD6@�Υ!��T��@���T�}��xn��C�pK�Uc|��I�ȓI�7W��\�����p8�6I� lzr��G��+����?o�i-��"��d����6��&�PB*Fvf�Ѣ�}��֣��!����oNg��@�*��|%^���-�@Q�%�i��
,��o1�]"^K���5�>���.�/�p)�$�]"�;�Զ�H�puA���btD��7��B�)��|F��:��MHbES��;�e4|�d�J�`���y�=���3�]�wO��Lp7ܗw��Ū�w0�y�4Q�lɩ�2�~��89§C{p8��8��q+��]`���觧N�s}�fY��tK�^ �����m��2�r���5n:K����p8���g��{M˾�7}�_���m)lx%��"	N���_�},��?:�|�9B+Ej��+mFgȐ���o�+�w�tGt�?Z���'�����I�%��p��p����k)C��mW��V�p9/�N�1$4K�L���<�8��<�T����dv�o��l�H��kJ�����E���z{�B��66HE5*��[ʨ�,>�$оNpW�/�K~�p8�!*�� ��e�~�!��\XWQ��s!65bBݟ����8~I��E���#��J��3�G���}q97� ���_�7sP�Vq�	p��c���bC�Ē�|
���p8NTi@�a�� 7g���}�RВ*ND�'�L�;b��_�H?/�<a ��"/I�~L4��n?8�Lb�s��MmK�|f�vl��w���{6K�o����[���%�����q|�5�Ġ��̸ﲵV��[�w;E���3�KXFBcMJE�����8-�vAW;�^_vSQ�q?����%�`ǵ�()1�S��u��&=|������������5}�����ES9�c�,mhG�O�ī����Q�b��P>2��P�샃��/��_���ȦQ��5�ߒ��xA&�ũQpw�큷\ReZ�o�P(��;���p�M�2:�b*�1�g��_6aj�0L�� �WC�丮�lj�B���g��W�����"��U�#�<���}'�#e�!�va��:��:�����y�e:�H���/�<��=B�����!ۆ{y`|�0l����9i�E��R,�3���"��	�����??���:����
U��pb*��`�F[W�3G��gN���0�}i�N&������ENKN�;{a�%��GH�|%�v�Y��>�v�XR��yR��]+�y��~���Gsu���D{��<.\�J�}@p ���SR�!s=I�����ac�p+���p�Ƈ�{�Z��W�H�C�8�IN'e�w���َ����ljHy�T�Uc|����-�ah$�y��p8FVQ����1�U���x�9�}�|1�M$���̞��=�E�7��/�V���T�:��?��c�_V�dj퇓G눭���q8�h\��Ͳr�:wIg��� �]�7i @_�F�G~���C1�GWd��鳓���������+xS���
�Ʋ��l��ߗҦd@p 6�?������ަ*���9������ZP��<�cfd.�� a��z�g�4\�t���IU<Uu��.w�9Q�{1�%���qR-�]��n�ñ
�]J�C�z��)mBpo�@"K!�J��αf��p���`$�%-e���é�������>���?���˙y��O$���Ʀ���G?O��ё	��y|��}����gp!-�7��1dRӛ���u?W�O���}{�_o�搡�����爁x���)�bW�6�C.��P�!�ؔ�0����Y9����Y>2��^����Q���ƴ_W�B��l�z��հ��ݠ�@a��/��4�6CO�Wp�pӘ'[�ϭ���	�vn)��p8���kI�IHE��@��[��~0>�����\�m�ve�m���b���?hyK���n�L��6���p8��Z������Jf>,�K�^��������c�����%��#	�/��{�l�mM3<�me�o	��Gch��4����4f���	��z�kM�������`1՘������+��0�����ѧ�ǌ�������J�O¤�a�<��`�]t��qrԘ���{{Ga��˃�]4�pjEsw{9��?ӝ��pn;虴h�6�x|&Rr�_p���9p��ok��pڷ�̕� \p�p8�
����z���1��3+�əX6�Y���k����/_�;���cb��� w�/;:�������������:�xaTx�v����|��-��wZ���3�mߏ�WX��>�l���!���>�Bu�i��[�m���]���q̯�1ڻ����������呓*K��ႻuA��`77$�if:�ws�����\P�}	�l�~;����x�J�e)C8��PX\���Xم%���U��=q"Q�w�UcJ�;����\�YL��H$\p�p8��^�J2�����j콖�&���
�f��4�ނ��M�F|�I@���|�e8�ڲe����'��]�.����yw�
�����yw?_���O��#]�8�����+���w�&�x�7}ޛ8Ҥ�+��DU3;�o����XF�`����5 ��N����>޸�[G�n,4���Աxz`�8��I),�]�����P�AAy{��	�i�����e�?~/*j��w���h�+��ox�����e��x%��v��m�I�8��|�_���D�o���ۣ� ���"�v����s8����)0����Ýc��^�P��bWpK���AȻ���S+�t���,e�\���4%�� o��)�9;�5�h��"��AVK�ϝq����'^;���0��rsEK��c�L�y�"�dSn��;gO[t0P̵���#��>h��p8Nk0��u9�����ۃ�Z�?{�'E}����z�\�8��{��Q��51�$�1!M�ƨ�h�&6����{=�qp�������(p[n������g�c���������yL�s�ʦ�j�ڽ��#5��Gñx"""""�R3Ý��^�2�cI�DDDd��n���
�Yp1����1SR��������p'���M����:�3܉��,�nV/i�7`�;�r�����%`:�]�_�j�Z�V��� """��WV�g��'�r�Z""g��k�y99ށ����Rp'/Qg�z���*���W�����DDD���|��0�����H�4z�p'��`�N�K�h��ZmMe�>DDDDDDDDD�\z��j�f��.�N���k��Tׁ���������M�60�Nޡ�1j���htY��V�U�hp'""""""""R:f����7�m��OT�o���������H�T`�T����u�e��������j��d�z��\P�ew??��԰� """""""""ecw"���z__��԰�S """""""""EcI�*��h�i��%MS�ה+M)�!~ """""""""E����N�Am>��w�<�"%�קcT�o�Ś�X�2���gQK����b�S��T��@���S�����t:��+�0^vü%�R�R����d��HW�I�����0i���^�S�b��#�Zw�w"""""""""�RyB��K/��^ 88�d@@@;x��K�_,�����
� �Z�1P��O��/O�)��l���������O��[�D��Jzaeҟ�e�Z��WK���F��I��		����a�Ƿ�����~��j*}4*��;P���jT��hk|4j�� u�����A���F+��U�|�7��P?�Fe�[��4��5���N��V�?�o�tz���u����gf����y(�����{����4�ml0U��F#��:��t>�:��SY�2\hj0|jA """""""��xH�{ox�NW/y�M$�7ɧq8��>�J��H9)�˕@��lhh�r��'NDJ�h�*g���FΥ�`u�g���A2hPo��/��BA-�֨u��;4�Z3�j�*���FZ��T�V��5M���O]@@����_�/M�+���s��8i��""""""""+�PϦ�J����z�H��	"�$�#]��2HT[[����k�t֨+t�c�DDDDDDDD^A�ew����L8&"���P���������ț��*��J�&�n4@D�FT��%"""""""r�V�w�6�j�:DD�@�w"""""""�+T,)�(�!�w"rr�w��������H�we���/�j��-�Өa�DDDDDDDD$Q�5�E��5���M�Xŝ��������'�:��J�*�������w��G���������2�
@� �	���aw"""""""�Kj�,)�(�!DDn¨Ri@DDDDDDDD2����KxU�]�
DDn�h42Ý��������2����
`4�T*K�����p'""""r��@$�A�Q�bU-�ʪD�G���3�]iC�F�a���\N�w""""���a�12=	����*$�ۋ�k��ޓ��}��ׁ��Z����w�1��&DD.fTA��F����܋F�B��PąIS b��s�o��*�P�ף����ոPV�s���XUj� i�&G� E�����+O���֡��E�2Ε�uNI�-�I�_��/�TH�^u�ե�z�N�нU$���'����D^y���e��< �=))�tY/M��o4�zi�5q=L]��hZ$�/=�ALM��������鴥��C�����������*�J"7!��z��J�W����L׻�G�_j�4�KG�ML|5ͯ�'��O��`nv��Ǯ3�8UT
�Ix���MD�V���	Q��.K��l��ʻ��9Ҕ���P�༬r�ш�@�&o�a��4�w�DRD(~;�����%f��Z���N��Z��/`4O���",,,��ǧ7��\̈���5��V��3R�)c:� *(�!��������C���׉l����b�4�8rƩawաU$n���;��{b�<�a/�Z���0y�ܵ�|]�N/��;�E�p�bɚ���gϡ��9TT�b@�^��=g/���Z�Z�Q�H�ה�Q�؜������H�z&�➾�0�g:��Z�9Ãq_�y��k�����v�1�>z��&N�����u�����"�)Rnj�(O�'�|��{_�:���Z��o0X���9�	�bC���ODD�Q�(~�5w��^١������HD����5�z%�r�k���k���r|�-�o�����}[��AiYO���Z�欉�[L�? s���� ��E��g� ɥ����4�̀;QKSU3� �p'"�b4r �����	"�~���xvd/����I���&�s�z�m����}�Wp�ͱ�Z㥛��[b܍hx+�0��_��k+w����fϧA��K]i�۔nұ�|.R�c�3�ND��ԁ��+�7�W""""""�Q���=��I��w'�ޟ��9��k����J!���a�@n�w'֍)���5�EY��/���A���j$G���=#5�)�h-��Q����z��Pܕ�5܉������WǸH���������ώ�{�e��K��;���K�����<S����J"^��;`B�4�m�N�{�~��-���R�wᶑC���'�r�v�DDd�<��i�R�F�[�Ǉv����n��b��Ό��ѫ�����J�n���	�2���P����y�`9���V���2���t2�ӓ��b�A����`���y�@_$G#2�a�r#nq裕&�h��Hۉ�K���:t�K1���(����T�Vס������T�����.V(~��5w�%e�Ƚ�l�LDDD�M��s�XKO�'�.����a>�r�-���a�x���1��j<6��<�`=��}��}�J+�x�qL������+ļ=GP\�9q��Ix���F�A��� $��\�;X�;��N{np?[R�3�ҥ��q��E�&�'+D��^�>�����JD
��!"""�U��X|q�x���'�9_��&ܜ����Y�.l�*ʯ�7s����D-��9Z^�~�h��LԦ���Fym=�to��h�s�\!V�F���@D7g��E��kB��E�������"��;�����](����"��)���<��:��� �V�R%�(%"�`3܉���;M��s���2��!럝�{?[���[��E���ů��S\�v[<:�:�E��O��AuSvd�aO���
����u8WR�������xn���I���*RpS���@iJ���g����{� O�ǏG��/�,c%����]����$"""""r����o&7���!�X��T��`>۞�"���+g}O�orS�D���4����9�@d��*,q�s�zhj���&]=H�����kp�~����:� ՞?h�J����&C�$`h�t�����C?�R���ѽp��
?ffc��l�?���g(�����5�-;��PI�)~7BDDDd�'����&��{b�W�j4x��H�
����,Ƅ�`�x2:�E�uM���'o��9�[Z��ykk+�[Smu9|���#��#]����Z�?o���. u�ahE}�t.]��j>1+2�o�H�M��vu�0Jk�P^S�u窆4��� _�Ӳ��Â0k`gy�+���v�w���
x�ΙF̅�i�ju��`𖀻Nz� """"���l>��^��M�^�� ����o�:���_��5j�ٌ@�9h2F!����a-��F�}?�Ĳ�1m�r��A��^����*���.�*����K�J}�o�z�9\Z�-��oG��7�������]c�ָ�ZG��G� -*�Ll,zl&����L��JٱP�&	��y�++���s�'�.$d������I]�0>��������8_Q%]���ty�����r?���z���(=uej���C��B�}��nR"B����K���*!,H�znTO�;���ߏ5'΁�A�5��=��^_��������Y�9,�5"�� ~d�+o%��h��x�VƋR	%a	�M��繵G:ޞ1�E���T���*�V���F����<�#�v����j]��5�O�j��W84��9>�,��q�M.�yQe-*j�m��e�/�R"C�L���&:����Z�쀚):� 9�����c�ƞJ���1Y���bs�x���ɼpYEe�..�.��bN_,G�{2��v�/&!�Bq���[�%D�S��Vк��T�9D����$y�y6��ڍU�r��f�^Z³�d^p'"r'F�cHDD.����_e1����g4�]s}qQ!��1�D���9z��¿f�rzY P�x2N�����w���櫊�h�H�G��hi�Š6	��"S�����x��	��I��܇'!<�-�VZ��O���\쑖���B�Tך}�(��~�q�6C�&8=?#>
�33?��������rZ4�����]O���K�=�:bBF�������e�"��)���"��-@n���^q�s���43[�������r6�Ęf��J�ӹ�&`��^Z���\�gR)>Dk4�j+ �_������{�x8L�u:�m_�����5Q:�����9Y�"�p�|��V9#gU7���{<�X���}\�N��q�Z�Y���LӺ���0�|����!2�["�^YW���0�ql:�'r4�x���O����c�u=�cq{����#�i���;��᷋7�5Ce9�s��Q����>A�]��
��}w���wG$G[�8QfSV6J�qy��J'Ww�͗����#m�0�K�ѳ���Y}��[�n���T|�#�q��L{r���^�=#o�!!"""""r6����AG���m�E����]c� ���K��]�0g�~�w����g�3�)=&���g �Gg��3��|��`�����`����� ��}�.Ӱ7�@�f��w�n���셶��p4ѰwKV�>m�<�Ņ�1��,���A_Q��[��Q"��޾1�}�UY�b@o��\l8����w�x~	<]AE>�zX�ҢBqw���&&��~W,���N�H�oo���'�!<"v+��&�NDDDDDD�u06�C���������޸�]"MdX���-r����(,��ně�w��G�tsJ��SҼsJ*����z\|X�� ��5�%�ӏ��á,��(_�8�/w�3�EF��3�ߞ1{�(�Ul����G��șD�!C��m!2������� ��?[\��G�bYf66e����Jԝ��x}��ڽ���2�"->N,����m���x�2t'�VÝ�F"rF0=����ܓ�rMq��l���c�☾}Mg����7��R&-���Z����<e�\��^�29%���p�U�������u�k)����m�thSWk��3_�:���N㥛���A]����wf���.���ƪ
40�E�T�<?;��N�"��M�p[�vk�:fa��38|�"�Z�T�W���=�1�k~5�:����8���9>
�}�ʫ�`����;T�YIDDDDތ��d��R�Ci�!�t��o�In�(��³�ֺ�N�����rMp�ud�T���q�����B#<���s�Xt�"����7 �ܵ��k�����)|x�X�e��N���Ts�+Рn�RT�W���&�/���R�^�/�wNI߻,�(,Y&�z,��ǋ�����w7���9����Ǻ����W`WN>�3;��J��������ș�����ExxpW�i��!��>7�\jĝ�:zC����}&tv\�f-���x�~{�\bƔ?M�q��H��x���Σp'⌆���->�k��'9d��N*}�9r���0TWA��8n,�<��jq)n虃܃������n�lXVQ9��=�OyE=vg�w���P�0�?f�lvp�Uh ><w|���Z��0��ح����Y""""""�J�o��� 3,�/�uL)�����;*���=�.�#���p�c���n��?�����GMJ���O���$����x�����>��{3G㶞�v�O�����xu��f=Ψ��|�/�L2/�O��Pi=ke5��:e0��Mh�vq�w�O��='�����~�&Uux~�&�x�>�9������`���åؖ}
�k�We��o�4y��")��I������ܒ�J��f�����^f� �A��s�P^ܙ&����\���n��;B��h�u�<���k���7��#�:{w~�T@pg�l�G�\���Z�,
{=yS|��̷���z����s�s�/G��u�pu�_���zC�0��aձ|��8�9#� '�Y--�Q�~�/�'��7%�G���	s�%}�e1Ý�����Q�!%*�=��������F��?����nv?���`w�7��xƽ� s����`��sF��ؖ��O���-�����6��ç��W4�I�DiQ�F�Ra֠.v�Kd�>3�'~�x�Տ�:��+�d��p9�^_'�hP�ԨP||�h�L��������]G��cJoҩ8�Ҳ����r{��X����"0?�.��q�*2�p'""""jB�����qX��$^Y�D�B��L3FhDֱȨ��yF���Rl;����G.\Ĥ9��iHsL��o�n��["/�7n�Ԩ08������W��J���7���,FuH�k>���k+w�Z�!�z�5��gq���_>3�ji.��MBL�u^d�/9|��8��r9��B�l�[>\�E�LB����&����?_���K���J��s=�4�������A����S��#gBz4#+��n�n�g��h_Ʊ��r��Re_,�K�,y��N��D]����/��t�.�BdͿ��z(5X&��<��2�v�D�>��{�g�_��Y��A/�X��q6 ����˨����qQr07"�G�K���#�f�	Wׂ�CEm=f|�˥}NZT�����h��zw��v��3�MS�h4zćFDB%�ǭ�����C�`���Aw"+�U�ܧvk+�����g�ջ�tYEe���"���4�عL�-�+5���=���W|f�h����V`�S��jX��.xo�>��Cd�˗zB��/@r��׍P_̙9Kg���;���Sae-��|9V=u�ٳ��8q V=#ߟ�O�MY��{e>Y�A�~*U�ǀ;y�妩�����OG��O�v�:�F�'8�_�i��E�MET��AwGY�yO|��c��ޜ�c�n�8�����0�k�����߱�23J_��d�'|��������/��2/ㅅ�����M�G44aT���&�3XÝ�����#�H��&�7��2ܙ�B�g�ZpO
��v�v=��V�@NI<I���r��ŏOsh�S[m=���X&�cq�{�v�3�{����:�����:���k��:�o�ۋ�Ŏ���\�wI�/�C[����r���w�(��2zDL���hT~�M4D%e�b&tNń�T����G��q�S��cK�(��(ơ������̋��D�/3�ɋ��W�cB�4��8�X�`��� <��3��6��G��u�V��ϖ��pg�CzL���|���S�<���_�mǜ��m���m����2�Z�U*1��5�j&V3&g�H�� _��7�0���E�12=I��_����[�nK�w""����@""wu��
���"Y�x�b}g&���ߋ��%l<�g�3�%!�����q�g�PXYO�������^�i��Eٟ�ɱ�m�N��� j�Q��Br�����̑��o@��]���K�t򿷜>�������G��`�ٖ�F���3�v��C�ug��TbΦ�xvDO��������e;�6 � ���DDDDD����ސ�Hi��	�p?��I����*k�ծc�t��~:�����-^\�{r<���L�x�!�v�M6�ct����4r���p��O�)�뭯�.��Gd���v�&l>�r<(�gP6��Cgh:�mt�|n,K�i�T�;��A]d��Px��tM÷{N��G��h�&�]4�Q��c������+��6T�cH�"�	&��`;��w�wβsH�������;�b������b�x�o��&��l1���i��2ܙ�Nf�s�����l��0?�s�2N'ʵ��4����4}lZR]�/v�cC�����npw��f�Y\�������+�`�G�'�6�h>Bзu+��k�,x����׫0��-R���b�����e5uXr�4n�n��{&�@�V�^���RK���8�� ���R�J�84�(��c��vd���j�$7�=0ܐG��,)CDDDDt����Z�p��?Y�x}�X�d{��|Y%����R'�[{���� �ͩ�#�=��jw�8ͺ�gm���"=6B�h�J����%e�wNkUrέ�b��f�,��l�l��~��J�G�K�?�����]�&�����ᆔ��6�Uwiâ��\Ol{�=""rS+�������U���M���Y�?������lŰ�$������|;���ۈu���cIR�6ѡ�**��:%osߜ>	a�&oO����۰��R�$}�%U�a/�<c2�.�Omŀ�i�j�G�"""""G)�����>j��{4'E�ud���s(��HԬ��UX��t�jl�oʶ�yxg�^x#q����r�ظ^�E�@bI����2�T�_���Sy7ܕ��`��7�6l7ʪkq��E��45��p��-�מ�ŋ�{���[��`<�O�e%e�W$""""�j�:��������������}�k���[4�K+A�	�Vf���A [�+��>�k�MA��:'}�_^��a�;�[�w���/G��#�`��߬1]��3z�c|FZ����A~Z$��X����탋Uuf��ʊ8QP
{d]�=��m.���o�7�Q��\�~�F���ƣud^Z���
^w-�vw/�cˮJw�q_�O��4>��^�h��Ps2�� ��ew""""�k��l"�t9�(�J���c��~�H9wff�%*뚦F��4'�`��]ۘ&8R�b��ı�|}�.�ң���j�Ud�rm,#.
Ӻ��{>C�&Z��������)�=�7��:��<��Y��S\$�?4�a��`�AT�7�p���r�;�S�)�VΜ���Ǹ�Q��˖>��b����m�8C�ɔ�A_��k��1�3Y7�ț�9Z��k�u��f"���������O�Y��.����ǆ�[8cC��gxD<��E��e��M�3�C�uXd5��t����s�yR"K��RC9e�&�!Һ"��asm�� ��m5��"""""�"�Z�L��3�=�Dl%�"5�:�˨��5�s�`�	��#ݮ��������׻]�ŉ�[�XW"I��}�K�÷�& �r��׻�#����n��R�����.9����|��0i�W`�>df�]����^xD�N�A�^�lD����}�n��O���R	vekj��L6@�2�#����_�W�5�O˶�Y��f�_�Fg~ ���-����AZI��h<�4��������L��N�=�t�4�,���~�����=���6	���9�vv����P�)1<�=<�?��zs��W��J��@_-jt)[biw���I��L�c$<��+�±����-T.Hq�t��N��<<�i*��W�Y"rk�!""�Q�T5������� ��m��V�ƴ�Q�T��&bf�v�G��xg���\�<h�g�c�>q���i��C�����q�	�z]ni%�l8 s~9�'&wI5y��~܉5'�5y��C�at�d���KS�债|4��Ax�?"��_��w�u�D�+��-�����X�=ks�)�>��D=��ok���B�@�L쒆�qQM���Won���;���������/�Y���#p'""""""Of����*�M	��;�d"`��m����G�t�{�Û%���ؒ�:+��� R�צE���k�{���r6�9I���Gb����M7�N����d�B磂�[b4����u��x[&^[�۪}�Vm~c�#)���	(����1�G;�h̗���^����𶴽}k�^����W��o�<�~�ע<b��z��DDDD�͘�I�����z�U�5ZK�
�;K(y}~nT��	w�<;~ ~8tg��0Q4!-��)(�ոk�_YB�����j��Ǩ������鸯�k�ے���N�=�����a=pK�v���Rd�/6{����0�C
޻}�5g
XKd�4�/F�O����Rڟ��~�"�f��:4���(gҪ��º+����"��<$"""��2��.���_�&Fc���>�^�J�-1?�����>�7n�-v�`�_W�'sD�������-���p���"m~lA��@FʓkD��)���NdW��p�bW��`,}l*&�{��h�~�2ܛkJ�4|x��Y�H���N��9QXiz ����A�	0y�ْ
�#���J�BQ�L�\OO�ʥLl�%���)�(%3g�(�Ă3�uŇ��D�Uh�]g/(�ݜY}k�0�_D}o�����2�ʝ0�����з�,/���1[;$�~E��0|z�L�`�\7�)�>7��8���((�;RyJ�ݛ2�/� �)���t������v�r ��?����I���������r��L3٢��.��6	v=�p�c��D� �DC��ΗU��U����э7�iQ���
kM4m�8(�]��edl�bPZ���;��n_���t��Xi}1'3�m�w6��^s����!19��s��{;����	18�[o1�}�����9�~���Q��;���	�D���T�+j/p� )�Vul��ā7\�ʊ�r�QkYzi���.>t'K��@D�!"����ҥ5��z&ǚ	��q�8yu W��˥����S�ʥy�ٝ����8���QTU�V!A��OG̔&s�QϏ�϶����-��.֗��7�ݞ�r���#n"�����DDD��v���}J�6^pe �uǨ�u�������d�ӟ�lC�}1YZ�l�����?8A�O�B�Ij��k��(,�׻�7k>j'n�V=��w1y��G���{ǡwJl������������/�ɥ�����ם%p���܉7V�&X���N�aөsxGڎ�Z����t�?��+k��� Ӄ
b vwNܓ�v)vcw""""""j��OD�{��+����.�-�������"Yخ$J|r�8ć���>3�'�`���N}�2��\��jos_a���Z��sl�Ml?~9��׿�f����Z;ʨ���D��2�|iJ�X�=,��1p��G�6;�������ʝ&o�v�q����z���m=ڹ<���P�gRm8�g�sp-�g�5�����Y���^�}sVF�7�)" }G����LV�'xe�n����+~��3c$�����"�=���#�|�#���5�u�p'Gq����H
����|g�@��R�ڎ��#�F%����7��q[������q����u�L��)�!Mޞ��`�T^s����J�	��O���i�1���������P�Y,��]��ms�]xzDO|��(����}���v�Cv���냯fM��Ε�t�`U ɉ�}:�C�H�J,�]g/��T,$!v٢��>ߖiS	$�5Y�NfnS ���Gqum�'\,0}��;�6�(��E�P^[Kj�uxy�&|v�x����:9%�q���K�����z���l�-��ܙ�MD��!"""g�ˏ�O�S���I�����]���i����ߧw��@rD�\����A͕ѯ���k�2�=v��Z�ʁ��Iې.	Q7\?w�	��gOIG}C,�S[�6p�������d�]g�妫�Z*��v�� o��9>
�\ʫ)��%b��^����*���OD���9�'�-�����\�hdP�+����r1Ď�)/� ��~���"#>
�<8�6ַw4Q������׫,6l�O�g�=�7V�5�~=���6��}�k<Id�#��w��p�u��q,�Ħ�i-45WR��Xkߵ��5A~>M���X�oSW,>x
�b��N/=aE]�� 5����׸�x�ɀ{ZT��Yz��&v���צ�x���[S��J�b���܇G�D�����Yw��ծ�v�C�}��-Cq�?���	�w�L�k�����M��v�C��D�-�-�%�]O�i�<��*��d.��A_-_�S�ߘ�������()c~���۱`E)�vѦ��a� 8R��04����W&D����Sy�~���gyD�D˒2DDDDD^���d�5A+# �yߟ&�k��jR�6xjX��~�,1<���ؐ@��O4��d�a�˦\qWߎ��������^B�}��;G[ Z���L��!�4�}R��ԥv4�4�����+�m�ݤ�w3��� ?���--2-iZ�6�5������b��+�xUI����؉	5:|����Ǯ��~�@��-�F�f�`���ME���-"8��+���9���9�O8�:�g�?;o�"��"p��}��Ɔ,��juzy0��Z ӌ*�|�F5ь�����r2��Bsk��|]G��Q�x���__�� ����3QA��Jw��^��h�=}���-�
۲�����W��X�fO!���YIDDDDD�x���P���=�!�q�x���ޜ(I�V����$��7���r�]xn�ztO�F��(8���3�`�s���ef����1�}���#��Ǹ9��7���+�+K]oT�w�9�@\m���ZZJD�5wK�m�XS�B1w��,�9�u�xy�VPˑ�g�^p'"""""�S34# �"�noMmq����'cʜ�q�|�`h�D|v���پ��Y�c�����o���-���f1�b���g 1,|�\ȸ;���שCqo�Nv�Kd��c��^��+A�^���X�{oN�]�I��̷���&��[X�����T���-%"{���y�3��in���� ̛5�!����ۑWVe��Li�����]��Ϧ���}s�n��?�~v�Q�x�Sp�'K����=2��2e����(����W�n�d=QX�Ǥ������c�1k~q��?r�"ܕ����m#p�����\i���/�8��)�����o�쉥@�����~��75�"}�tpYk&����V~��Ոr+�]�����OS�zT�7�N_۠���ז���X�9a��`,|h2�D[._��d.>ݞ	�;3܉�\�#v"DD�@<��fi�!KiM�Z��'��������ixn�:�o�Q�Ѵ�����;t�e�2���kJ4���i��z����K���ʧ����b��p7b ����`t���O,��g���	M��m*��Kգ̕�X����`�0�T`���|������H8UX����&oOă_�3�Z�p�V�VX��D�5Y�oAE��Vq�:��jM��w��������lÈ;Ybl�Ok�k�~�ֳ=��5��V�w��I�����rYw0�}2ޞ1Rn��H"(��+�Lvs^Y�]n���`�h�����J�]�|�Z䗻G���ɱ���q��u�����յ���Ȱ�c����D���ʦ�U�3�5����گ������WY���+)#�9W`2�> 5#ғ��r�gY��XSRfDz">�{�\z���������8��R2���DDDDDDt���AQ�����[L���\�*�>y�5ؒ�W�	�+S�`z�t�����o��#g,�O���vZG��_j�C_ø������˲��|{���$��0����b �96���W���	��ZG5=�Thg����|������~�L�h��o=}w��|nd/��M$\ai��!]��*_&��<=wv�͇�HKA�m�DDDDD^������/۳��u����5Pm,-*L.13o�	��b�\缥�����C�ə���;���e��x)V>s�D�9��D����1k`���mXu�L�&uߜ���N�ЬvA�c~���x/܎�i��Y�2���ƾ����l��������6����-:t�Mbr op��ҭ-�;p
�`�������~�������{;��G,��n¼}'�D*��Q%7�U�Tޔ�2��/"r���j\R��C�W�m���I�G�3z�Ǵm���L��a?N;1���u����������;��8Qe��K����v7�m�(�탓p0�o�ً%��,�l%>��S�ܨ>rG��/�e�Tr{� zX4�W�A����`im����5U�<4:�'��m��r:�2�K���c9���j�>�O"��9Sly;���=�1�k��n/�[p�X��n�Y��&���%�Āɳ6����>��<�V���NDDD�h�O��Z��^N�2^�����3IkeV��q�S��i�P��J����"��!_��A�
���2���mrƴ#�EQff֠.X"�n;�G�:�)�h�9�kL랎a�+�c��=���m~�������ݣ��LHg����+��I�W4Vݓ��l������}: =6���U���~�d|���̱s���5Y6$�W��:۳�/��o�j�;��K��zSw�����8UT�,ij*@�����)�6�b_���[��;0w�����F�Ӻ��-�ۢO�Oq�f��e?ٖi����̟��71�b�9� ^�_��2+ʒ������I+��ӧ�`,)CDDD��ϓ�J+�`�,��J���~H��\
��tU�!���~�AUh�aQP�B�o�AÀ��bĝ���3�������܇'[Uw��D0|D�$y���'s����>����-f��KJD(�$Da@Z��G����֦,�wO|��lV�5v���;>Z�y�r���Y�`�#C�ɓ�]{<۳/�@n�Y��S[ISnJOD���p�y��d���8GnG�y�}D���h���pw�ע�Dm�^�=�2�銲�:d�I��EWk���-�K��ڽ��������I��W�Qe���5h!g�7E�ޘv����l����Ԣ���dY2���m���\i%��|���<��hxL����2�9MDDD���됴���i�B/�T��ґ�^ ]���hI���p�4c���Rz*�z��Tj�.״���*�t��\"��n�J��E»Z����U@SV
M�ih�ש��Am�C���6�Pg]�I"r�~�;q/~�A�	�L���N��IA���8[R!�=.����`��!�䇎�"�lRWI9��j&�f�3>\��fMtZ�{c����G�<]QPQ--oi�W��Q�
���#���V!Ah�¶�s��W+���o''2W�9���չ�J���_�u&^ú9�v�ڳ�¤�cQ����=�p#�����I����6	��xY��_z^_�����6hk������M�-ܗ9�'�]+���)�P=�������s
� Q�ݛ��DD�Q3�V�Y��Q(�F��C@�W]��ue�d_?�KOW_��c[P���(�aO#��	��'[#2( ���?Z�ʈf��n(�s6��K�69|Qo:��i�/�܇&��(O}R�Dv�h,[�RC���$r<s�۷����"��[Z%gA�0�[C�����T�9������=�7��DVyc�윇�Z�E�L���|�U[�ҭ>��y"��z��؍��%4ٸ�TwS��b�&�l9䉇v*�J����ُVC��-Ý���Hy�
(�������l܉H�ƪ]���ّ��DP����z��"��L|o!��5A�(�VG.\�-,F~y�Z������z9��Ti���H����o��G'�Gs��-���9~�pz%��Z[C��Zݍn;�\��/��簆��m}��~�x3*j��^Y�z-��1����SRfk�y<5w������VW�}�ۿ���3�ӭۉD��7�Y��JDDD�r�e ��]��d�\��t�\����ۈ,�'�Y%�w6l��y�⁛10����b߹���p�B�E�q;J�#��U���"��쀀��3�������7�	�7�o�i���}��㐦���ǽ;���1�R->UM��d|�\L��=�Hˡk|4�!��͢-ؖ}��}J��S��x��!�{�z�%eD�ۿ�ڍ�wi��כ���;e0>)�dBA�����(8@����z�D�B��`�[k�ȧ��~�0��O�}�w}�o)"�|�����iC�����[�r1��&3LBŀ;9�,7p�h_`����r0�͹xad/�ۯ���*z��3��-�y�"��x1Fuh��삑�S�M��o�9��m���������7&�"h�ΆXs�l���/¸�������#1<��`�xQ>��͇�ƚ�V5��$*#���;ڒ7��*)�5��/XDDD�(fGAD�@�?�5G��%�1rD����L�,*�g��CTP <ي#g��W�\�ЮN�ǳ��aÉsx��+��D#ZѠW�og[Q��I	D����7��k���Hd�/��9
*j�������}xaTo�ݧ�٬��ϡ�� ��V���MV�ANi�\:��竬3$��V=#O�z���	vZt�ܘ92��������d5�?�v}S�0�K��n��	��.�/���)Ė�yXt(��l/Y%��ܽ'��P6��d��<�>��<��2�-�eT����ީ/}���R��^WÝ����(��w�������O�b�?�⃻G{d�QB淋7��]�)�n�I��)�{3GbP�Dx���������92�@f��Г��i���p�B4R����׆(7�=�43[�����p�z�;�\�'{��M�v�qy>�k���9��XYc���=j���[������N���0OF��ߒ�ُa�l��u%e�F��#"""�Q��z%���~3�+���9��Q����Sbf��<<������8S\.-����M�����M�`P��y�x��p<�qHӌ��O�<r�L�6�W��z���N��~"�oiM�<�{�3�+"U��g?��Aw�+)�R��o$"""�Q]�xC�����
��r���[�C��8(�������ri����L�|û��a��,�:u&tN�R���פ����{Ѡo����{s
��uS�Z��0n��M��@�
/�A�G�9�.2ܽiO�~G<DDDD�Ph�]���ND�Eۚ��p�p_��zl�&�+���q?��f�s�u:���r���R�ꐌ�M�n�1P
����)�^�E��o�'���iDc�}�
�3����χ�d����J���L���5�.�!�w""""%Rj�6�^4�R�'�V�'���O���='���xtH7���]�@�7{����;�[Z	�Y},k��`j��rI��&�4�Ѵ�e۱�}����]�y���	�M�GuHA��8��v�w��uf�WD�]���p7h4�������3(4��j9"R7(;TYW�W��˟�l@g<:��.��*���Cr阋U5P2�q/�J����'��Ĉ�IP����!�O�u{��\��_���=~�<�_����m��������TyqvWYM�tz�E��+��2�[�]�94KD���LD�%~Y)p�at�x5��gB���J"ʳ��n/��a�tl���wƨ���uA����x��u�fAgp���vG�"�]L)����O����Qa.y=G/��ZL�6�{q��y���ErY�IMg��J���7uÿ��)_tp ���;�=��%�˫@�P�,�"ҿ��o���n3J�u� """R �e1�{"�qü QjfYf�<�3�;�bb�6�6ѩ%g�����9�:z�d)>��Z����V�'Q�}b�4��HE��hh���� ��#g0o�q�+��r�oy�O��?on������mԡ�� e�	�3�{��A�ࣕ�S�1�+I��ΰ�|U����b�l܀�܉���I�}�UL�v;<Ɋ�N�j���c�$���c1 -N�����p�h�?�'2ֳ/�#�|�\#|�|��������ʓ(�#7�ţj<�&D�kb���mk��z8�R�i9�;~N.��m;�o�2o�I�q�@���Z�|`<F��@n�Jʑ�'�vǽ�:"����x��|*g�UD�]���XR��0����Z��9:D
���L"�]k�t�V�FRDR"��`pdP }��V�7Ie�uh0PTY��U8_^��2�^8�&;��ip�X����N��w�� �߾�u�F5�:����t������b���"βy{�>�|s��߿o������k��Q2Q"��a�1�[[y�nal#�����ٳ�qu��J�]�g)7�Rw�D�y�="�fQ����A	"�Q���R�z�<��@��ܹ�C������l8��vF��������cS1�?�Y������uJ����.���y�l;i�|���ݮ�k/_�n/,-CDDD䮔Z]�m'S*���""��kq�v�Lst9����l'޻c���u����ǧa���SRr=q��}�;��H�i=#�"���wic�7��p�^�����%1E�Hy����,���,'�|��(n��c:�6{�6ѡX���x�۵X}�,�婥�Xz"���	��������[��A�J9��.W��ADDDD�I�Gj,)C�DJ��9Q��'d��}���[����@��Y�sgM����K�z}�疒��=�1�O�������=�Wљ  ��IDAT�"RU���w�GZ������^����GD�LJ\���5�ި8hFt=~-�Dm�Ǿ^�//�7G���^���x<���<�r<QWr�4��3}RZ9l�j>;�m�!uh�{��DDDD䶔���Y�x%�~�1Ý�pf9�G��O˶a���Vݿ[b4V<u+�g���-ބ��r�}��C0�k*�uk���[�%d���Z+2��l���Ւ2���Y�DDD�L
=�72�K�h*��Bt#��go7��vR#�����3.�5FtH��ێ�ߛ�TQ�:�l��ɱۡ5�tJA���?'������R����o�;��9���NDDDD��_D�sM,��DM`���h�<��l��F���v��1�����uƪ�g����X{"��GMh$7>�!#:$#�B�|G���1w�IUՂ�A5)��K�~{����W�^��V��!"���m������W���˚,i��e�;�e?m;y$O�Z��� �˟��:����ԬǊ(c;������Xx �8�=9�V	a��.��0�M�ń���W�5��G�����-�9��0?Ղ��߾ՙAw�j�*��������؋H����N���Ȝ�I7A�_�[�3��x���6�f�D���=��Lq�efc݉s�t*�u��DA~>rY�^ɱ�)]�f��!.y-��h�a|�������RTF�g�倻Z���w#��DDD�PJ������gB��w"Y�p�md^ˮ�X���J���#��k�|ZG���!]�Id��9[�-Y�;�@�Η)+�Z�^�S\:��@�Hd�E#=6\�͕��l>���O�N�!Y�#�}�]��On��9|��JI�-����ܙ2���a&�5J�T1Ý�	ܷ�i��n.:���E���1r涽��{�'OW\(���sE8r����8*]����p�������F�"5"�ҥ4������B�̒k��:�r=�hg|xE�\g4R������LD���D�l
��ss�~���%����p�ѻ��m�� _-}}�� ��ǾZ���2���Ҹ��

@Ym�<?��E�Z��KY���BYM�*kp4��.�Da�U���gG�Dy��`R�� ��=WV���er J���=?��5׉�_\U�?/�n�q�S�1�����Β�!^�[�]]>�zmծ2]��iQ�7�W����n���)�N�5������ZD�����"g��D��z�^�jp �O�b��S��u\yF���v���1�_��=������j�Hq�A����o���^�/�נ����ٻ�6�����v���qb'q�ك�f()�P�@Kݔ���JiKK�e�2 !{�A�r�#���%}�_bǲ�%[�u��W�w�i8>�=�����b���M�Ҷ�������/���[��יo�b��!5*���@#}�c�&���'�|�1/��@_D�KSL�?�<(P���s�݃g���L���H�e!>XU��7nvg��W�����u���{�l���^���"���-��c����c���9��[����`��lQ%>:|��9�23:�����+�&oN!>=v����s@�?�=5�j�8Q���ힳ�l��Ru�����)åp���~�j��1�]%l{��S�����oMJ��T��+:�o5��$�Z�^!�8�#ZG,7��|�t�g�1�c�a4��`7�d��[q����5V���o���C�{�1ŉ����.m���J]#>;�%�G�KA�Ma�u!u�+��{ݠ�DDDD�$Ӕ�C�ɜ��C���M�S\
�M]<9,&�[2�MK��V��Ƴ�p����+M?�7?�d;6���~��m��/r{�}�}"�����M��J���~8{4�8p�5�+������%��Ȝ�N�^��^;��q�Ww�ڝ=��Y�˖YR�^�s���'�����ըo���K��p�:�㖓{�{��{UK���L�4p��&�v�z���Rs�������م!���!1,�{��y��Ӎ���.��Vn�{OۼMWۼػ�� ߝ'?��������ӕ;m.W�����9�\
�ۛ����7���Ϯ<Oџ��;9�R���Kwl��ǜg?��qC�Y��r���fl:{���ºӹR�N�%B����U��������h���JD��{�D��ۛ��E$;��O7�����ݙG��'��ݱ]��b.�>����Y�M��!���=s�,�U�bs�E��*�oK�]U��we�Ļ'��{N"�����������n2�cfJ<���O�f�t�֓O*�D�(<�HBlK>�:>������Q�a�;P�*�K.U�I�����ؕU`�J$�'��"w��-e�z�*oy�DDD�����H�O�3q���g�T�9i`�S�Mc���E�;���0 �Q���4���J_S��*��Ŭ�xl;�g��ק`^���D��k���O<ޓ7����}`�秴��C���� �����v@Q<��!��eu{q���Sٖ�6�^���p"@���&�[oo�Z�J��㋦H'I:zu�Y��5Bס�T����aV��ќ�.��+)�f�N�Pzh�-�+kNfKSjtn���C%�D����Bl����s�8YX�]�~��{렩,=""""�`�y����P�-����%#���A���}-��F"5:�+:]��͋������e5�]�@��j���.��N�Kӳ[�"�W�������N����$����ž�B��*;{:�"��٫�}r���u�d�����r�᫽p�3[�e������r�,�;N�=��-�Zs�*l����G�E"9"��5p�B��R��#
총+��c_��o��m�6���1Cpèd���ۉ�u1�������n����t7t���2<�#"""y��^���"���a��*ܗ�[���8�_-�dU�,O}zc灻=��p?�a���c�;�{�p��=��ok����2f����v�������u��=�{;�Ӳ�X��*��%
'O)�7�fu{���f�.����HfI@v�i�B���Z�����m���Ӊ����풘~��.LM�������'�pR*d[���z|}�D:��<�/e�N)t���<�'��)��?mp���Rƫ^+y.n���e�N�«�S�MUv?l�!B��y������h������v�^��z���P�-m�*��m�ƈ�t�R��GZ-�[:��s���
w{���^�~jbb��H��v�j��D hK~���}���l0���N�7�����A�'���L����Vh}!'"|�s�P��P?L+�{0}p�c#\��x���x�����e�W��19��1)���U	.��^U�΀�����J��7D$k
ׂh[��l5���Nj�;��*p���pdw���n��UBAu�K�ᨏ���b��{jT�`���������V���x�ޠ��}ǀ'aݙܶAa�}��"mοXS��y�u����W)|�V��-�Kޣ��P��9۪��r�I�T�	Ǩ����H�k�}=g\�� ]�58WZ���)���WV�SWt%t��
w""""y���Ox%�	��q7������/\�猳Z.����������I*�E���D�ltp���r������� T]���[Oc�����k�X� x�P�l�C]�����4����'D�{���W������U����k��:����Zi�O�-8|�D�ڋ�3�}�!>41A~�	DT�?B�}.O~b�5���F_��� 4R���fi�Қ�f��7����<����?7"���Uu(����C�n���^��x�,yn���e2�n������A���c�0.!�j��s�w1(��*��c��:i+cg��1���k��nI"l<�gu���QN���8Â��3��mڍ�l�}Զ{���]���o��m���(�� �J�Ǯ����d�A�\�x���
��ZǹG��v"t�2(�j�㵀�.�R�~�\� \L��?I*ޣ��x�J�W�5�ۮ�!�"t�S�>O��?n�,t�������H��[�,�g�oqϟ\�
������L���B��;��Kߋj��Ee7��6C�¤��g�\�r���pLO���Q��-�j�6�s���j�z�Q��ePn���T��
QWצ��K^j���̖�x��������F�[�8�G�e���";���U��p�ń28��B9"*�U� ���@��ZD򡸶N�y�������<�@DDD�%�
w�/!��+��!��I��տ]R'Z�ڝUh�׏�0p�WU��y���Y/�8Wt�9nv�߽c���κ�|�D���=�B<�7���C�G"%2�b�g����2�Z��Amuz�����v���^���D�;?ר�_�:2D�_u�{U��˯�[^+�#lEE��6?�����f��!��H�n���N���K��L�\���x=i_v!6f�t����@���
�e��h',=��W���`��tv,>�D���������-��h�肉N�����J;�u�z�OP(C������)`�:��;Q��8t���2WTy:����dG!׊:w�<�W��Sw��&���B��X8| �*�^������&����@tL� F�������,����]._@��@��#�ƙWn�Z��%<��a�{=�Z���J������U'�����0!ѲE�7�uj��v��u'���99�J�6��R+���cJ�
_Q'�����%�������
܉���d��A����h}�I���,��NF�%M�X�>/�<����7����91����p�
���N�Nh��U<�܊Z�ybP@[D����6���D������J�/�߮ه5߽�b�J�\�/޻J]������ ��Mbs~Vy�B��Y�1y �D�-��Lگ<������v&W
ܕJ�W�<�@DDD�%Ӗ2l�C$?M�+3E����n�G��q5p/�m�#�lC�V��F��]�����X�zY4|��e;�_���۫�S�.�I�����i9�s��z��L�=�EX&���t��ű�2��`5R� �#�N�����뼒.=uS=�1�4 "o����kY�>t�w������<�l�����	�Ad��' �5kh�|�_�9-9��~����w[V���h�w?܌A�A�`;�}l�$|v�ݶ-v9خ�?mB�|l.���^}s���j��xD2�=p����<Fi�k'=����W�_�����.�e9�o;p����� \��OB����jOv�����1Cpl�/��*w�Ϩf�N�},Cw5������+�Gb��y���u'����kIz2�A���<��}J�/��"H������ȭ�Q���'ǫ{N���:FԢ�v�yZ6���.����ÙV��I��j�E�[-����ؐ@V[��"_0�˓t���,�_g�I���ز#3��k5_�R��o�ĭom��� �A>�a��AY��s��~lQ)��[������	o��	�cdK"/����5��2KZwo�p���IDN��O"r�l{�s{�I�^�\����^���# �90�[���.1�j��^oc5��W+�}�P�.o'VL��l�o��������]�j���u��g;��]m������C�5;_�,N������03%�;\���_ۭ�ߛ]h3p�U�p��{�_U+Uw�T���%8~��f/��
��{��~<w���]���Z�y� �W���@��i^j"�>��F�7�����E����<�������П7��)�ӸV��;� �5���ѳ}nJ<r3�2�./�ך�;5n3)�7�8+]��w�R̺R]��7��իQq�(�laK"/��L���C���NDDD$Wr��M]h@=������[n]��BQz`�l������}������ןε{?��
��%J�g]��~��j��V���Od�Q���QA�xh�(�s�a8K�Cyi�<�o�;� ��9ew�����SFH'*lI���#_5��v�'�|4j<2w\!�������'��o��ۂ�ڴ���Ү����I��xj�!�s�l��E��G;�����w8�?}󬶰��K}7<�tW�5*�0�l�@0�vAJ��e����I��*i��߉�C*�M��n���DA��Ź��ޢ�7�/�������8���*-y$ADDD�$�@�^ A}�Di-�IC����e�����sǏBa�|�E�tv�0�0t^-�4�F.G!&�J
�<���e7m�P�n�j��̾�=�Š�"t��J�yi	������{�7Z��Ū��34�6���h��������+���o���6�Ta���k�|A�a�=⽱�v��ٽ��[����U��zwM����[{��i�}��C�-���w?܂Rc�"Z�,�j5p\~�����7��2�=���o �������!"""�%��&�p�=���>�-|x� ��E���K�ՉCQd
��,9���9�{f���H~1&&�X-[62�*p���������͇�ǥS����+?�5O�?w���o?.��!og��x >|o����#�x���v�7�ȝ��� ���3���[��/�Os�������6���)#\�omc3�`6�ͅ�ĉ{�g�1>��f�GDDޡ��;�Sȴ>������7ᥣyH����ϔՁ�]D/�l����I����\���}шAЪTh6\{�UO��7ڜ���kbR�����f��+{NY��qE}���L�Tm^��|{���/vagV>����꼭OfI%�X���������Шw%p�������x��t$G��������Xs2�[<#�":���'��5�PP���N����q�5�������""��x�/�ȵ���a�'j6q��D�&���um?�7�-)�.�|��7���Z��⣱��z���'<YPn���w��N�T����Q�k-��UJ�n��F��}ĦY��5�ȯ�s��ݑ��r��t����ُ���� iP�����un�d^����?�{w}��b�Tq���۱�g�1|z��ż�f��WGb���oƘ�ȶyUW��T�:o�)#O��'Fa~Z�y= �$��/�W�@N1֝�E����U�\�g�+�8=F�	{.`�L�;7p,yo�p���ID�d2ɱ3�%��Ű�;�W�XY+M]%*�Ws�
Y�ή�*��&g�˛�N���]��br��'�k��U���u�~G�K��;_,���"���w�qi"""rM%"""������
w���W3A�uF��������h�5/-	iQ���AnE֜�����m�~vj"��C�~ί����#��J<4{,�uM�lhDFQΗT��K�����<�<�v�A�QoJ
�s��Ǭ!	V��1�3��w׵���[SGa�蔶�[���w�߮]��V�ǗNo���='��g�@�J
�M&��sr�DϨa�NDDDD�g`x0�~9bC��f~Z>~�,}�3��;v��U����lh�磶xZ����3��]�T2q'"""�T2.�0�����|�¶�]T�����ffJ<R���n;1)?�7Oo<�p���O�+;��x����w#w��m��y
nx����*�T�b4�`��� """"�w݈dL��sVi%~�j���R��S7���G�-�ެ�x~��7饟mE�b�ﮟ��/~&�lU�Σ{�-e������,�<
�<|����Oq��DDDDD=��)�?g�^��4�L���ݸk��i.k�烹C���d����Nm�5)�?|6��a�;uF��2DDDD�N��iQ��%�1����I��G�@DDDD�n��}f�� �E5u?7�[p0��b0ՙC��wS�+K�#4*����K����\hU�����{���Pt+��B�{u(q�D��7�be-
����X�NDDD����~?st|$�����zBBX|4�D��Jju?'G��}߱Z��}'q�4�b"�b�p�+�u�8�1}p<��I��@-�Q�kĩ�r�-¶̋ؗ]�&����DDDDO��ퟹ�F""""�� ��t������B�}����1cH�^l���M�/>�bqV�;G�O��&`ńaX4"����a��׌�xi��6�[��t>��,6g�JW%��֖2 """"%�M��;��KYDDDDD=�`��g��ҫ�=�eH���h�?�~?^�{��stp ~8o��m����a�1�N���@��_��i�i*�k�w��
]#��DD��ǜ�\`RkP8j>4�uP7Ԛ��J�k�0���ڷ�yk�)Q�����159Dr���w�ŝGAD�GQM�ռ���[�u�E_�VM5LXs�<�a|R�4oҠXP�D��G�ǃ3���=��~xl��q_�{�tUM�m�-e�[6EDDD�ϙ�;��������P77Bi����&(��al1�k�R��Eo��7���%�
�Wv���+�?
%*u��&�F��&���m��*-��2��ܤ����:T~��J��l.������z�y����U�H�o�
���v�O��S[u,�3���E�������h�q�Rƒx;n��?.�.���U?�=�O���ߏ����yDOa�;�����E�_�_����k��-��MB�|Шoqz�1q�(�5"��Υ�3�̙��E��p&})1,Ȣ:�����/�=���f�i�9��@�>jU��"L_}���������a��|��{G�⽙(y��b~Z<AD��~��6>��`#rʫ{�q9h*�U�����ȫ.�)P��Wqv��5�
���#�10"��}"���A���V�pnV�DM�KU5*%���N�?��g�1����|Q��Yc� C1�ُ]~���m�z�j���MGBX0t�z��h�^Lz��5HӅ�J�.(�[���9�Kr�%���F�;���j�C�����3���%�k�a�%ѻ��i���1!2��� U[�)ټo�j��l�*�U���x��п|�k~x�U<c�ˮ5�b"����fʠX���7���ᡳ=�x܉���<ؤ(�H�!C��r8�����Ve�/9�Wcu��Q+��TJ��j�r0b뚭���7�H��:���&��}�y�ilF�� ���c�[[��Pk^M^� >�V��
dT�#%G�ⅻcx\d���h�q�u�p<�����^�~F�	eu��D�>
wLHë{N���[T��0����cΐ�f�������I���د�:���MЬ�$�u����3#\�]z��]���.nu�K��ŕ���ɂ�-�(=���f���:���Uxv���ŵ�������GVؼm�y�����e1Ϫ�L��#y��p:�ғ;܇��wg����tx|��DO��y-�&D�7_���3�ї���DDDD�(�W�I���uP'���Px����Ư�~� �a�'��h��*���.��M���7o�y�`qɱ=���c˦#5&?�h��?��(�:Z�
��y��X��Wȫ���1x��k �����s.=�E#I�A	�;�a�6�\�,����C1:1
K��tMWO�|~<�*�,U�����`�{�a����;b���Ҳ�6A}�g�KDDD��������e�6�X�7V#��q��Cf��ڽ�ּ/־o�ҋ�v��c�\�=%r!Z%���w�:��U�p'"�&��^"����	�K<����`�����w=Ŏ����ˣ���7�aRr�����ΗTJ�Y��,�R(�b2�RU=>>rwNL�n?,:�{�=x?�;��2�ǳ��-�
��H5� /��_�ۼ]��X\
��tƈ˩C�{�'E��[�җ۵�?�l>��o_�6���MEI��-��6Y����w�	y
����mR?�����c�B���_�������}G���Rp�5�ud���G1<6U�� q������1�hq�͉� 7�ӓ�޽�p��{$t�w�R	""""��xu1��;���F����g*Ez��o{�S����'o�gb/x�]\���#��v�OHm���X0��6/�t-�awܕ������O��pW�����F�75c@p��/��ƥ��fLR��:>;���,����jqn{/�8EK""""O��l�4	A�Z��Lg��rH��C�64�H��>�bVL�_��J���=Kp�k,z���DDDD$[��q�0#b��1ĕ��*�!�B������[fK�a\�YZ�/Of��Q�m.ߜ���eN�O��-}/.o��a��{ǋÃq��X�5��t*[��}�&Ł�+��K���"*���dDDDD�Ι�������:lo�p� ���xt���������{�����
�� m�+
@�2!�I��r8�N�N.��㎧I���-u�%��7�#�l�����\z?�3����%#O�Ԟ��/!<H
����ɖ}6ϗT�\�[�N��NF���j��;�H�;y�;'�O�MD���18[\�7��t���G
V��a�z�!����J-�m@���c@��>�҄����B��{���}	��}����74�b���r�t��g���i7���8�C�'�v�-L������FX,�u.��jD��Xߝ9�b��_���	""""��a1���-s��<y�,��.ę�r��������8h4�0��0Z�拽;������q��U�NջV�����-:�9�� �������V�{UCL&8�q���j��� �_�������oBD0f�%��$1Hj{����\ۃ�
���U�5jxy6�W�3���q�b�k#�*�ϊ�X��'n�������O���ǰ�T�������S�V��oh]���k�s�u���03%;���r��]�LQq���x`ڎ���S�q�̱6o��L���'|�~T��|��h�x<�AÈ����£�H�����h���l?��u��S�`�z"""�O}��4�%��
*�=��Ե
�Y)�V��_4	�^�<p2 �b��E�����p�Ri����Yv�MM�ElH��e�_3
ϙH�k�ADDDD���<<k,���/������(��
w��DDDD2c4)����	�Kh�h@�b4�^�.����l����Ha��̋�sǤ�m�{N�����w���X6v(��FZ��LA����5y��e���O�M��V� ��jз�d��_��\T54����:���k*h�*i<���0j=�D����������y���<[j)�߅�������5����:B#""""�5�4R��I��V*`p��P!�R��2��_��R1:�j������A�m�[4�a�.~�����NF�}j�~��o�g�W^��X��~t"�,��J�Bvi��:�}��i�ж��-���Y�;mdۼoO�o=�'N��ڦf�ϻ�]9�;7��/b�w����Dx��U5���9l���×��U^i��b�904bqcz*��P?��uz=��bwNvg_�~�h.~8cJ�='dx�Q�����)�����l?�������;�L5=�ʱJ�(�`����v�!�=O�UwǴ*~9b��ŕ��'ې�߻I��&&Fcᰁ�p6��zfI@|��.�jJ����x"��V������*���[�_?(_9g����R���l�y{-6��A����&�L�`�8��� �5�؝�9`7=RPdu��S�))ï�mŗg�Y�l�xi9�U��ɉ3R��7Ǥ�fbH���խmj�Km��.����""���M�7��߹f�Ӆ.��V��񸇈��ȫ5+|�ijuS����o#�Z�0���p���H
��ϫ���o��Z[�+��-�]��ݷ�+��h6f��VF�lo=wo�;����XPS~%��c��K����{����m�s��v2�-���jl9�'���O�"*������gJ:������[#!�D����v![��`������-xb�N<�}�����7������)|g�8<�t���>���;Ϳ�m��r>'����y���DD�n�y?q��xqE��7�>g��-e�����&"�4zx^����I
��(r�X�Z�8،����'}���|��(��:����,{����E: c�"�tD2V�ʶZ���R�[Q��[�RծU�{��M���}�W�]��QatM��ۈ��&$EKml���Zlo����|��}�c>n���F�����]�"�G���럞8��g2q��
rV�k��7?���|��W�Di��ؖ��O�u+ң��+(��'Ϳ���p�R�l�, ""�}�Q�F��d���X�a��YR�T����DDDD�M<��]����ag\9F2���"����MR�{��j�{���9��5{���6[E�-�Č~�������N�W�s,��#������.W����(�#C U�ט�w{�g���>Ɵo��%c�`Lb4��� ��RO�ិ��j���3}��;��'o�����sێ���|���xa	^�w+Oe�����]Q�E���̲�{�����7���;05���v��u�������{ɭ�����%"�l�~>�a�x�[ǥu/p7�L��#"""�����t��E�
8��� ������ͧ[��mVY5F��]i�QGD+�n=�vÌ�q��iT� ,|��Wպ�|_�~���T74��Ŕ=�R�V�:�|i%~�fw���n>��)�������8UX"wx|�6|y&���u�:�UJf'��ä
���i@���F��p�R6eeccf�T)o�8����p���������g��.^�BD��KO����V��]�#w��M%"""�+�絔�I�#V�h�?h����zl��s���Z|�V��x@�����g]��YTٿ������O�\( ��H����r�/��s��>�I��	���u�h�,����B1!>V��^߬�+��o;���N�eC#n{�3���R��.2�@DD�aI�`x�`_-&&�`o����4����H��j?x��
���1F9�����y�SťRE�#Z�
#c`\\��EcHD��!<ѫc���˂}}�;n�����'E���)R�~�'_H��m9RP�W̏�����O���o#��I�ǘ���S4[�	��J@DD�!N��MM���2(���]a�+܉���dJ����������a`��z��U�v*�ADd��˫D�|�%�Y�		��h�|���Tw��S�Js������vL�Хu����;nş6���6m�y�ط����^��G����'=�D�c|B�y�5�^⤐=����?m��܈��s����ڞ{�	��t?�p'"�
��$"7���맀��:�� `#�G�>��{��T����b����k���q�1H	�\����iJ�u6��q��]�[���f�����u�j��������kg����͏͟)��͓ەN�b�
���ͤA1  -�kc��V������Hf}����LQ!.�]Bj��bWRi��Q���!"G��(}MT�������;������u�1�N[��u�<>o����]q}z�4�C""�5<ڽ�n����`�������!"""��P��܏�_Dsc1b�41@c���/�X�ND^ൃG�N;�����u�c��U��9���O����U�<sέ�+�։�d')<t�}Zd�?�k�]�M%"""�!�I�0�^\�B%��q��� "��D�nˊ��H
q��ݔ����@��Y-{�ȉ�ܙ6�NR�V��c�.�l)CDDD$/uF�>�;"6�.!H�rx;G=ܛ���$��-��gJ�l.�o�yLq��ui)x��1�e[�r�b4B��^[��`w""�	�〩�B�|\�[��P��o����J�׈R�F����f�H��ID����ٜ��I=��S�l������+�R��H~�4j�e�.|�I��d�' ���}��j��x]�+܉���~!������{��|JR��e;���&p�&��HvD�r��+��^��]�����A�7�Bjt<LM9o㰇���DԿ+,�9r��@�F�D�W�FcK�ղ�Ŷ[��4O���Q�3""o'���|�&oP����}��]�Tz�'``5?�Ɂ��]
��ЛLhlQ�� ��YP��i�]c�M-}7i�Veq��Va��Z� ��6������5H���J�[ՍMȫ���lB|L�>�����E�V�N��/��lɎ�,�
�5]ܽ)�V�z6"""���F1�ߏ1\�<C}��碰󕈨�ʭ��[==0,��?52�f��QZ��`0�~3xlND乪tM��J�t.���ZʘX�NDDDDDD=�����|�B������6��57_n���FV��NAu(�ա������.p'"����C�*���� t�!�v�������*��&#��H^.U1p�ʪ�r7��+��Z.oz�DDD$s�>&̉7b_�:������:�&j(�- "�D�mK|HP�<~T@��ee:]���i�^K""�\��f�mOs�bI���u�
6�#"�x�%9��u�ϨQ���jT�`R��(3/k��.,D�.P�b���s�R�X�6
!�>��V��Q#�G_�>j���+�ֻ>A>Z���w��-]����!�G���$=1��Gv��H����'"r���z�����z���r��k������7m{����ܙA�'	(����=�MA�MX"O�~7m`�	���<]jiB`�D�����9��Cp����O#�3p'���^K�J�+�`?p7{��K_<&u�٢
T74!���J�/�q>�K�U_^��w>���`K""��^�Dm��EīK`*]��C�:x*b���}���}���DD�QI��
����.8
�}Pm�
w""�i1����Q)�V�
�P\S����J����<�ˈ�r�� vkRT��egc�f"����V�;��#��	�i� "�Ꚛm���]�TviYOa�ND$O��xu��剬.�׫z��L&���;yn�P0q'j�tbk�l��>�9q0c�ЗL�\����KS���k��B��Z�8
Ճ}z�k䠩DD�������ͳ�Q�}v�\���u�"ty6��!j�P8TD����/��l(F�NG��/�Bg�[���p'���^���K�������_{���DD����kN^��q��6{�p�����o���-�u
w""��`!QE"	�f�,3���0%�/.u�G�a�;�_�Z�4�[z��+쏑��R��;�ze����uw��+�Jo	��(CD$<0#j�ʞ�J�D@�IBXD��Ġ/�:���e�;�_~����t��^y�ʆ�˂�"pgK""�:|���05�o[V�&Q��թ�Z�����9�o(���������Ug��Z�A����x�FG!Q={����E����D$?�>�O*����ۮp��h�d��AS����Ok�b����-�ڰ��'������hT�zitx""�̈�t�r���I:�pW�4�t�!��ӢQo@s��z4��6v�%D�����
z��M�÷W�\$�T��p�j���N�c�њ
�(��ټ�J�@��/��\:���A�������V���F��Uc�Z�Є���8x~D�(��vyo�*l���}�`䕋DDr��B֟�������X��G3���
�E���BD���"Gz#pg�O2�٠���������w��2�p��X<8{��e�&=*u��T^�CAu
�j����6��)���{�X�{u�q�r�v���ń�h|������GR��^�����`��_��=oeq��/��	���Cay%~���8-2�N6�������I'	�q��/o;�U�3�i%2��9����W�\Y�����C��a��gED�~�j;f�����g�J���sw\��:h������2�gS�����AS�]8?l!cr0�޼�������S|X����%�|:�n��ґ��.9��\����\>��oN�����X.*�۳���'F#2�r��ؤG���z
��<�55#�����a�����1o� �����L^�^�]��I���v;����������p'"�?qU�S��˦��zn��+����p^U��We{��""Y�QG;i���i�)OZT��}gL��ٗu	�2r��l�J+�~qz��<ѲfBR��ީ��z�AV����{�
u]s��5�_��fǁ���2�샍xz��ǱE������oDRx�˪@�͆D���	6������Uy'�Jl.����pDD���ۏ`nj�yJDs4�Y��m�k�p���]�
w""�m5�H&��i4j!7"wQ)��� �ߛb�,���3F����`�˖�Lq*pf��WmY!��Jѷ=����M���T�����wr^��#�p2�?[<ғ��0��̋����6J+��3$2��#E=�/,�;h�Ԥx����DD��8���6`�OoGT�?�1�ѽ�C�� wi�p��Q����Cw""�fR�����, yp�/�Z�� {�&�������q�뫥�S]�t�`�ˮ��߯�m5_��	�^�����[�tl���X�klw� X�7u��E���o����'���m�G�-ەy+�� YK	GT` J��L�/�=F��c��γ9_�OJ�C_0�Q�QR�Ê׾Ě�o�������W�u���R�[^+�l�z�<0�H��\��S;c2�e����_}���]Xv�������0>)ߟ5N�@���H�*,�����~�\��>	�q�RF��*�F���uqoXT������]j"������D|z�ղ��.��co�α9rb�Ǎ��`!�,��+��o޽�j�SN�>�C�ױ�|���-}��F��;.`u;yn�0�z�Hm,
��3�92�3��{���8�Wl������u��/)<#b#�?����V:�����(�k��8%��;�����.[�X��q�z\���R^�C��6;y����|yΕU �0�mjƺ�,��n5DDD���|�����]�d�����6b��Y��+�g�Y��Q2t'"�l&w"�(=����5ɯ�]DLK���V�5�R�~$��?������0�ru���B����c��uS�I����6췸_�Z��Z��ol��@Wu����[i�����.J�N9�t�<��z��ܽu���p��s�ɳVW�����Q�@DD�N�����	�ܱ�v�#�f�T�/N���AS�w*�u�ȏa;��T���&�iFT�Y��S?���E#K���ظ���������M-�55�G�'���e.�]������b�z"#�C�^�a׎{�A�~m��ua<���l)C����0�<[�r���~�~?64*��x����sDB����������Y�ᥕx��e��+���o�Ƒ�%=�8���7�1�%x�k%"�H�/q�P��׌�M�9��pZ���#9H�������c��'�G�Ƀb�����ჰ�L����$D\= }����p��M--�e��ve���� U�B�,O�t�j5tx�����l^o}�w˟Y�BԹ�&���������i��X�
�������i ""�)s�0��⵻ajr���m�������{J렩ސl�� ��������S�QQ߈J]#*t������'[��I���$�pԺC���tQ)m�a��L>9tF��Z��6��Y��%�V��5$��zU�z����'���b�����l�e�.�����
�o�7&!
��B��e;!�]m�h��_���]z��*ܹ	%��-#�!:0 �u�V�~�q;n���s����W��y2stl������'T���W�g&��'Z�7ԗj��{�ڞ�v������v"��s$���&J!R� Ixn�ad�^��
V��q��=�½���*KP^]
��
��2�ٻ��ہ��
�>v����KK��YT��8z���NL�A\H�t�Ҫ���b;��	i��{�
���j��[�}�C����9�]{�;ދ'-�:�Q�g�Ͼ�ZV�k���|��߹��]?y*��}�{r�m.��u�x����z�h���ʼ���-s0���G}A����h&�r�4�Roj�p���`�8A����<�Wn��:蓖��C��D�m,|5}W�^ר���� Bی`- �a)v�u�[ʈ�tW�MM����钑�������]��Ř�m?�<&_ϒ�:�'
J-~6t�pW���6m�i}P�Ԍ��&�66������)�Dny�����w�AS��s��qx~�!/��:�_�Y/�����B\^�h%��U_᭯��\~��t,f�DQO�(���/~&�T����02.�W_�n<��'���G�-���7�Je>l)CD�w��+�����a�p'���_��O��Nlǰ�f��g2�'����|�>("D���EP��s8�W��� �t�$�0�j��f�}�.n�$}p��b����������΁SRO�V�噢r��`0YV��'����?�wϮ�mwy�_���;�S��-��~!������E��QϾ�?,�������F��:�z�f��O�lDFi��ۈV6Ϛ��������4gh"�9��Z�s��b�����˻�I�_���������ZiJ��5q��j+xP�7���p0jj�o��:ī�t_���_���sS۾�z�"]����������|��o_�o�O��]38�������c�X�>��Km����6R�Z������֪��c���F��M~il)C=eթ���j����_��7>tx�/Z���eMJ�Çw܌2��;޲��rqՉ���m7n=ˆ���X)4o%Ƌ8QT������S8Yd�b/@�����@T��wWI]=����n�U���Ъ�Eo�v�~��]��K��ǳ��7f���<��TL�p��T,9X��uG�.Bv�n�:f��l���s��	�MWFzby;Q�zz������D���KW[4>��ڼ�I��I���d��U�o���,8�u	���5�(F2�u��*S3|�z�Қ�Uڏ�����&wѿ�����b���o��3}t�L3l���E���d�w�L���߀�����qH��l7!&V;/ e�'���8@����Us��zJ��o����$mG=ލ�inyZ8��ux��Q��)��ᅽ��I=��||��Ij��^|t�rLJ��;5��CeC�[ש�륩+<!P!""���5��]ǤI�����Ic0>1C�¬�y�H\q�WQ+��9q�L�O�:�H<�Ӵ�ް�̖2DD���q��#b#�S^-Ue��)�h1Q�"MDt9�n�hԠ��_b�c���@O�`���]^U_���JT�UA�X���Z��P��������̺}xn�A��F}�Ӂ�Ҽ�y���I��H����x��r�]|}�	���$R�b�0i��u:�/q��Ķ��} U���m���UCu�������s}v����k󁎑A�(Ok95%�=��8}u�R�j��m����=���,���s��yZ��'&���WUM��D�4��ը�(��j������>oqm�t��\xM��R�l�C`�ND��D�.&"�\E�_� $l�#H��P�d��B�޽����vtD[��No��;Uk�6���$Ч�$�y7S	u����&ȼ���yx:�7�t���S�����u��4���8�RE�۞C�8�Ѕ���U�'Żm]b�����bVr���+�VV�m�3�������3W�鍮�ӌˉ����}��
����&��&"�D��>��Ď�Q�w�t�&z�
��]���s�xo:�'��ANe�ÅQ1Q����X1:=y!wK?�p'""�)^��J�I�B��������Hv�F���)�|�Vw��\�9j7��F_������������P��Je~��q�ı�~!��f⫳�YV���&&�bQj�y�ɉ�荎�b`��N�����+����͛w��!"""""�`S���[hTJ,�,M�^�Pj�u���U�4���"%"�!!R��ޖ�o�DDD�9��9h*y� �Fj#&"""����]$�&����֖2��5QQ�K��*�vX!""""""""""7��]�T�����9D��x�Q?�5�{��v�\DDDDDDDDDD�v^����Qj��I�~�t�ĝi;�]k��`�ѿ����DDDDDDDDDD�n
�	�
�DDDDDDDDDDD=D
܍Fc�?��!"O�my,��_g|�/"�4�U+�7�P�܂��&4x��������Ȟ�
�~���;�cj��ą`F\0���C����g�uX�[��f��������Rk�C�����;��"�Q^߈��f�1,CC���V�P`td ����P��Н��.{}�I�?�"GT*%}4�G�K@DD���������
���DDDWD�_�ga�����M-T�P��]��<5�A߂�&��\o0��];��b�p��
�
�p��ƶɈ��}|8DDDDt%p���l)CDD�%�1n(�z�t������Q���銚�f)H������gqM=�;��w�@Y]����������777{�h܉�ȫ�j�o����-�7��-3��
p�R)�J�PTcy�[T�?�a\� LI����D���H�D��O��׌����='��w"""""��IƄB��:���j���U�F��#
�Ң�(}�|<�]^��}Â�
?��58[Ta���Qq�U+a0�P����vWZ����������;y���^5d@޻�:�F���;c�!y~�q|~�j�h����`n1^�s�������;$Q�������34|�	�W����=4g<�v2���ѤoA^y��-ā����Gqu��m�����I��ԑ�R���P^^�q�?/�-�����	Q�����S��R���_<��Z��`DQM=2K+q0�/�8"]��]R�����ϙL��*~�\DD�UF�E`�w�!2�򀨗�����=Xu"�˕�b�d��\i���?-��iɱҲ�#����WWKUDDDDDD$_=��w��h�3{�U�HNJj,�vq���o����������W�'�l��̋m˞�~�?{������G�� m nxi%��m�;�|^E�TY/��E����&ań4,~�S)�����t�hx�DD�5��;1_<x}[��ugr��7��ҹCy�X���j:��l��;XS�c��p�lV%��V����>Ó����A�6o�QX��^Y��Z��2�R���Y����|#w�>�gf��{_���l��l6ɒ)$��H�(�������?��w�@ !!�����I6�[�7ۻ�޻�.��;^ے�ʖdi���K�6imy��|�a{ek�����N�[�ZP��kEMGo@�����O��6��u��gb٦��l2@�d$�Zp��w�s�ֵ���>��w,���\�����K2R��[7�?��P�|>�{v��
�9Y�gB�z""�!�r��
�����=�VDpQ)�����]ӌ�|�:�&���J��+�W��������.~��:pۯ�DEn:6�.��n�8t�8��~ḭ]��Xs>���_�m�a��q{�����%C����˟B�z�*�x�m�����(���8���ux��;��(�~a��/�2�{��f��P/7#�I�d7�L5��,E϶��=��p�f�&j�Ee���|;�����p�o��K��	�ғ�+��C�8��	""""""�"x���Auk׸��Ph�a<��PЯ�� kh^R��I"d�@Һ��l�2���ܲ߻~�����,)��k��b�tmmm'�f�~I�\��Q�#��%ix%��D��C���z��=���N�><�SWI9�:fu^42��(RQ�'�֮��:�����w���-VI}��~�I}��ϥ�=h��H�A��8��M,���-~Aa�~����0���{A���;ԋQ�&�s������ns�����u�����Wo3���NJV/Ũ��.�����y��<_�o������n����U�Շ<�<���کy��e#���gADDDDDD�cd=���Ό�X�F�<3u���G�'�Z�V�i���h�m������8m�}>x��w�Wtd�.�r��P�.�	��Dnݑ���3��(�&�i�d�'I,H����Wx]�������냗Jp_̢�7D ~��uk����m��O�:�m��=�����s������l���ψ������l^^8�豦�I��g{�~����s�����Ճ#����+���l�ϕ���]Ϩ�G�z���U�M3-�S�I�(Q���(B>�t6������v<shr�Ჿ����KO�=�.b�NDDDDDG<#z������ow*8=m`���s8q��>�G>q=6Uݞ������م��{�WvbdK��*�S�pӒٸy���j:zp�yrF�^��OTQ��-�#""�F��b����	j �H�0�q��Qܯ[P��d��ކ���c1�q��2�g���j�NӮ��Q,��iwy0q&� ��@��Q��������ŗ�\���yL~�������xyg���_&�b�._��+�r1����v�<���j����f��Ϙ~$ADD�����yQ5�ԡ���K�A�����r�<1�
6�.��O���.l~^&��u�M������u��[����(�F���n�!wV�eT+�`_�g����N�YI�K4�7]E���r�*<w�
��[�|��J�i��5M��cxl�q�Jw�wx��yQ&��B��lš���0�u��γM�;��.Iz�ꛆ�o(g�ND�$�aT�.���߼~=�7�c{e�����j�G�����'���K���^8�2{��/����
�,ia�'�.�W��e������mx��9�e�	�����d��_va��$9�i����P~r����M�&��n���[=+DDta���;*l����s�Qԍ�p�h���g�cw"�dЮhż�wA9���`ۡ��l�"�(D����}{u=~���n@�́H�܋1Ȳ|F��""�8�y~�T��5���Ce�%Tut��rà�i=܉�hb�ӆ-��k2��jݪ1�hԃ���(�F�p����aS��u��|�v}�b\��o����=~��Aˋr�����v�h��V��o�y^Y��쬡���8�[���m�n�?��A$i������D<Q�܉�(Ne$���O�u!�D��� �o�Bin&�MFE�-ODDc�!��6�]���׾�C��������-�n�=n���<.�^7$�C������޲�5�9^���n�Wѫ��1�}������Eɧ�<����.Xn��� "�����"'�gbMY֔�����}-���賡���������C������`���I����Q�g���EU[7��}���Nu���k:z���q�rܬ>wPg���[������5+Q�?|F��@ݿ���m@�`h��$I3f�{�^?3�,ь$F\T�
w	F�==Z�.6����0""-��,�ڼ�q��~��o�����.[�T���wv���=���v��{���hU�3�&çn�ԯ���tх-+�ŏ�
9�o�'k� �N����[�,������]V��g���s��{���y�=<�����l�f1�����i����s�>�iבq�q:��4�X,�e9DDDq*#a������m�L?���߶��yޠ�J��h,k2+��������?�ި~�z!�]�2�@D����̓�Ѱ����<"�9p�	���/XQ�����P����́�2N�;��=�618醟�_�j%�Z�@�u�x�H��zf��ƀ��iF}wr�,���b��T�QkGӠ޾��n;�����^S����ns�^�pl)Ӈ@Q���DDDq*�4P��P7l�},]�/��&�""
$��9��U�+�Q�␩��u'�]8DDta.�;��i$��ju�^�k ��7�ֿ��6��K�Q�����-4mdF�:��}}��}�c�b:�ڃ@��U��p'"��e�T���"����o(u[mC7��DD�\�߃��I;ġ�~S�v���tL�V?�ߩ��U�*^���[b� >Y�G������`�Y�-��b���j��5nc��h�z*�_$ ��M�O���]�כADDǌ��@��~�9���ep���H��>�_��a�L�b0BgI�>1���y�� ��]���e OqG�k5$hg�9N8��`��n[?|�)��}�"$�|/���B$��鑤��Y&�r�^�?�Ni�{\���3�{~�C[��u���2��IQ���dP��<��hR��+�Mz�����w�U���t�}W{�mrtu���%,f,�~����`���۫3C�Q�{{���_X~��3!��"Z�ܴx6n]V������xl�qP|Ѷ�L&S�$Io#�x�ޠFVS��{���8�RR��JIꔃ�2@����x�����m��|�:/[��T�2C̫S��i2b@_��S��V'�:�dY֫�Ɖ�e�:ec�L"��x>����������(���DD~�აƔtx\Ρ��]�T�&(zd�^��P�-�0��0��	F�:���]�n�3��D��dug?/��l��8����¡��8�V���'�����:y].,��vi�Io Q���Ϋq۲9Cׯ�W�9���/n�mo\��7ʲ�(�}>��S&���l2���&�s�ͻ05����(Hl�V�<�ڃyq6 �*�' R����m�w�x�Ӫ˭.��{>z]����9R��NgPV̲v@CN?u������K"��F���R/�|��������Z���ҟjP�&�3Šw��t�T������|G�10�� N,�o@7���g���;��v��lpPRQ�.�'�Q9u�[����uDDS��uނáyP���N�t����7H�͎$qML�>�Ð�3;���h:,+��}q�2<���5����_q�o�+A3J�W������4��޲f�q�A?b�vE��V���p%��q�����v�k[z�9��5-��g7�� "��|N��+-����W �݉�"inN�����3p�#�?ߜ.
�8�z�>�[%�	�%���s�P�j6D5p�v6�#o"""���-w��&�m�0p'�Hk���\�c]���N��0�DD	6���r�و������`���Ȟ�DDc�ڭ�W��M��B �DD���Lڭ6d$�n'��}�v����N$�4������$å3F���+��冷��]�Ex w��S<Nm��$�&g�iL@41p�`���,K�Q�}"�a���T���;����<t[�=ڝȈ�b��6�s���P��jX7"�)�U�����-�ݝ�h�
�:z��WvboMS�c�Nr�N"��d���4�7��EgF����;e�M�^����������j�ne�� ��)��w�sg��H�����$���D��?��9Y�ND��ܡ*�h~kK�p���j�G=&��u�!{#\ǌ�^�:��M'PS��	�N�)Xcf��SDD���g�ZR�������|����C���;���F��ĝh���ܹ�BD��Ts�6�$گ�:�i�u��0��Pq�4,DKNŴ�.w
�O�$WE'G��W��E�DD��Z���S��˒������]���ԕ�h&�o'#D}��h���%Y�ND�${�(�܁��VPxI�w}~�aV�-��>~w
�"��u���h
S���%Ѡʶ����d�IVd��φ,���l�h'CDQ!��k���#vrAD4���߅��9�U�(ڭ+^��:��Spdy̟)�w�XDD4�ds�VE.��TQ�u��֊�̡�;�6����F���hD�nTd���D4���PY����$��,\3���G�u�SPd��c�Qw�^�NDD�D��^]+֔�bQ^&�R��mE4��2f�]��DD4@�FnF3p'�n���M���h�ha��w����>y'�4%�3� R/��2u�`̟Y��	wM��m?Ӡ�H����G���z��_��i��=V�W�~�DDC���k��M?�烤���v���G�h����OI�.$2l�
��5!NCdڰ�/
E��]�y�Q�yd�	�w�2(���]����atۦ �Ĥ$�&k��;	���\�S20�}}�|�-e��B1��{r�������j���@ѡx\�uv*+6D��w
�Q�>z' *܉�(Й�<w��,.G�ɀy�
|��ӾEy9ڥ����0�`���o_�v�'*mAD�Mg2���%%DD�&k.�ډ��om����n�DKNEؗ����"I�1�j���!�}�""�o��K`P|����Zـ�������X^���X�������A ""
�d���f-ѴS�F�R��Q��V��1$��(zRr`7%�u��)$2��W�K>��!"�Xc~��>|����r���������%�}iy>��ka�)����O��""MW��������(*$�A�ԫ��DD4���>��m�):|>�W������]$� "�Q����rN!6��#�l�s�ވ?�2ޭn��k~r����V�{��;] "���W���s��8܉�A� �,�嗁��f���2�SP$I������<�:��DDc�x}��O/�O݀��9H4�̽7�[�'������D���66�����?����ZADDc��fW^����EK%�N��� �'#"��t���1p�����Jc����""O�݉��E<~�uXW���3���V����7���UZ0?U�	�w�%���E0�6+z�׼�7����Č��W�!�E�l���j3��.���(�O��E�<�������z����N��E�%�}�gϾF8�SO������2^K����vфD ���>�o]�_ڴ��}>/7���f|�m5���)<��4����D36�)��KթX��j��]��ӭ] "��tz$�|/��y��3U,�;!��{��"�b�#3��2�9�.A{/搖�h��S�unV�S������b���=܉�.������؍�O���ׯÊY���e�������n��pc;�7u��ώn�C}�O���l�cvf�kϑG�}�������p�y,��h2��t�Id�;�t�̡�VDD�MGZ.�F�&��z��H3=�z�nD���="�`m�n��~�nXP��o\�5%yC�Z	fl�]�M�j���='��G��mM�ؠ��.'ź�ګ+V�9�p�⛑�_K,1p���<�~�N}��e��p'"��x��m*�H�mK+�qv>Ve�b�_��g�{�Ve�<Y�W�ׄu�U"�K��������"/VjW��Z����������z��#pw�b ��M����>m��+�SQ����d�-&�1�v�.������g������w'����6,�Rf���V�SplN�#i��G����?��(�>���������(�H����Ex�*��)(]�.{v��Q�{hC	����@DDDDt��XeKDDD������[	���7�-e�Sp�{��9�ɣn��쩈��� """"��J,�"����
�𮃏�;EIe{�rEyި�G����#""""��I��HDDD&�!����ñ��[��6w
ʎ�ִ{V��C#��?�]�'��r�#"""�J�F-]�� L��0-,B|/�og�NA�q�e����+��|��.��V��z��
w""""��q������!���=6�XX+�)��_������kV^�^5��N� �]�E���D���="�����]�c%p��`#��3p�Iy�ȹUn�o[����"""
�,���I�D�X�NDDD�K>y{X�K���>��?V�����{N����j�_R�����.�����܃ם��=�������z¹>6�g!��hRJ2S��`��sM�I�:wX��MNr�����߷��fI��=_"""�i#�<Zۭhk�������N'�b�#5Մ��$&���ȱ1X����ry����aG�ͭ�AQ$$X�KV�		�q�1Yh)#1p�)y�T�ruŖ�l^P���$<��$�Է��8�~�U��g'\ޜ�t\3���r�vLsO?�U�c�:y�D��U�q���h��Gk_?��lh��Cmg/�v���=� �M�و[�T��+���N�m�²�D�}�Z���[mڥx���e]W/�����#X?��r\�����[��� ���;ap����B��N�5����,����p�d�RM(/KGNVB��\��g�u���o�}��n�v�x�x/e���β ��}�/��1p'""�#�K��o7m��O6����$��9�P������Q�'���;6�������i�Ə_ۍ���u_v������=v'ޫk�ן~'�;	�,��B-d�i�l���<�<������{����k�����G�֩�qPk��,.��?�v!�u7�hf�;�Te��t��>l��c��-pw��Y��:���V���]�%��iW�&-pw:Cl�)s�T"""��8.*�Ǔ���=��E�xp�{�Yz���1/7}�6��U�msLv�vyâ2�������/4U߿xs/�7�c�|f�-��8��r�#�߼��^	V������Xɡ�1����n�u��;�-�j�n_�k��߽v~��^�<��N4�H܉�����l����T5���ٴ���N��H-��!�C$����M����H0k�+Jr��������uZ��ܡ*|�w�ms������ڝ��WCu[�v}˩Z�n��/n�B���`B���1b�sD��On�\�=����i����_���'k��9�u��3�:_������P��XJ�.4����&�ߋ�=A�t�٨].��u�`�hqr��?y}r�MW�ʺ��}�û��׬��Τ�#����v("����2Sq��uJa������M��a�N4�Dw�h���%DD3M%""�	��2���W>�Z���Q�=��0>�v�֣\��K�q������LFQZҘ�{�W�G���_�Zʜ_��_��v|�����wߛԀ������eڼ88Q���Ϳo^	2͓�̉�"��=""""�V��D�+�mΉ���;�h�^����n���{q~x~����bg�G���}'�^��Y�����Ӯ�C����Vj�
i��	������p7����pӒ���㯍����|��_�օ�?~T;H���7`~nnYR����p'"""�~Y	�2���_������Ǫ��߭��`�W7�Ү������q�����o��'��v~qە�fA�֚F�*1��h�t�p���R��������ϼ���=>��E`��5��?�<���?�ލ?���߼Qk+���h��ւ���hڹ�	7�DDDq��ٕ	�
w�7������}Z��h/#l�W�w��O�ԟ_��ʺ1���YQ!/��~���j���$l�]�^��sd����R&|������s��4O�4#I&~��͘����_������T�'�C���I�.��D]������"���(J��GD4��&e�}�܉����/�6��?5n�zko���{h��Wׂ��yfg�j�e%��ħޏ�|۪�/�N��8���ꚇ�����U���kqŜYx�h5"�?Ò�h5t���C����g�j$~v�&�JOƿ\�G��⑱�ߍ�ʆ�|�
-��t�i弡�oP�����[��<�K\���þ\�DDDq����O1�|�I���0PQ���w�e�m�e?�����K��!Z̬�����yt�q|��G�����e��!p�̠�c���Î�}���~fc�b5������l�6����;���
w""��g7%�5{6�Z*A�לS8h*M�Ư�HEn����M�Qw��%���]n��3�`���C���^�C�u�Q��7Wz�N|繭c������]����H��|��!�j��ǣ��ዛ��"+M�������,+����\��y��dіID��DDD3�����p�Mȫ?����t�g�!�ő�n�Vq.z��oA)���w���8y)�C��4Nj���Du[7���&���¼�q+��.�c��9�	�c�@��z%��J�����lG�v)�-�c�p��Ҁ�o���z⧘�������X����?�:
"�s�"��"��ל;^�oA�a�{h��gKWE��]`�NDDG�>N5w���,g�೗/ǯ��xL^�p��lä_C�)��<����C�s�|��o]i>~���H6��}����4U�����9i)�9]�}�
�	��%7i�,�g����y��e�݉O?�
^;~v�>�7_�*>+A�qg�N4���LҚ3E��sԭ ���ū~�ճ��iL@�0p'""�3|� ~�����7oX��e��VY�UK��IǦ�����Z;G�p!�=#�d�Š�Y�C�٨�E�����klǟww=��,�vA�V�^������0oD��GwG�-/��]���W���#�2�j�%x߼b�p�����A
�	\�d��u�ݎ��k���d_شK
���N���F=��Ƞ΋P_|nb���e����H0cqA��r���ַ�/h|��ƿ�x)>�q)6Vi�#OD��DDD3OGf	<z#��wC�N�ȇ&ϭ走�ߒ��a�NDDg���8
ӓ��ͫ�1���_�M���k�g�Ǩ犊l�"�+W���˾�f���'0��ų�i,��ͯ�9�߾{�V�����-�~q @�b:�ډ�o;����9h'�M��)J�uQ���[�����e��#��|��7�橚Q�]^Q�ǋ;zaT����o?�����ۮ�<��iQ��8h*Q��w����;%O�˪v@��A��4XP]�A�6��š���/��]�aqa6R-Ft��q��/��['΍�\�K\L�)�4�H�������Ѫ�߭�s0TA��y�h5lN7zN-��S/ۭv4�X�64U�]���8�֭�`q���W��N�V�]6;�z���hT'1�H�}V��n�u�J݇���ms��~�e�v�`mi�vpB��W{�'��DCw�"��?��~��|/��9�}^�,�`�N�X�NDD4s�%e���2�Un���3[��nJBU���iy=�DDDq�hC+���-S~�z����z�O����Ԧh�[ӤMSe�;��ېl6��jՂ��<ޡ��������7��o�n��NQ�c�;ь֟��ʹQ~�]�]vPx�'�kg�uL��;�6�S�"a2a���>�(�1p'""���dT�݈�S[apr Tݩy8[�>Y�tb�NDDDDDDD3�uQ��Q9wJ�wA	s��W��/���$���5t]�y�ۼC�e�3��I�ù���E����;Q�p�85o��uH�m��ާ]���Z[��Q�Iz�v!�w�ȁ����"���2�z3l�X3�4&h���ۼQ:���;Q�ArVK%r�C��A҉��m�/1�����O'�DDD4JiF�6h�D�L$h����h���ɘm=��K�kC⩭�K�BM�
8��3p'""�czE�¼L���py��j�BS�u���d_�j���M��O���Z&�E(��� Ei�p����۪`w�_���$��I�;�msh��s���o׮O�Q����!�bu�Š�AQ`u�p��DD�4�i"�.��˘�fK_;ʪvB��~���ۊ�G_G]�Rt�Ϛ��f�NDD�Dh��+W��/��v�m�x�H���6?��y�XW�?��E+���-B�k�Ǽ_�߹n>}�b�t�=m.7�v?}}z��QϽ}��yci��ǻUuxx�1�}�6���D|^}�￤\���I�g��Vl��� """""����T�����C��/>�F{��L��2p'""�3"l��Ǯ���Ƽ?�b���K��0��9�'���;\Z)�+HMԪ�]��X���Y����FRd	�赸��_}~'��g`yA���b�D��}��cSEn�ݳh�����[.$���N��֥s����UZ�x� *���V��������p�������x����'"""""����v����x:�uE��+�g61p'""�37^R���iU��Z�f���צ��i�iA�D��;K�E[����_5�X�,P3��������ub��d��,*���Z���$,.�nވ{}%���<�T���j�4�	�	�^f&������J���.�ۋ��_�ً�����n��?o\�UŹ�}�ܲ���>�؝���m-����zDe&{�*�3l��̖*x�/���ň4�DDDqf}Y���ܴx�V���.��f$�Q���͋����r�?>�7�h��իVi�M����=���4�:ro�{=�d�K�h�y]W���Y�O1��7p������E��� ��2�}/����Ok���-�m�����~�DDDDD}:�e��C�����R	���֜�}�DDDqf�Ŋh����7�G������TE��������`D��Aˋw�Ap�h�"�����c>�W]�ｺ��}�v`@�����C��w���4/g`=�ky��9�������������O����v��4}���nJDoJn�^��;Q����MEX-���ڵ�8��~�m�щ�e��g$�����䪓�0"p�j����=�֙���K�3w�~x�$�XA/Td�a��1G�p!�_����=Q$I�~Ii�.X��@�K���݋���`A$0p'""�3���'y}�:�ŋp��B������{�5���T�qh~mIn^2[� ���~����)� w��Ks����A	�����I������2�D/��>z��c^x�p%.Ŀb��D��Ý(*8�M7	>�:�I=͠�P�N�T��鹗��m0��;Qz�T������Mq����D��[�g���������^X[��M1�+ܳ�C����q��a�\��hזi���~Q�˒
|��K��!�<�T��A��{��p'""""�����3���Q�.���M'ќ7/��f�NDD��ۺ��?�����߀99�0(
~z�&����ן~{T_w��u1�h�_h.�q1�d	�Ɓ`�7AY�D��Y~���\�_@~��R\��T{���2l���Hze����w"""""���i5�ؐ�x=�����N܉����'�a��Z|r�%Z?w1���_�$�����p�U}ۜ�y�W]��#�0;��m�������?4h��ۙ	�-j�u���?�+��p�Y�F�^o���U����y�DDD�휈hqw$����aBo+w"""�<b��T_=~�~��%ia�����ͽC�k��]o춎�����Zp-K��� �Xc;���:Q���4<8��ma�������C_�
�5�����6�Z��W��;*���#mw�ADDDDDD$(gؗ�����h9�ލ7N��'�.Ү��*�l��o��s�G�J/�H�kD����x�%���D�{q�@vܿp�:���~��^��vAj�?>�+W.Ղ���r��8Ǜ�/���mw�[�.�"�M?���,�DDD3�s��]���M�T���[����ܟ>X��ݰ	�	[ʔ�%i��;����`�lG�viw{�gJ���BR�J&�u7�y�����-���H�]���w�������%�C��%�(.J�M�}�N	�E�֝u�E���4�K�BZ�֝5!���ρ�;Q�Y߹vV�䡶�Um�8�ҁ�͝�n�҂�5�}7/��=��φ�G�A�;�����s��3~��L#nZ<�~-h�>��i���+��������p���U��=?��'��r�Ͼ3j��Z��Ăb.�4ྟ����Rq��C����6m99�э�~;�,&V�Q �p'���Ѩ����Ѡ@�W�����;�C�p�ś��Û.�?��ER�w?�- 饣��{��-e�gU�?>�m}�Q�=��(*����˗aUQ֘��w��^5`����^��^��;�>Q}/z5t�qQ9nYZ����D����3�g2� Q�`�GDDD�-��hf[?��NDDD��x?c/�ݰ���k��u���/ڷ�x��ܲ/�Պ�'�������A�rީ�7�����Şs����Vca^���"0�t�V�~��u��J�׎�C�a� ������Onل��.�`�.<��0>�b>:� """""�XIR8b�X����^B��DDD18�`��N�Y�����]ޘa�����￴K
�ǽ��CUڔ���YiIZK���Nt�.z��ͽP�$�X�W��^9Ok1S��5����6�m��
w"�U���$""����_��m�x/���e2p'""�s�G�&�w���cԶ�Xc�'��G�z!���^�/�����z��/l���@DDD�.�"�IG���� ��;MѶ%���]�`��Ql��]N"""�u�h�q{l��w"""""""""��Q�Qw8B���5RL��	����;�L1�M�,�+��R������(qי������p)FF^��D��;��(s��1$Ԋ)�2p'"""""��X�����"���aX���p�2B|/>IF�1p'"""""""""��pT���S�.ˡ�ݡV��"�a0p'"""""""""�0b#,�b��L�+�}��pc�NDDDDDe���KDDD�#�#pq������m6���`w��@]���h�#-͌�LL��X��������AK�m����\p8<��|��$���bBvV�:ozN��^V�]|�1f�`H���DՙN44���{�]�v�5�����,f��!5ńX���g�C]��9��ͅ�;�zq�T+2��{IGf�%�;+܉������M%""��t�@���6T���s|hj�jSɬx����!���)�^:��� ��ѯM��Ip��!�+܉������Rl��Q�c��}����+Su����б�sQ�*�p'"""""""""��B	�cM������n܉��������DDDq��c�[և}��i�,=��.Q�$[<�0�>H�i�~x�F|�٭�s8ADDDDD���7""�xǿ��ǣ��E��4|x�|<u��>]"""""
]�C�є0�"�i$I��k�^��4I^5��尺4��;Q�|<�sX�NQw��2�rUI���������(8>I�&���kb�KgDOJnؗ�����j6bvv�6��8�,���Qȸ�MDD�<�5��0�z$�����Y��ֱ�hnn[M%XY���M��es����������u��W���J�(j͙����,��;� 51����ञ���7��S """"""""����
!���uf+ݣ�79�"�|���1�����X�FDD4�t�ς�@�;C�icMHÙ�5�Ir�^��;ͨSBz~��"""""""""��!{�(:�(��d��� ��H��;͠����S{�	����"""""M�^6ьԑY�]2t�,�)	Us6���#�Z�)hF�p���o���> """"""���8Q��]�$����=D�~z�ep�M��z�)h�߯���؉��������¢=�Xӥ���ae�����2�u�i{M�4%܉�������x���MPT�xN�l�TTUl�ְ]`�NS��xADDDDDDDDD�ӞU:�^��0t��~K*�E�i��@�����v���<�$��= ���������(��2K��d$��a&��:xey��^Y$e��nEI�Ǽ�79����c�NA{��m"""""�0cK""":���Cf�Hީ�t!�OVi��#{\�/G�d�s���{�����+��p�nJBwj�I�Q��DDDDDDDDDD1�ഡ�Ի�%�KL���ڔW�i�h(�N�y�ׅ�;M��D���eADm�U{ yܠ�B�G7��Y7�J��e�YkWB
l)9 ��Z���hf�;�Q~���![U��uH�nBm�Jt��O��3p��]�|>}�*m��w���G��+�N�I����@m{w���F|��uHO2����(��+'<U�(\z�*��-e���f4�ˎ٧��Ȱ=lD���]h̟�������)h	
�S��ճ��wQ�����"�b���6��ߏk�_�a��L3��_��W/����NDD4��b���b�uQлa��

7��C�3Ӂ�;Mɂ�����t-l��ҠSd%�qmQ���m�82's����hFa�.Q�|L����f$�ہ�[a���"'������P�8�����������3��6,.��ݠS0+3+}CEm�@�X�DDD3{RM�v""�G�vb��wa���"/���ϋ�YK0�8T�����l^~v���%�rn���@!��(��z�r����������P<.��~&[7h�d�V�+I�/Z��`�NS6�0Gܗ�U�٩з����aAi�6�����h���~�I`�;�L!���S[a��M���*�$9b=��S�F���W���D3�2Rn/�JEK[�6��_0t��}n""""""""���[�lg�]���h�S[��0
1p�)�W��EE�������r��*����ng�;���z]��I�2Q�����z	�NP������`Fc���.��;m�NsnJ._P6�qi�7%᮫��9h*�ÿ�D��CTDDD�N��`� �����[tw
��K�y�G���۸�MDD4��?�:�""��"�����Bb�)A?��DDD3��Q�"p���;M��]��;0����T}I��`E��L����q�5F�.����������Q|�h�(x��!""����w���v֦X� 3	&E������x/����S�a�ɘ�>�N��kj���K��3��_lO_<]���z�~+�br���t��rjS�����7h�l2C�$B6'B�)iP�i(���H��:�t
�:�dI��KP��)����p����O����W�1+c�;j���;Q,��v""""���(KGQAJH�ص��~'���4�E�!-c����)?�-e����Ue(KM@�|�݅�]���xs�� }-M���b���æM޾�Qw�,�X�z5>x�&�&!ŠC�I���1�����S�7#"""�<�'""�3���C�Rb�.�hԅ�^BM�}���S�q�c3�6*2r�ڤ)H�-��O�
�݁����dm#�4�����==��lp������О�s���Wk�.�����6��\��ݦ�����	��/�
d�^[��hR�,�0[,HINFFZ
r3Ұ���υ,��7:M���D��x�9#���D![?�nC�b���,�c{���I���D�G0�cbM�Ɉ�.��M;$E���M��ǂ]""""��
��\�l��B}/��Nі`��{7�GC��?;�������aIa����nU=����8X�:m�x1��8�/Qhx��h2�gǗ���"'�6�c���ew,��4�	�.���+�Ǔ���� �W͝������ۧk�e�S�L~�\""
��g""""������:5��2u^1O��~Q�:�@�o�^���uM@�>H<�ww^��?�3�m���c��p���̞�DD!��(Q��iǗ�""�OM�p�����"&ΈeK���3V������}(;��r£���˖"/%1���=V���(�HAv��X���e�ד�.1�ODtQ��� ��/DDD4��#o��;+�)�dj��
?�2R���ދ�9��+�<VT��62���ʡ�n^R���.*2w"��H�"%""""���B������;�8=eh���O��8�pS�)fc�c��.m�T�jf�%�YZ�W���67D����>�EN�7)Q�X�NDDqHl�JKFIF2���Ku�KN�I��2#�^�'Z����n���׊��Zq��-�R�ل9��(��@j�E�ۅ��V쫪����ȡo�a�Ǝ��t)��T
�Y���H�)h�_��u�㽗��71����w���z�6o����ŀ�-��]O;+�)L$�AQh�=J,nvQ<a�<�/���Y�XY��t�iJ˲�=8\ߊg���j�m
K�m�7�4;+ʋ1� ' �4+3k�⩝�a������=66<�8��a�NAG]�t��n._�
F�~�vq�񾿽�w �6销e8��������D���KD
Kv����f1vߝ�����$#� 2�UŹ�tߦe�l����ϻ�����rsS���Mk��S͘��3����X��c��z��:GT+�{8r��?�|�)h�k��#��?���ׯ�z�m٧��3ȿ�]�]�p��3��-e(L�Ý�(T�"%
&"���h��˗��Wd@�0;+��t�z�
������c�N���3��c�M(�ʀqĺ��p{<HM��0#5l�;XY(&փ�;EQmg/ޮ�Ŧ��1�?Tߊ���'�6�/�W���tpz��B��
w"��k����(n-/�����s3��uE5��o݄/���?�V�>�p����Ɖ�f,))x�Γ�Z��w���5���]��
�`���������N.��	a=`��r�Ӥ�/�Ć��d9���n���s���Ҡ������}�.�4-	�]�pJ�$N12�[״G�G<���[�|}m�"Td��5���>��v����|����ь"� """��sâR<p������%2"��S��$o}�|�����3A?�����8R��ۜN쩬��v��׊p	G+y�6���E[��6X�����Z ��2HM6!;+�pK�Xi)3V?z�Í�>tu���eC��pNv"V,ɏ��ca�N���\���;���VkGm.7�{�{qz큿 ��S����Z�y�5�n�w��f��[�u<P'��z//�A:���[�+P�����!-�����;�8>�� 
�< ���M�=�^�~�1Ɠ���ĻV�y]�z<�����'����ǃz��/p��h��B�͎$��஻N����F�զ�Qأ�.a��9��w��q����=�v��RS��� �2P^���tK̴��ο�ק�g}C7�;m>G���w�`��BJ��ŀ?l?�MI&��{���`�ۋ�����h��b�]\>���3��VhM�&œۗ���7m)zq{���S������uB^'�aᗷ]��ܿ�;y��{�g�[�N-T��K�����p��;NVk�wY�Z;�����P�ۃ�G�Q��=����ݪMy��2��Ⳮ�����V8���(�߷�<�5+
c�)w����#���_nه�&sߞ�D��A����hJ�7�(x���HDD�G�p��ۯ��Qt*��>��6���Sk1�O���y�Z?�}5�>V�"�jj
�O�7�GO�P���ӏ�0�����~��F�"|�DE|��w�a�����*�=!���]���;J����Q�W�ğI�!l�A�Eb�N4��IDD�,#��G>v�6�Y��U�[��i�>�aQ������q����>��E�"X?Z�p�^�a1���?�B���M]��ñ'J�kB}/b0ՐIl)C1LM���9�"1p�03*�?{�G}�}�;�M]�d�W�c���t0��!r�܅�]ʓ<$OrI�r)��rI.�r			9�!�^\(��q�&�V׶�ggT,Y���f�[>o^îfgFki5�����C�@ ���c  ����+�t���խ ȹ�Շ^v�}��ㇼ�	�e��e����;�r��ӆ]�*��:n��X0WuM-��=�u=��[w�SW��w$mޔ�Z<w�{��՛�ʆm=�j�lm�S�����;{�N�:^%A�o�?�4����#3ZQ!G�`P(���* @�Z4s�ۻ�+�aW�:_~�W�q�r��C�����_Y�U;����ߖ�գ�y}K�L���k7�X���Q^��>��
pw$m��*]}꡾Z��aŅ���Η���_0g�.9�}��}��<78[��U �T� �y������LO��_��<��m7��ECݝ���/^���P��4��{|����]��`s�Rɠ %��R�bڨ�_���}~�8���]�KB]��t�����
<�,OZ��
 /��  �jWΝ�i��n�:BE���\��hL�~ߩC��gO�1zy�Τ�w�R��v��0�Q>0�1(SGV����)���Sf��0R�OюQ�ˋ�]��/w7�8�d����E^   �(;��9��7]p���=�8������PC��.���7�U���LD�;2Da(�1��QW�sgר��Н_�k�j�ڶ����[���xhF����i�� �](pdv$�\W��1�����rٕ�dx3$�KΨ�Y�u8���ħD'tw����Ń�ϝ6�Duk]�2�m�d%&ӊǞ�J<P9����c�f��r�E�O�1��������Z�x)��0�%<�=���6  #4��+���n6�{_A���M�
/Fg^& =]{Ҍ�lײ�K�~��n���KN��q{>p�4����Nؾy������xL8�m�p�TN�|���YcGh�;[�p���7S�}f��V����k����+N��D��D.��i�����n��5Ǆ�)�Ƌ
��X�?  �B~���;%%۶p<���ro�䔙��gVd�!PS�pm�v�j6,�?���c���Ꚕl���6s��>m�
�=?�T���C��=��rwНҵs�[�p�wl�*�B'  p�{�N��hDv�U�w�(0�Dh��f���k�jN���o��xݩ��4{�p��U�L�R\���;B�XDH��c���Q�S�}wڬ1�u����v��E����9�m�7��S�L��  H�y;�;p,XAWl�zw��3&{�׺S�x߻�4}��W�����3�+w��,��;kꘌ�-Eôa�9���E�mBz�3K{G��]R'wڰ��^��;9������=���c�v��z5�ء�]�Բk����)�ȊF�oc1KK,+k�-���cU^S��G��I"  �"�+�_8&,g����]p�S�h�W�ۭ�eE�TY6���������"}������;�Ϟ�͛�yѼm��)����R&
�jӌ�5e�"-Bj�5C�G�J��!pǐtos8����H9�;{�S��p��W
��-�����~'���R�����w**V��46j���[�F�׬V���Ao+TY��U������*TQ�|u�[��ͧ���ڗx�����3��@ߏm� �3�#�Q)B�p,X����V�~h��.'����˶��տT�
Cz�ӗ���|P��L|v��IS0M��]ϸ����+��T龰f��m+C+4�B%n����/*nRcϨ��5���|/wd��pT/o��ɶ��������S��w�2m�9խY-ۣ���:�u��˵���4l�4�<u�F/\�`���8�ծ�Vm;HX  R�AS�cιؽm�O��rzJ
�w5U�TH.2|kg����15���t���/T�nvk\}B���~]��j��{-�T�;�~�}Ʌ�Ή�i#*�Ξ:e�H�Pf���^RAk��%C;��}#�*]ܑ�'�ڠ�����-��Q���u��U[{T[�|R���W�'�	���;���.�;�\M��2VW+4Eb  H��v6�;�v���t%�m+.����ѕI-�fw�.��#:���yС{�F	�gM���z����q5G�����so��Ɇ�3F����h��35e���{!�h��y�/�����$<S���N��,��/k�r��}D�=�7E��_um%>�n}�	m{�)�^x��\}��F�T.k����| @F��U�웁���񚺟���a ��Y��rN�y]K��>�����<�G>}�&W�����;�q�#gM��>y�ۮ���b8'twں��E'����DجL�q�ٚ��e5��j(�������ަ[�&��[�9Z����n{��={��Sq��w.yQ{^{MS��F�.�4g+A��p  ��#ܣ�H7�8lL2����ɍ���8G�^���c�6�}7���J����бy���)�s�<q�����U�g�*{��3T��e�4�
�qNV�Kݞ�N�^[]#���X��d��0��e�Z��Kxr-pw�Ǭ��m{�ie�x$���S�^Z�9�p��jj�K�+���p  �@K ���EC��F0( ����*��>S�]w�n��)=��^�����Ǖ^xu��p��}v��w\��z&���k<:��צ�gɌG��|��P����{��s�"��V2��;�D_<�Μ2����6�j�{�������杊6p穓F����N���n}(�{Q�؜�J��͛��O�Km�3��f�֭Z����O|J��;O���%��/   ��,�P�n�
�� ���(S��C�E���O�����z�	�/�����/Ռ�W���n�Z}�//�y>z�a�cTY����3����9�o3�1 #J���Mש���Ť�r͛8J�=�$l��5���U�4��L7,�����/�yw�^ظ=��Ϲ�ȗ#�/w<��޾��n��l`��Zs�oԼs�f|�:�B$�ѿ  ����= ��#p/(��0{xq��	tT��xϳ����������t?R�޽���_xK_hi������:��=���"7Է(�C�c@�P�{�~�a�!}d�,w:�>�Lq+�;���}�7��6��ge��yDͻvk�g?'A��Ys���   ���  igw?�U0���U�+J5�:F����<�mr����������������2N�~��u� �v��45��P{�H5w��'N�����&��}ڈ
w�՟�6l�]+֦�鹗2e�ā������O<�l������_����[)�J�; 	�!pdN(��	p�X�w�
w�U]2��+N���kϕm��V�_q�#Z4c\�ǜ���O��$��%l�TY\@��� pG��+u��;�qK_��Yݱ�m�g��j�~�%�Pٻ��ֺ�x�i)�	dy�����������?��y��/
�(E,� @*u/!�s�n�Gk����84���V龳�Y���N��-�XJ�vGQ ��D�"pG�f�<�g뿞Y�?��v��o�ا����^�҇{���`����_�v1`fo�K���{�>�\��޻z�'?ּ����,|c�Ĩp  )d��8����fw;L�+N���t�[��}cӐ��U��(���;��0���p�v�s��t�7�;����5��9f���^yE�O����uz�~�?�)��[�   R���1����=drAE�7'�����:��;���̓چ�a��� 1(҃W�V:4Xꄊ2��Y���#+�����m�?����S,[�4mߦտ�uNd�y�U���C�|���&�x��N  @&8��ݶGf (��?�i�e����L�/�)���:!�)S�;��a�����G��@��}~�+V�o�2L%��R�j�-�J܏�J̰��hD�s?S,ܦhӶ�m�� H%A��:Cwg|�G��2�u��wy�;
�ĠH^iHZ��қ�_y��F�i�p���r�b�~g���.;C��݁Uw76k�zm�w ��1�w+ћ���{��6�s�*f�аiӕ-�q*� @
u�poݿϓM�E%*>m�
���1g[2cQe_,�?�;��m�!�m�ZV>�H�n�qO0q�
py=6���ۯ�P����[�5�u����_�s������R�B���uܝ�Q_��uzb��}�Ο>AE�����ҋfN�������<���m���{�v+���axկ�3~�ì��!p  ��U�=@����<[�����170��T8c���R�ݷۺ^V����xL $3c�}����?���H��vw����"��ܑ�҂��9;��N�����x�+bY�s�Pt��)����������+� �T*<�
�
�����v�Uv,���H�p�~ؽ�Nmm�:��C2�d�V�,��o�x�a ��|
�8ɝN�n��w'��Qv��P�n���1W���cl��ߑӶ��9�Z ^){�)���u�O�Ֆ��~���+�HI��(�"=x�!i�CD&���N�m������9?���ޚx���ny�a�;�<��LG�  R)0i� �YZ�N�|A���Lo[�t����1lw|��eZ0i�f�����{�.��;�����o�Tb�\���U���
N���pT�}�О��tp��#+��{����~^�.n3h*     DSTx�����7}����ilѕ�<�Gn�L5U�>��0א�H�_���N��!�w���{�U>۵t�&_�~���LF� Cdd�%g   �5�}(�����79z��iG}�.��!�C��p����`�#�ԇ3{���7�Tӎ��k��������?)��    �Hk��L��/8a�����?z��\U��s���B���s0�w��6Pjv���#
Uxߗ�+T�    �I������၇����7�O_�I��D�;҄����^���_^x�Z��#���\���ի��^�^Z�I�]�Le��    �?�0v�@��UC
�;m?��Y�ޔ��;ܑ�U�;>r�'�Z�i�2�Η_�me��4�������    ��ކ�!o��g{�a{�gj�đzi��>p�T����^�8��e�}��'V��yQ�t!pG����]�L8�i�v��}��q�D��*     5�4�i��~q���ۮ�Pkv���;o������B��������:�rp��az�#=ܑs�~�5M�]&okS��MBO�^=cw     �ɞ��A���W�k���c�a���Mt���L��-��}o��O�9�en~hP�����mҁ�9�0���׭]+;z�}�M�ж2��    ��m
��
�}'l�ja��H����3toK<��׼�k�����/P{�ڦVE�d�&��9%���2�K�R�n�Z���M�ܾ��a��fM    �'�޲�^�GV&���,Y��=�\�~����	��:�_��o\�����rN�H��`��t!pG�)/�y�c|x���w��⑰��mS�ģ���y; �a  @vY��`ҁ�����Wz��+�������n�8��?�X��q=�v������������_�M�k4n�"���w32p'o    䛍{&���/�ї|�߰���_��͞���2����=�l��<W���N5�1����ٕ��5���n�{@@��#�L��̠����:��a�o-{�(�    �͆�����~��;>v�.��;lw$���ilѵ�>�g��`�8��3��V��@���O������ղg�п�ݙ��5    �g��L.��څ��(�7]��;a���_�o�~$��7���oyĽ�����.Ra �hs�n*ܑ>��IQ�R�؈ک����O�r�t#n    䛷w�Wk4�T���s�4�X"�i�a�%��2��|��=ne���>�[4}��@���i)�t2ܑ�.F�+�������}$��&e"*ܑ�2k	    sD��ܾW�M���<m�B~�����l��T[�~W������/�ﶫ)�'_d�l�nE�q�B����2+(�"���e&BI    @�Y�5���qݼ�C���x�M}��e�|}�pƸ���7n�N��I�V�lY��?bm     2ǫ���g�91%�6�I�����]�	�������o pGz�#'|�2�a)g#~m 046��   �ҳ��-T�}4=�L�N��[����҉�i�7M/)���/_�w�+(�g�D&�;     5��z~�v-� �^J��w���:�4#pǀ}>]s�t�9e����il��ww�u[��ݫ���@w�q��������om쵌׹f�̬
wQ�п@i�2Qf��     H���ژ��=�hqG�B�����	H7wHa����aMQ�c��g��p,�6l�]+���՛�e>���I�U�XϹ�4T�˰�䂊
���i  �bȖ�D�%[�l>�  2��olз.9]#J�_D�E��֎}Z�s��t#pǀ|��9���N�N��Y�ܩ%u�߻�k�ZhiK�s�ZVƵ)�!�/S>�   	~;��xD+*⳨_qw���:t�bfb��t�Fǭ���S�p&�;  �8���}y���x���=����Yt��)lw�����kO���r�����Z��ǖ*Z�qe���*�O��
���L�� ��AS��BVDe���~�sB{�OL�W�uc�ϕV,*b�G"1j��|AE̠�� x�w/����9IeA϶i���Wa�ꝵz�͍�w$�	�O{��O����O-Wms����{��鶎9�sF�S|L�M�iy�[���6LS%�ǫa�f����㔉�� @�l�>�5nZ��A�mB�/��b�p�{ˊ�9I��h���
/�V��  ^q:|�����Ug��{]1g����E
��>�ڷ�٢��H���`5�˻.������Ow=����_^��ְn�nq�uZ�1}��ţ�n��W�3p�0e��I�	��b�6u�2�I�;  �Cے�^��2M�3��,�R`�l ��߿�Z9e�N�M;ؾ��<~�n������mخ'�np��#iS���oy�^����z}�ʳU]R�~���և�l�n���ڕG)Q9{��?��S�	�(���  �0��_P۫Ol%@f�н5
��3���`�����l��m���";���&Ŷ������_��r�  �Bܲ��??�'>{�
�G�^��N��8�ܑ��� �Q
�z�i'SlI�ܶG��Qm;Шt��(�W�9�m-c[�pH�����p  �E֭T������0fY���JE�2K�;n�����XF��}�4T���� ��ƃ��:�����1w���F����  ����3w=�?\�>�P���W?Y��(lw������A�1d�#i!ߡ���,�+��RK�}�('����g�}ޣqKonߧˏ��-���{�S]����04�ڙ�KKU6y��7m�>�e*�� ���(r�m�Uz�MnО�0۩�w&�e�4������{߷K־��^��� �W|k�~��
}����wk;a���@~ӛ��gϾ��W�#�X#pGҺ�z��j-���mK�(nۺr�T�2���U��'N��k��_{[����*o�9�k��M��+��P��*e�Q�-$p�&TY��)�T>�"  ��0����e��U�v'�<Y  ��w[��ϧ>��!m��sk�����Y����W��}Y@& pG���5��\�v�¤�^\��c͑���9 /\3͛A<RaԂz�Ow�H�Ɵw��f'SQ�    �!�-}㡗T�ܪ���Am��ic�酳=	۝���V�ۏ���2�;�V�˥� �t(�Gf�TUiĉ'i���{�7ֱ眣LƠ��Y�L   0?}v�6�?���\/)�@�Y��s��Ԫ/��=��=���I۟ؑ��}���q0=���2�e=~�"���CA�pe2M    �oNO�W6�ҏ����[���kٶnm����R�6�
�4��L"�8c8S���
w��'�t�D5n٢|6a�be:�v     ��T��p���7q�>w�I����)+^k�����7��Ͽ�{�iK��;r��O/	���Or����?���U�qǩj���tT���H   /,߲��k��뚓���5wl�B��e4��[�d�N=�~�xs��"2�;rJ�4�)Ӎ�7OæN����o�ARg\�1e�v     ����^���rw
�LMQ�)�e�2�"1SuI�*�B���Bj�D��,[�mj���M�Zר-�b�^��U붐�	�;�VUZ���Ebq�5��%�zl��jj�h���=�񙆊CA�$v�v�]R��=�-�\�f}�Z��oȶ,�1g�������P�#  �WѸ����w$�}'L�M���޿��7��_�z��)�4��T����=���5���Sf��W��C���/)}��,�n�T6i�Ɲ��=���E��L�>�!      ����2�jX��O�<Z��ׯ�|M��]ZX����3��Ȍ�^��իռ{�r�ah�?|Z�aÔ-lJ�     0 �HZ��qB����X�ĉ�U�냧���~���P:�b������4�3�Ѳ�~GV,�\6������S�M� C�n   @�!p� :j=�LA����>uT�ʋ�+�?x����
w���0����̾Q.�M��"��oU�*�\�i�����      y�;�ֽ��i�2qx�6��)��v�wV���s�����j�E�i�Vm{�i嚢��tʗ�,3P��� �-   ���I;<z<e��}L���p�<=��m���]����go@:��T��Q{���\��м������ӷ�;+{_N    �V���*��*�0e�����?�U�`'�w�g]_j��ے���åU��ɮV���@���^�{�Ա�{�[:������Pןy����J��}�E-KY�45��?�7~�S�{}��]��������l�    R �|Pf4���	@.!pǠ�1}���ʒ�^�}��S�lӎ�?�h��$;mWN�◴�W�ԮW^Q�*9R'�����F/    ����e�����#i�a�N��M�����c�z��J�h<�+�;>�����T<f�6�_���Y���/~I��re;z�    �fȖ/�}�����\�t pǐ�0qt��MQ�t�����04��kT4z����[��ڔƞ}�f�SY9@j_,w�(N&!mx�  �������I%�@Rܑ�lx+p:�D����.0��*�<Y��+ܸA�*XV�ٟ��F�?U     ��p���E�;�w$mݎ}���+z���
��c[m�ҡ)UeaP��x�h-�ֿk�%Z��;��W&��4���',-U���P    �?�W��#d 9�Hڪm��)�5Fb9��Cc�:K�'����ޫ�O?u��,;�ڧ~���s�rm7     ^����F#�!pǀ�V�]�����q�@q�f}��tɥ����ڞ�����|�T�\y�F�|�r�->L     ��fk�;��@2�1 �A�����/�S�j�Ĕ�
G���D5W\���=�mO=��=��� PR�Q���1g��V��N���#  �ňdg�;����c@>0��M���aڼ�2Qc��EE�t�%�Դ}�j�x]{W�Ё��r�u�ܹy�~2�����L�}j���U    ���֖2T��ɿCr�ܩ��Esj��gWz������W.�d[+�۩|T2n�;M��r��Lû�y�N5mۦ�;Բw��maţY�H�z��B�ʇ���ZţF�l�d��LQib[N��|v��1����fينb����UM��LӔ�4���ϐ��-��U� q{�ʍ�e�z    �/QV�܁d�#i!�O'N��_<g���{�0T
x�-�ϧ|(.V՜9�ԟx8,3p�a]��*�,-��� �K �'���  �ɈG���p�C����=�m��8a�H�(+�ކ�ؙ�����8�y���y    �Όgg+\��H
�;�6����i��Y'j���=�qv��}�"kj���ھ��{��6*������C���s	�|ľ  ����p��w$mxIQ��?s����m��<�T3M�ĝwx�!���    ��cZqe%���#pGҊ�C�n��	����+��މ�_    x#[[���H�;�����=�����- �
�U�`��  �Y[��g; �HHZ�׳�w���>��Y��Ñ^��������ieg?4d���B    �#K�k�b
 )�H��w��=n�:���)1d*��BW^$ �W!M8&  �-[{��|��A�����4�o+Ƚ�eg��2T]8����!�    88<r�;�ֽ"�%��-[,θ�C�q^O     eknaS�$��I3{�;��mٜ.�gl�' �`e��$  @Je�g$� 9�Hگ�]���vh��*���n����.�[��P���|4    8g�9� W�#i�[�����l�'�Mxd� �z  z�S\K�.w�������inI�     ��K��F��AUV�ڦVŬޗ@9�ls�Tk|E��hЪ����Ԧ_,�����`s�����~��:-dJC�v�y    ����a�'4��E�����&|��^��q���^��Vw�{h�&}����;��m�f��Ϟ<ǋkF�S��]u��� 0H�  �
w ��c@���T}�����X�g�>�(=p�U*
�d�9StӢ������9�|� /�k�     /Y&���ܑ���%�����N�Z���1��������N�;�$ݺt��44+�
��q�ڢ �   ���pr�;����*�oS���]�63���E�(*���}T^X�a%�nÂ���'_K��,���o4�c    �K�An�2w$mn������|j�\�7}|�ex����WKL����bwwd���     o�>r ��#ie���юv2S����/]�c�w��W�@�����+�ᕫtù��q#��<���4G� e   z���m�Hځ����Ѹ���ԯ?rQ������Kj�m�9#�ܯ[��m��/�i(n���
wx%�    �����6w$m��}���r��-K?���:e���<��V=�n����	%M.hL�0��p,=��	�ᕈE� CC�;  ��,q���G�^�Y߽�,�J}TY�>:V����1��_�~�Y~{�>\S�/�2۝��})�nw�i)oD��     o��F�M1�w$mہF���}��9}>~[�[�t}��uљUho9����iy�!�!�1�     o��� �.w��\�i�:c������7���Ǽ�Fׅ�&��W��o^z+-ϑ�2�
� 04�8	  p�����e���HTW�����?K�gOV�gj�������������=YQ+����A_��j�����/�Zʼ�v�44��{��qll�|���J�
��q#�k��j�}�}�
w    �ײ�����c�b���}u�;�Ϟ[��{�sj
G�N�,�p�������wɊ+�����9y��Ϝ�k/^�y3�*S�Z� ��b2���]}�t��VIol�+     �*���e�H��w�?&�7�M����|'��v�m+���9�������Su��4e��WT���J�e�*-+QIQ�[o��[�L�$�V(dGn[t���dLiA�mt�����e�o��2w    �'܁�F���s��
��Amk,�x]A�"1ى��xL�榎�QM����I�HX�p���� <��ikm�o��w��@�y�J{�0�w�z�e�u��í:@�}w�t�N��wO�$~fEU*,)9�2�=g�����u�et{N�߯ʑ�����2�>���?Pa��U
����g�zZc�K Zs  �"pr�;Ң���8��5Ž��{g� �*tRri��4��Ж�r�g}��h�-���o��sN�����ݣ���Ӹa�=�M�    ���;c6�	@."p�����'��yGiބQ�3f��+QA���e���O��7�@H���a]{˃��'.Ӥ���cˋ    �l��A�Ѱ �wل�2]z\�.�S��F��w�'O/'lG�[��Nt��Z���i���3�
w ��   ���q'pr�;eڈ
���i���?���˯ܶG���k�����w/�r'�ij|E)W�    <S;m��XĽo�����9��N�{'���(c��@��j: ��#iN��2ӭ�uZ�$�%Սw>�h��mb��w�� 0��D�-Ŷnh������������&��T"a�m͉��cj���(�����m���R-�VFQ�  ���b����CWs;m�/;~�Ψ������紹�ca`0ܑ4'h��KN�������e=��oK�q�A   Y�0eV�P�s�+���#/uU#�������|�R2

�݆��bQ���HV\v����$0�D]|��@P  �	c���g�q����mvƏ���w$����K�n{�!=��˚0z�~p���?�n���t�   �lg�U���O)��-�>}���>�s*л�w��`�*<�r��/'�  ן:�G��>�R�L����* C���5�E�}̲mىi�i]��Q��]O�� 2���˴�)ٶe���$��i��-۟\լ姺�)0m���f(�Ƌj[����c���[��s�/�� ` ����|̜H��;������%g����B]�輮yš�.�;U�y�  ���j�  C��k�_�м߿[vsC{e�w�/�í�rv<&E#Ð*<�2��|�&�W9R  Ɣ������	0p�H�ۻ�t粵���ɪ,*��؈�J}`�^���ʳ�q���q�   ��c�-9  YfTY����}rwڈ
���j
��1��ܑ�=��统��4t��1�tΔ�T��������߽O�~~�[     d�1�%G{��(D��;,n�Z�i�;}�/h�J]<k�[�~���N�OE���i�/���z     ���r�w�wٺ�u���gWhBe����i�h���#Ǽ	���Sg�_]#       �A6�;<�����ə
~-�<FgM�3���7�w�}�]�ml       �w�L[4�g�ou'�S�^�%       7�~"m�A6h      @�"pGR����2C�=�;���\��%��6�#jh�@K�����6m?���       r�;��T�l�q:al������{l�~��r      @�!pGҾ|�sz���Q�gh='hn�6}�W����      �\D���-۲[7���~{�b�L��e�bq�6�hsm�6�;�U;��u[��@�        ��c@������k/Pq(�5OC����g����	       ��;��76��t�G/���G��F��O^�xl�����nh       �w��}u����O���\v�����>q�.�=Y�x�uwp�H<.       ��4g0�-m�B��`@s�V����Jw       y���R
��W��V�w���z}������       ���6sT�n��M������Ϯ�O�Y�p�62       ��;��#t���Ұ�P׼�e������g������ض������5��m{       ���I;n�p=p��UV�1�o���is���]����zR       ��ܑ��ߧ�|��^a�@�       �\E����3\/nڮ׶�Ra�����~�u|}�0}W}�        W�#)+��q'       @��       � �;         p       ��        x��        �       �w        <@�       ��       � �;         p       ��        x��        �       �w        <@�       ��       � �;         p       ��        x��        �       �w        <@�    iP�o�B���}_,�����zF<&ò��&�-3�#\>Ru�N  @'w    H��*ݵA��?   ���    ��RG�H�"  �G� @J8���J�O�/�?r�ο3��5����w��?&Ӷ$�6���j�B���lw  �\��G�  ��)ڿ]��<{�el�_���=߶e��}��X��c���P���Sٌ�ۗsv��X�헜�]�ϖo�XÈ�@~1�  r�;  �IU��ʅ�5��PZ��<���a���ew ���_,����m�F�u X�����B����)  z"p  C�k��y��w}����Iʽ��|�%��g(p�=�  r�;  ���ԙS���w��i���״���'��~�qB�;T��
� �a� ����(uC��C��9'�K�7=�f��ʴIh�|DK  ��G�  mJuE��/�5IcGT=YF{�n���G'�   r�;  �Q�E����ڴ�^k$n��3h�ӫ��mTN��M��L{�v�	����s��   �!p  �v�ko�S_��)�@P�hX�,���@�$�@>��  @�#p  )�w����RH���K�9��9  8�;  H'p5�	N�v��� ��;  @��	� @����v�̮f���'��   9��  ��S���U�nЃ �O�l�A�N @O�   e��"���T����'�   r�;  H��{�[�F��)*�s�S  pw  �2����!j��,  @�#p  )������&l��   �� ���M�⁐|�6A�zɐ�y��n   ���  ���ǝ���$A�;��h)  ��� @J�C�RS��`tD�$�@~�-!��;  �#p  )�T� g �����R�-�^��;  H�X�P�@��5ZK�b6 ��MS?��\}�����آ�_}[�z�h��"�v�   �,HPG�N��3�x ���/��s�*+֗/���U냿�� �A�  R����݀<Š� ���W���9���3�� t"p  )��v�A�;����"N� �ĩn/��z�o
G �� @j����ũn%t�� ��&W��ړg��ؚ]� �8  )E���Pg}+�&��VR9�_k�2lKF��e��m���bXq�X�yf�kÊ���X�}܈Gۿ�w~�<U�0��~�_�~�.^x�B�CWq�޹O Љ�  ��i
�(n��,�U�k�i��c�N|��ў�ʭ���ŉ�lZ�%�C���UX3[��i�Q3V˷� t"p  )E5wo�L  �l^��òSX��	�vm׏�Z�k� �;w  �R�Q��	�mQ�
 ���y�:��p8� ��  ��e	�:O>P� @f3��WU��brR@?� @JQ�~H�O�� r��e�����#�* �!p  �e�w�Hfl  2Vd�r�6I���# p�w  �41��  2Kt�J�b��#1l˝l�33 z"p  �E�n�M���  #�ш��7J��S�n����� @J�ýS���A�;  �(�w���I1�� �p�   �8`mg�H r�q9Ǫ���� 	� �B�  R�
�F�O���� ��3n@V����d
�`�:@� @jq�ڡ{K!KL>L_]�@���|r���  wٱX�=ެqt���F�  R��@�ŉ��S
���p�&U��__:�F���A=�a�  9��Eo�8:*���  ��a�qR��]��?�+lw�MS߾����� �U���t�A2���  ����C�rG�Y�����7cde��~� �r�[$�AS��  ���'�u6?�,qҸ������5 �i�I#y�% �@�  ���٤�0��������aݼ�M��e  p���;  H-ʁ�u+l7��d��ߧ_�����_�u{��ݝ
Ǹl@O��9˶x��ѱ �w  �4h��M;�l���E_�� 䙮�(� ��!p  H�Ca;��  d8�c��H��@�  ��p�v۽C �� Y�?Z$��	��� @jq��? ���sg�1� ��   l�=��8 ��g�$p~@_�  ��= 3�޳�جx��k{ͷ���I�7�m[�)ۗK�@PMՓ �U���u��qd  ��lu�p�ƃ���*۵A�.ZXF� ���8�Hm� ��  ���v��s0����J��
  ��� �F�  �N^�yH��y;�Mڙ� �'#sNg�7��-�@a	��� ��‵��J&{{�S���pw���6 �-e���e��   ���`t�|��c3N�t�eX1پ�  @������ @�ضbj��J�����3��2]��2qwB9��j���;;�j�N ��  ��]�[�A���V��Q��W�  ���xH� �� �ԩۭX<.8���j����f]L^� :��.�]@rx� ��  ��}�V�hDhg[�;�fY͈��`����h)�{��b@8��7w  �"���F�V\��/#�Ou��t����PvrM �8�^  �;  H	;�&Y�7b��y��y{GwK���CӶ�s���% ������#)�XD �� @jĢ]w���aO���V^��}�8uB �]ox6�|H���@o�   %��L����G��
���6n��}���b�� Q��{�r�H�  }��  ��q�mJ��ƀ�[��X6�<h)Ӆ
w �e$�H�m�z��;  H	�[�_���s�j7p7�'1:�& �9o�� �v� ��}G{   +��u1v��hY�-;W�PV��;<�
w �]�=�-��Hm� �f� �����cq���勆叶)ٶ���j��������`��=�; ��  }!p  ��3]jmj�Vw�)�,�/P �x���0H,�b�ţ
��2����:�<bu��X�{{Ӷd�c*˲w&���w�m����wZ�3�L�8v��ٓ@�!
�M�`�--���Zh)t�=h���&찲�N��L�I'��mͻ���-k��%���I��I�N���=�{X�"�l춍lV+	6Y�f�Y�d5�f� sk3e����@�Cw �x���X^ �w   P	��[LNc�)�V�I�;�R��҈KM'J�".=K��$�c��h1���@Bk���]�QX��1���.�l$����)$�U v�b�204q�;('z>R�� ��:   p   �p��r)Ng Qo b�t��'Kדb&X����I�[(�����NS ❈����: %�  @5\٘��1-�`i� ��;@�:��ay �   �'�N�B^
 �P"�� (@�    �����]C��������{��u P��]e���e�(^#�{�q�^R{��gJ>�J��IӦ��u�|�s�T   �>��5��wX| b�v  ��]e� L�8�w�C�1�_nQ�_���Emk���)��%    ���  	 �;  DD�2^"F�qN����[kZ�^1�m�Z�NX-f�I��b2K��zn[�J+D�.���   ����C5 ���*"p ������DQ�P��՟���ѿ~|��y�C�M'   �D�� ��l�Y��� ������8�ӈq��P{�l2�    w���׽�.
�  �A�2Q�:D�j����)RA����l6��8텺<   H"2 ��A����=��5  (A�2VRƵc���4�ˋ͌�ܹs����<�j����F�J    �{�  qA;�� p��]e<��}I�Vw���\X6�    �� ��   �w�)���� ��PwR�H����     ��� ��W�C��; �"�*c��kH-�a�wÙ����j7��"�D��O��ECJߦ�hE����$R��M��y�&l�d���V#o6�#���6��1�m��$���gE�dxK^���N�qε�  �&���  pe㎈�<  �C�2�s��8l�N�P�io.& A����$�Ә	  C���Xz �]��:���
���| T#"pW_�����`�َ���4���� � �`�   ���,QJ� ��4M�V�� B��h���+�]���� ;�z!PXv �vס�� ��*�y^��[,jnn��5���A�;��|��6��㥿�5%%�0A�H突㸈�4��koo/�Z�y��ٶIC���m�j�mҥ�`0ؤ�4��٥^��3����CX��Ɇ���S���ٽs氍    j8>  B�2Q�q��DuuuOt:]CQQ�D E������������=�%�  Y(���2���G�T��"  %nT�q�&J�X,�< ��z���*��	t>�:�@  Y�!P"�<����5�� @�����p� B�t�" n�z��.��t礋�@��q\ @D�M  ��6 (@�>%i糞�8� 
�Zm2�����D��hR  "�O��;5Q  �v=*Z��p� (@�2���Die�ٚQ^@��Y�u��|��I @D�ع� aɉCX�-|�  (��*S�45^Ik�"���~�9���  DR��� Q_S  w����K�C�&�ɪ�� �I�L��[C��K��!�  ��C/�p�� l�SX�-���X���*�%�RR�j� x����ZmЉ�F�iE� A<O }�� V$��;  ��������b� xd0��Zmj���y��   bD�; ��'I�?"w�V ��������l:H�gz��S���v>Z���d2     �%1��!XXN �w�q\�4��X,� �t:�tt�����h� ��h�A�ٸ��   \!pW_��Z��~�<NE� =�9���m}���=N�������|)�E_J���P�	�}�&�33*�a��Xr�$Mo��)��ǘ�r��A�O����������z�Ҵl�X,��`��[6�R+�K��#���&  Dj�C f�  �.� ^`� 
��/a��X'�uuu_HW��u-+�#Z�z�t�:�d�)ǱЖ�,ev?T�=8Bky�;&������Z��Zo�Xڤ�Sl�4dHߕ,�;�/M��=xRO  1"��!����:    �՗P�`&��B����D�g��l6��N�*��  �,�3 ,5 1��a;��a   �*Ei�,�vʤ����N(�"�Պ�R ��u (���>�7bo�N >a� 
����yNL�0�q ��֐�^O��
 @4�b�K�(��   H�՗P��Y'�<:Pd�Z��  �() vX�4m��p0 �!pW�(���Y Y,�>`[d���  �P��;D��7 @��k 
��/���D��x��K	����| @K��;�2�
����]�p�6�S@w�%��$� @�~�l��`w��M�{ ?�0�2 �����sX׃o� %�U�6.�N;�V	�g,p���t�Χw�.�V/  �%e Xj����/���/X ��*�y�k+[% � �  1M���b
�c]~��  pW_��Jk <��<\�%�= ��Dۤ�u}!��)|��{[�CI�J� ��*K����ߋ� /BԱ�}��#[x  a�/BD������*�C@w p��]}	��) oX�����9ԓ �0��! ��� �k  P�pT}�vX���Y;��  � Ċ�2rw�^�f %G՗P<A�2����ɱ�E4e�T��Y�OA�s�F�hIT�	*����x��Z�������z�:�{n�G�R�M��j �/A�b��-�]a�#�V/_�m��y=��L8iS��Z(ڈ�kC��y�&�PZ�K�8�l�|�]���*���? (�^2�Z�Ͷ�q�����)�E�(��!_>��Z���f
�5��2O�S聧�޿����J�F�Wr��TiH�2���{灂�Q��)�d%A/ڋ
A?��U��38=Fp�E�^Z�wzy��^+ͫk>lǸ�h#KG;i����M �@��mDvp:2JWL6�L+YLF�;�ue�5� Qo�]B�؃x��J�m��#���;5�o8��ށ�F>�A�z@�O��~��L�W�z�� P��]e,DM�#��ߛg�X�"����Y�Q��vH��MZӥ�D�D[  �c<:Mrñք��}NG�m!y�:����ϐ�h%%-��ȐB  �@��5��:�u�Ld�h'sk�Z�l6�Ǥ\v	�$u�gj���N�o�b2��{;Z}?X���%w��?� �t��A�e�v� @	w��<ϡ*�Y� ����f������h4�㬕�4�i���m�%
]��h2�u��N�E��|�7��!�\:?�
�V$�Cdm�#��Eyb���W�~�T���3r(������z��鴃GP�����O�Ğ��|�,' � ��ʤ2��!-�EV���綴yD�՞�y>_�>�@m�o���Hx�	Z�G�����bCԁ�k��!��=A��t��gOʗb[�!�4���-#O��B����K���d��EBs��N�����n�8i�4��C�\�T����P��W��(�����]�y��F������M�R�0U���p�� ��p�#�8��g� D9���J:*i�K(Y  �4��w�!p�� B),�V�A��d��{腨�}�¡�{T�D��4^��A+��K:(�  	��
P9�);6���; �C�>�ktV�u�4�V�u:�tu"AH���T�RU�݀(¡�L����i'Y;lA�`����  �������C���k���ȡ��*AƙL&�����,�C֑r��pܥU�(���ECi+���M ��w��K��]4��D��4���J&+NZ�
݁;w���� � �; �$�x��H�f�N�+�F H����΃� ��&�q��4`$A�(*c�����Ki鸡���G���K���?�SM� ����.�p� ju �
��ʤi�Aܰ�lSA��j��4�Li�.��;lŖ�����(�NS#O�x�`��Z�C�>����80�~~���� �ŧeʗ��6] �B�2���x#-�)�e��j=���-�X�bW��!-)�sD`Q%e� ��]-w;�� ��o���#��3@4���?XCA��2 �������(��&�ɢ��Xk������q]�������p'B�E�EZ�Cx`����Rin��}FΒ��~�DZq(�>:��? (A� �б��6��u�ʚ��x��P���7x�p�&h�y�U���v��C��+�{���̱n��nF�v���ђn�p���lZ (A�>�B�c���L�s�a�ts�G�h�.�¡�;��'���{ĉ�9VJ����,�����5��L��4��s- �A?r
�����M�� �!p��E1�h4����5<��!P��ݱ�L/d�ظ�Tΐ̦��1�"�C���Cw|�`��E�ݰ����R��>����*��m� �AW>���:"sxbMN#  w�a���l6���t�5���@E}�u�SzG��;��Wۚ�s�:�<�-5g8A�a�q"!pWJ��BwA�NU�������C E8���t�����5	�; (�@�Y,���(��j�Τq��=ץ����GbaF[CᘶyMU}Fa�ɼ�Qf��A� ��4-�U�#��8�[ �;�_��h� �Z�3EQܢ��X�`I!��{�P�	���M�*��ړ��	C$y����p�C� �8�z��bH%  h� ��lS���:�n�t�eB�&�bJ��FC^i>Bb9�pW���ݎG� ���GP{���	D�46��}��'(����)���l~hY�H�5$:���sP��m�3��V�$g �����)$4��6I�ج���%�9�k��̞<�{M��}���HC�&,�=��  ��2��D   }��K}�;��g��.�8n�V��I(Q��!p�8�!p+��#5�U��I/�f!      %�Շ�S �k���8n�F��G0�=�p�-��^�E��w<���]E()c�A�      pW�N�Y,��<ϯ�8n&A@DQ4:ޖ�K�E�E��A�pB q�Մ�gE�     �����8���q&�i��`8 }7F���>q*%�+p'�a�
>Q ��j8��gǣ�;     x�� ��`6�3C�t=�; grN)�F��y$d���&���zD��'�      e�U&�,p!�b��b٪��J7��m�\����?vz���I�#��=��:�R�.�gŦI��<zizE	��i4��h��.�>�[�����n�w�%Z��cL���$�.�ԑ7V@a��=�D,����     �w��<ϡ��;��6ET�(��9%�ǹ,p|����ݖ�Վ�u���]��>���D2�P�]=�o;��     ��*Cw %�N!��������V�##�;����     ��  ��5@����{X��j䡤�zD��gg5�     ��  1D�4�G�z�p+���2����^�L    ���H�ӈ�\��C�iɔ�l��1�F3��6�mi�c��h}�jj���o�*�8.�?~ ��`�	N���uL��'�y���$b�q�Ճ�[&�2��     fxAM/-�C�i�*�����:M���Zw�}Yu��m�h��  ��v���mbADI�ppR�j��J)�d%q�@�̘U ��     ����t��
iFC�g5��d]6�T�}���ƎC���*�mn�HC�>4��X�k�sg%_�qE �*��H�o�����r�n����Î�YR3ɒ�IVC�\��6]�����k��l��c�,����J��6k��9�D����-FҘ:Ik�$��C�Ե7����4�}}��o ��A     ��q����i��r��T�*�G���G?^<���UE\�=���� �WP��(�����y��y2��'݀xgNΠ��Pr�Y�=��m���FK�9�d��#SF?2������F!�$�&ӕ��XL��h&CG�Z���(M�u�=̩Y�P:�:�$     ���z6�*+�s�4<�0i8}e�pZ����uTs����; @x�Ɋ�h_os�3p'�H�j\C���*�S�����G(�d%��s�=o0�g�G�Mg [f��
��q$���������}t�
    ����OO�;��!M�J~���׌+��#ӟW���NF���%v��b� %{�`��;&�Zs�t�bY�AW0�J��@eX�C��b[��C<�*��%     �9���^B���tZ����t��r���r��p@� [k�����!Jj�0��v��^M�c�u�g�D(3��p     ��Z��p�E��œ��+��9��w�B?�p=�s�n՟�; @l���O�ރ'*g;_<R�߿R;�Z�IKz�      ���u�ܭ���)�����9r��{k%Yl�jυ�]}H_ �Q����u߿�s�x�(��e����&� ���8>      �:��%ӫw]I�K
(V�2u$e����Lm&3��; @l�[�N2�p�;B      -X���=˨"?�b͂�z�kW�u�~�:U�L����� �8�j� ��cI�]�a�7      �]z��޸���{�RL��u%����d��]��/� �H�`3Y{��<�����{���; ı{L��ǖ�^��g���m�����p�4y%*�9��;����T�� <X�BsÎ�v���6�5��鲑����):�<E��^ڿ	n��m�7M��ާv�E՚ᡲ�����6x�F'�F�r�4~@źyC�_�����ʧ!�/��  b��tY;$���rQd��Ǵ����u��[ܦa-�Z��ԏ%V�,/[��/5�"���O];�  1�������BZ�>r�4 �F?�p�����W͢Ye�/��8�v֜����y"pW+!��# �Ï���1|81���A �3�`��ǈ��f\�|��}ʭw<t�|��u��_/�J�s��Ek�hf����?p ��������a� @��}�l|}c�8�7�^5�v�:GW�w  �8IDAT��	��"��  �Ǳ6$�!p�4N�������QO�����B���DC�S�������!3ɪ��r����8�LHh�1����@����Og�џ��O�H+���a!����dA'���R ��=\�05Z��'FM�x�� ��谪<����������Np��(A�*I�M���2����L\E 	�h��U��ێ:}�j÷�y0���
����[;<��ۥ�(͠�xU�/�~�h*��A�+:���� `�S��N��k]��� �����'��z[��o>M�#�vC27-��dx������ҳ��5A�9i���g���?��
2R#�2�PcO�y:��J-&3e''Ѡ�L�?��)V��@Jʴ�ʹ�l=�CY�2�8Z��/4��׌$奥�آ|���P0Ymt���~�[f��r���.p1��b��Z<c�d.UJ���y�m��A��; @�b}D�1A!�8^@w�.���#p�IO����,d0w�Q�B�h��A����4��/@$��(]��r��������Pnr�dePiN�ɦ%#�ihn��ϳ��4�a�V���qj5�|*���׌JϛF2�^����������MI��߽���>���9�c�H��e���eZu���|X��5��בA��߾{�x�����oU��^���2l����D���wtA�WZBˤ�"�A2,]��X�n���~Gz_o{�}�:����RE�liȥ�����޽SYE_{�#��z����n��Y�P�yg�����v��B׍N/�x���;��NE���t���]���y�H����?��hً�٥l��C�?�^F�p^z�Z���ܳ_�]%�t�`�`�SZ֯U��rf�H�7��/WSMs3�n
�2�i�i���)4e`!��{���}�n����\�����۟T������t����o�,/�J�t�s�n�:;P�>�����o�� 6�u��.�N��}_~�h*}���͇@U� ��/	 j�;��{X�(gyZ�@��P���9U��"9�^I��B����jI�f&�o�C��W���&��?_��-@tĂ����1��s���mm�l�I�o��'ϣ�gLt����'I�s��5����[2Z�3��e ?N�l�4:ݾ�r;� �=-�v՞�߫{�J_�:�]8�rR�}�#�;m���ەU��,�fÚc'�����=k��Ǜ�e�����O���_�B�>�=p}�?����G�"6i��u9|i�~���=�i|/;�s���VW�����=���?���%4:-�p�ay��b�p����왽��鞷?��է�N���4�����;�B�|{�ߤt��_�Gi��i9�ъ5���K�c���� 6�1}4�rfc�Y6~(=��6�_��<� ��p�bZWGZ�C4<�=���fH&������Y#�l��b������44ӊ;�ɭ�\��l�o�'U���/k1����L�~4��}����w���sJ�h��Y4�d�C��T�P`*��q'������w+���t�p�	"����vy�o���eꅝ{|�޼����=cMP�v������~g_����A�5�khay`gI�������^���5�\�n/�狴��);��/��^|�Z�}+��Z��-̣P�o�`i�p@�m�3_w�4�\�v�M�M���c�5���ނI�H�٧�Ι@���y��@� ���<���N!���к:��@�y8���;�K� ��N�)Yd�(Z����ƀ{��� "�S���O��U�j�W�6�/�p���+7�)lw���V��AE4oH�}+������tJ��j%�KG�J��;����%����{�
k�}��ʻo�:�k��X�t��-��6����^��o?u���=Oc
��z���J��7��g��Mv�h�ѓ^�yw�������o~H�s:XWO���1�r�2���76ӵ/�P��i�8m���������x%m��-n��6�������E���R~�nKǕ�Cﮡ� �A�2�j, ��?%eDV�
M������e} �8nNTHO]7�m�C���Dk��������5F]��uU5��7W@��o�D�vT�Qy�ު�R,c���v��fN�̤ރbG�豕���QRLW/'�FC�T���ܦa��ϿXG��|�>nP�rmwG����?����z*�۲T���t��D��{�V+����_��N��ށ!k�;����J�Ւ�䯻�N�|��+Ϟ�=�ut�B�ǰsձ�����VR�q~���g�V�~����Z��K;�ғ�-���<ZM<J�/soS83���Ň�|\�ȸzg�a��UG���|�\f�;H�xX9]>��rS��LK��}�<}�����õ�h��'����=��Ҕ�B2H�3�o�>-w��cƠb
�?]���/�ȝ�����3ͭ��f�N[{�3v���[Է���kj��׎v^7((��Ō;���D��,�zl��� �; @�Eߛ)((^<ZWG���k!z��ϒo&/�Gl�������H�����NsE�ɂ��4���lx��|����-r���y���I�v�P��l�A����k�~���胳��C+Vѓk6�M��l�4��˩���ۤ�+6l ��F�|���{���?�2��qEy���;(�&,�;'���n2��{�'+V*��ys�!�{l�u���a��G�������K�{l��ϳ=�ᗴ��ԩ.�b��c>,L��ts+m?}�&+��QێS���!��tvi	-���q�ΘL7��-��GG��{}�~����CGh��5�~y�et���;s��m=y���9+���r��a��'���y��i;��;w��y��*�jD�S�-��譅;v`�����:8�N|cղqC� $���g�`s%\X�v�p�<�p�h#��	PR�:za���!6y�N:v�Ȃ�������~U�]���l�/�P�$��+����_2�V>.w��ڈ>>t��1�+�f5��_W�����c��)�N�^{�9�~����t#�[�,��Os.)�ԯ�9ȳi<���%%������S���cIW���>���cm~n���Q��}��>��J��U���������m����c��}ܮbgc}RuܯiYY�H��T?�t��8v������5pg��<�6��*����'(����~���Չ�ъ�}w�޲����h���SF�lFY��MH3���j T����G�h��wl$㹷H7j
�'�",�X��F�gf�A�p����3������q���TI���jH�-�!��<thP��9��b���\�b(:��?M��2���xp�T������p�to����q�E����һ��ſ���=pw��0'9٭�W�I�j�{
��1��Qo�Q�D�������%�x�zp�4�ͪ���	��ޮ<T���쳵t���A^�u*���V��#'�:
e�-�v�R��C׼�&���������%�)ܔZ�33P?R����54f-����;��߽R��]��y?����C�(ݡ��b=�4n8�tu,��#*�	�L�,Y���%�����+���Z �r��Ow��a�����f6�h2�y�Z���v���g7����6��Y)I�#�)iH����K�4����M�a��uK�Ք��C��iK*U߻+�]��3���s��W+��wזڻk{K=��J�����@�������V�/�'�K\ ��ng�Z���[<�|��iT_���u~�o���g�,��[��(#�޼�z��ye�iʟ�C�g{ϒx������R�s=韚B����X��~z�L�v_�$p�7������_��j�������_�@��7Ұ�9.���۪���E%��������*�7�;:�dS3��*���I�)Ӥ���w��,Xo����7�\�Q.�����=&��&̧D7cHw �x�������Oo���Ç�Eg(�h���z�w�8O�Y`]��.�bE�1���*��D�w< ���CKvO�r����O{(�4��sP�-=�$+�N\hq_�p;E��~)΁(��/��P�KX]��I+��+�!����)R��ʿ�z��C�SF��4^6$G��5߼���Tߞ�z}�����h���#c���Տ^_����������1#�����͟I�����~�����4�CKm%ϟA���s�q�Y���~�8*HOS|���
��������|�������~9N��Y_	?�;���Dc�bkk�Ipvr����OKqܙ��N{�ǥDT�y��ŋ��^D��x�Ӹ�m�Iߚ:^>�����ݤ�|��B$����yp���z z�t}�_w�uFѡ�5���  t�V���X�i�ɱ����ri��Z���P���?�s�ǰ�Q]w�⛵*�i��Z����wQ��K�ʁ��������{ǲ J�<�L��1pc�;+����khk���;�\>����b���?-�]�ɰ��ќR� �=F)p�T[٘���=�i�C=r�)�/>_O�Xz�bP�����St��� raz�d;��N�������_��T_��N�䧱Vun㛍�߃�m��d(����R.��w�y�ze�~�y�������ǫ��ۖIˑ�s�ؕ�v����+�����̱5* @�W(� �<��V@����u}TJ��陊Ӥ���3i��<�5���i��3����� �)�� ������=O�ٺ�ZL&�s�PU�^~"����jz�>�V��x����guc�AY��to�Ǿl���	��~x��_�k������|�==��,���ӯ�\O�khÉj�R.k��
9����1��ݟ���;�gi59����g\�:b�߯�-K�.�M�>���o�E�Ϙ�x`�ӮŻ�o�e���b~��Z:�ҦxF�s�v?��� Z����q�
�5��p`��C?+Iʏe�+�sX'N��������d�d���[�~)-GW<�������P.)�e~��ܻ��dȥYL}��]}��%  ��qk�疈���uP����yW�J������%S�����_���@-l'Zc��Y��d��"Ǔ?��gӑ�(��?w�y���+u.�cda��c�pD�����`��@�S��v����]T�}?�`XwG��u�����ZH	k��ّj�y0��	�=yu��-���;�❯*��;H���#����췏5��6ol�]g�h|�u�Y�{IE)-($Ϳ�>�x���;�u���+�w���lk;t�/g-�������#V{����r�:,4�Mu�_�N9^����l�'V��?kGwLK�\%�E�NS/6���ЗG�τ�·_P����G���dt)�LE�mA@�R �Sf�k�N"VAa��=:X��^�n�ҕ��o�KO�o��6����jP۩��M����}��l]��Dy�
އ��Ѷj�Nx�4��k�߮�L�`Zi�3g�����v[��Mo�R���������B�1kaY	}�d�q9IʥcNy��n����~V��1���x� r�SN�X��Xk��G��t��2JkɻxX�ܪ#+�s�߮�w��14��wX�۷o�=�6������a�|�P����R|�����{��94�ȋN���X�G��N����N��^�_7l�_^:W����K�������SgƁ�T��W��N-����詯�j����ۦp�G,���M��KN��s�t�or�6ο�q!75��KNJ���*C�e 1{�˪����{��m�<�>�Rny��S�|�.k��T��/�v*d�Z~|��z\9=�Ӓ�;p��-�����i�/(��a-�{��l�q�U��![8�=c��y��V�O\3�>�w\�Sȁ��=ʵ��ݭFҿ�\�*�ka����ն�ѩf�V�Ƶ#��_wnAz�����}�۬#�����})�hQ*��J���ե�`jA���Ov����W�<���k�����è���V=��XV���f;�����ܙ>���YN��w^?wX,���J���<�j})�N֒~C�)�i֝8屬L��A9��eю549��દ�Yq|��k��\~��#'�mL�Y�)���%�.XH�FU�[��ݕ��g����I"	���/vז u����8}F�ͮ�D����cN�"N��shh�-_K�]:׾Su�|��� �Z���
�6�o^W�=�NG&�s����);�@w�K��l��<���lY}��)t�sR$��W�"�$��Eθ��S�_Է��S|�u*�ˢLuZ����>y@>-*DW�(s�{��f+�_u�s'ì����Ν��������;�^~{�����h�=g��"�O�L�a�	­F���_ٵ��c�9�rR�nn����(���dxc����a%eXi�R?�A8�M��ҹ�ၣ-��;�8�5t�X}��c��+=�����u���M��I��[\��O��5Ј|�М�w�޽|OfR�S����뮳�@��U�<����6{��@-jt���W�f���>�qh������{t�+�{�C� v!8�ű���-P�'Ol̄�M�S�"͜�M�xv�^���OO�)�
��+6��) ��H��VJ���(5IO��.�u��Y<z�b��Խ�3�l�t�"x�������]���殁��Q��˼4��̼�����/!��0����/�F��ȭU�dg�U�dLAy:לr���>�k�u�=��&�L�v����]�̕z�r���'���T��n��2�P���R�j�D���n@f�\nbl~zh�j�i��q�7m�[9%�^��۫g%a�m����*�ά)�_���Ȗ�Ǐ�Wv�#o\�R����VVF)p�i�r�2���-pgީ<H#�g�����a�Th�?mp�S��Q��XZ��W?�d���6�V��;����m�aҺ����v��6��{�c�'iC��E�f+�w�!p�Pr\���J9y{x�)$j�����c�aN�c��GNѥ}Sk[� �rl�%�ЙbZ�{М���(�u������MO�S�4mM�rG��0Jz�=�3�ûE�˗���[�����vg2�<ׅP�� �х3��1͓�n�׏*���&�˦���+/v�˕h�Y�Q��~��R�q��;��Q���I�yrؿ`H	�����4���O���R8��1�dmW��ùQ]{;=�n��4�/4�?6�fN�x������(X���]n�b�,zc���S��qy�ە���5�k�2K�.���*��]ZBo�v?K๭����Ӥ��ޘ��n��u�󹢻�~ �0~$�a�{�+�����~B[��4+��a�!@zDZ��"��\�i�^>[d���,}~ܻx����ꋇ�% D�>��n%�X�`-�-�	"Ü�_wGg���:����p��y�
���.Q�N���Hu�O�e�YE�������,�O�Ȃ�@^�c���{�� D�`K�|e���[�6����˭ܿ:n���ڞ���^�`�������t��!p�X��9��!=�������^��;�?f���'��k�$���Ӂs�I�{�Z���4�c�=�u��B�Q.?�j���t��1��y�n��������(�����fӝ���ӛw�����������T���C�h�~�4lY\��}k�x��Z�o�9C_y�=�^��\�T~��={�O��n<��D��r=�3}i5<m�����XE�Ϻo۳�cl>��:���v�♓Oo�I'�Z��,���x*'#��{=���,d�^{�Y�!W��^zG�ζG�]���������Yg�_�2���q��i��=���̔�m6��w�9�[ ��>�o��SRF�XϪؘ	���ɔ�x�퍤�h!��-�è/-�Ԥ�ޓ�8�wU��PjeDq~��)I.z6�Y��9�ΡzAF��w���޲=;� ���I���wfM���Ե�;�g����1y��}�:��}��3h�B�yfbQ�|��l��y{��ǵ��~��M�&����������,��F����������r��D�ʗ(�.��E�=�{����6lw�_6����S&������3��;L�zL44��Z�@��C��<N��,lv�VV�5p�xe�56˃?]4��n���=3'�_ֺ�q���k����̽��:"f�Tn�<��ݲ[�q�<J��ZT1�*�+7	U=�7���'N�?�V+��p����	$pg~<o:=����r��=�UKۤ��wGv�������ق�S��Ê B��y�^鹉�2QƘ�'�x�E�y�F�`���K��s�����>[��ک��1�[}i��S�y�Hڮ�f�͇�2/����|?�N��J��]nw�������pN��5���$h���M��v-�:]o��O!��4d���k�ͰNS{x:�<\�-][�����~�T�8ԡ�jB�	^_�`���:Z�D =��2��MW���^�ZFA	�]���K�,7K�~�:�=t�wit~י%%YT.=���
ӕ�`ۅ�(��<���<d-��x6}���ݦ����tߴ	T���w{{�X��B�� �e��<>�C�w��ھ�@P�*��������k��/o�=�8���_���rq� v��t����:�Յ��B���c��Ѧ�S���r���-D?��]O~%�{��j:ڠ���||��4(?>T�55!�p6��[�6���r��Q�~�����f�VZD���l�s���W�U� �\Z�����NS#M��-^�m� b���R�h%�C����z����=;U��y��H��ޝwג2E-�X�v�rͱŰc�w]�w�.��R���>\#k���v�:���kސ��ίЍ������D��K鶉�=N3(3Cq<�[��V�J�{�������[M�en<�pw/r�	��m��N7� ������]F�J)�f5�WTu?c� ꗪ�2�������V:&��):�gy�Kxh�4����n��z��ߪt�Y$���	[fY�¥��L��}G�-�!����T��>���t������_7NMO_���\��U��J_}�]��O_�KM�P�CP�>�[ͽ��޲���F����=�9�����\"pWw ���l�u��-P�9c��{ �լI�$k�S����I;�";SI�r�huNaBqV�S9�ܴd�ec�6cdw�Ù9Eݯ���`;!��-�kf�{Z��w�B���/��|+=u�|�e�Hy`������'h����Թ��;B�q������'Wo�o�C���ӱБ�l���Yr�oe)�=�dz,���_[��MW������A@��Xl]��+��g^s��;*遙Sht~?J�VS���Z�{��>��b��٩#�~�8]=������s.��~���45M-���Y��s��t���/:�����YII�o���NӅ��TO�9�O��_������l��է�c��l�������~=';K`�n�w*��n��'�(�ug������!�h�t��T_i�ȶpgX��ߟ=�~�n���p|P	"��=��ɘ�'�R ��[� J�u��ʳ�116e  ��&��3�J�,YF��zH�^��D�m�A܏/�!JX˿���5ǜ|�Ёt��o��[�f��j{~|��:�����k�K�0�o��Ye�t턮 ����������V8AU��U'#��C�\:t0���)˥#�T}��`!����c���Ɠ�i�:�m�ꤛ�c
��-|Y,YN�?��m�c�vfɈ2:����묣���מZ8�~����7��ҵ��R}�e�+����n����,k	���o+���X�H��/UA����r+��;G��*���l��)��q#��a1[=������߬>�`�ʠ��tz��ͯR&�OM�K���	X�O�����R�#�ˇ��}�X�{���p���6�8E'/4�}��fPv&�,�X���'-3\ؙ�L���{���L�i4�_�S��Pz��k�R����\%-Cm?�̶��Į��F�R<�����i�Ѓu�{���t^�{�Qa�ɺ�����X{Կ�\!pWw %�����,�!�� @��4jt�4<I�e��,y���0�'y�\;Q�����7_����]�Lr���S�֩#��d��U�{��-�["|�������t��Z��)(�·�����nH�:���I_�>�o�?�7�6�YI��o�![�y;@����q=���Z�ܔd�>�w���P(�ʤ���|Xɟ��P8���ۈ�CS)�u(��� ѯ��D������۫�m/n8����*c5�E��
 ��{��	J�  Dݓ�S(:�<Dr�2Tϭ���;k�7�m������M�kƖSa�{+�T���H�����[{�4}XyT���;@��=	 ��V:�Ё���g��C�2ADԦ�P��'���x���gb��}  �u���^�T�y���,m�J�4�wR�Z���8��^��~��:�00��*�I%4q`>���ڑ}�����ͣm�g�gޗ��  � Ăwv��g��D���~,w�!���q)#�GA�  ��z�V��sCs� Z����O���ny\NJM\@3�����4���}zV�v��B�<w   �7���Rms����ո|�����]e�� ��c�D�j���  ��4vi�����t��SFГ��Q�6.�Έ�^ �hU��s �Xc�W���-�L���=G�:������+3�	�'zQ����O��Z��Tç�   ��/-�f)�YeŴ`� �3    ��kwѽs�S�.q"d�l�_nf\�[��� BƱ�;��i�];�~�/�o�s	   ܰ�}Ɛ"�U6�fKð���3���"YW   @M��:�V�wNM�����hmC0����; ��(�������s$Z8n�J� k�&}
 Āۧ��y��m&Y���wג���C� 3�Jr2���H���~��,�5t ��O��M�$��i�z���8/�L%A�>��Fb�n��y�!t��Q4���4����Z����G��=Gh��3d��   �?|��n�4�R�:�wl��[��w���p �/��n1��x�5�|eJ���} @tSܟ�[�|Z�f��[�)�ͤǖͣ��J��:�Z{����z�������A�����]s�Ӱ�\���>�hp�̱4q`�����g�8_�9��?����ٖv�����)��*�GO]7��*�:�0L�w��'j嚦    ��TS+���m��˦S�{f��{�|��AI�	��2r. ���K��f������� ք�E�ٖ�r2��{�ɭ�%�utɨ!�p�B+=�n7��y��z��c���c�'L��FZ���"�u�ۥs�=G�g���y�"�~�0�����.���>�w���⑥��m�Q�V����Mm���#�|��Z}!;   $����I7NNC�gS�b�s_�9�BI��� �(��Ԟۂ $�|�� b�ʪ2Z���d�f$���Y�t��}��.�z�J�y�Ɋ��ֵFG�~�̱na����t��U��ESI��ȭ�{�m6���_UZ'rR���K���u�nD~r�4������p�|Z%}���Ѩ�"?���u�[���u~��<�:u���x���C�y9�/��R:2w��j7���-��Y;�k	  b���+����_Kz��궱���VRs�)$�B�>l�@Hp�����Z�����v� "p�����jy�E����Yc�E�]T��@O~�����#K��6-I�t��?{{5�<y�"mɸr���W�T��wLv���yj�v\f��o���w�C[��"�WWͲס_�4}q��>��N44 �6f@�>k<�1�t~/ێ����YN  �v���#��7��'O��-���C� ��t��)�w��� .�+@��j�*�u��i�?��I_�Gn�i��*�e��_ic��m��d��E��xT)���E�����r��hpŨ!��Z��=I���];�iܱ�f�������I_�9�~�t�<��1e�ٙ�j�װ���:��^��G߹t�|��_�  6�Kږ�2����J�bg�9���C:O��C� v�������q�wT��83����|�����4��}v�>z�mt��HѢ8;�iU�ږ�ߥ#&����O�YE/o��h1 ;�~��w��ES�47�~��M���39lg��>�Ǘ̖�I%rK���"�u���C�S�H��<�Oa;�j@� �f�=�~&7*Y8��b����?y�*cᚈ� � �%����cf�; ĉ�����K�Ғ1enk�UGN��ﭧg)��e�د7�w���z�i\7��w^YA�	�i������Z�=F��}s'8M���}��Do�fv�A��j��_��F-Q�y�oiI���l��ڥ�7����i�n[���;�j2I��t�=:��  ���;^�����R�00�bU}[']�w��=���i; ��Ea��=8�; �6�y�.�J���֢���=�����I�Vy齁�ڪ��쎍3:����i���65Z�8���מ���~�S'�����lrz,�p5ݡ�� �)-� _�����/: H@m&3-}�]z��+hfY1�v���y���oRe��U&H�w�G�S�W��fc-�y�V��]�ƥ�>F��,��9��cmA<��Z����b2�Zx�_-vay��Pt�}\wG�l���^z?XR��ƧHӺ��'��x[�H;@X@�b��kw^�V����y�m�ܦ}r)�h���m	��J��@OV�:���i�C��h��L=M+-���u�p�g�x�\R�4��?�J��:��MR�t�1���d%�5Z�N�?-���e˭��[ Q��۞9��4D�N��@  �x��m�k����q�"Z:.vj��m>�������~!pWY0��� [-K�(����\��V�)��M�~�F�Yk4Ӥ˩!|N�?�� bSY�Lz�Wр�޺�,\g!�QV�ݛ$�Z�SJ��z��>g��X�vV�a|w`��j��Pms�om�ڦ6:��!]�J�;hO�9�������=c�\҇�p�]>�~v��i؎�L��������>^�Lр�o~}	�(ȡ'>�B�X�����A���Tz�Y򎤦�/�7wVѷ_��:-VHdSJ�� $0V
��/��Cu�����ڷ��՞����g?���Մ�]}�<����� �&�(�^���p���ȼp�b����v�N�\0�,,�Z�0�f5u���MFi�.���MƐw�����SG���� G�����>R*�������壆ȟы�_�TJ�����+�*��s��__Uu2����'�̡I%]�>z�L�a�0��+ik�Yy�-�g��ճ���0�M����d������o��Ƀ�����sg  ?֘��O�������7_*7V�F�m?(o煣�w�!pP&�FV�5a���3^B��`�h4�'���@�yh�Y�:O/-����p�]��Gr'~����P�D�*�;o|IC�g˥U2���,l�ڋ+hg�9�ǰ`��_�}��Wl�h0up!}u��q�
��'�_G�o�'ܹ��~G�+ҷf��?��A ��*}��A7fRi�|�� ����i��^��_9�n�2����6;c��ﬢ���s"p��0��k�����լ�' ��B�;���`��+�o>@����,�aЅns;��o��}�~�l.-W!��+�Nү>�D�N�S|Li�Ly��u�z��>�5u�9k��xV���飝Ʊ�����Ϡ������/�3�m�{�x����]d�^��z��Ľ���#�U����D�0[i��:zm�> �����ae�^����Y:�����|����^Q�UT @t0�6�n��c'���k�;����81v��%�q���6Ŧ0�w�#��N]���}s�����wo�N��gЕ�����3�y�^�j��w������ơބw�A�V���	��ټ�n����ױ�]}q� �-tO��eO�A1�# <��!A�%<�Â 6,������̵r�p�|(�\.���@>�j�c���
��Z�6���D�OVï�lb�|ZZ�(,������>�i
���p���x 3��zv���'\]c"?w�:X�<{|�J	|p���1���i	���At�n��{v�k��v��AD� ��y}L�̈́_�����8'@C�W��d��Հw�!�� $X�֍�UlG�D�N'�K��M�8Y��S�TO.���1h-��AN�Uu8SR��Zbg�%���kU5�:>�y�DzL��%���Ǵ��YX;�vȈ�t���E�),�v����H܉N����~v�жV�?AD�폿=R�ҍ�Ra��^pk�l�Grr���>�����?Մw�A1��� �����j���y�������}1b"���|,ݍ�.s�l�~�v���76�u�lh���y���9A�;�R��Y�`�� 8��6P\Q_l?�����"� :'�N]`�WK`J^6���FwO����v'�V�M̽���ǂK,�� �]a�$D��f�m�X,ás�8�9�W����Rә�7A>JNb�0X���& ��A�k�R�װ�<��������G�����nI���򼰼
�3q��_A����n�!"DHA�UB۹VY��Ե0$_�-��u�V���^�A^r��� 7)r�Ĳq��Q!������"�0F��kePP,$����݉ZqW�	���M� ��f��X,���ī��h�A�Grt8�8e$L}}��O� }ϣ5τ��#L.�I�^��W{Aq�ӭ��KWA��]�O3F�o��|Y(���񔍗Vn��{g��}'��X�u<��oP�ټ7{l<u6�8�,��� �D*�#���ֱD�ƧH�����f[ =g*���=��>�2�a�0F�ê�@�ǌ~9 i4��y��"h�.���7H�R��DǱ��,K�a ��RPf�,�	��AbB��G�X��M��5��_��+�r�L$�Z��_��M�������NhJ؞9�'�:���j+��k[��!�?��?{\m���U.�U�����=��@wE�~�Ε4�Ε�X��
�Z�..���*xJh+����x��=v�=��!�����AF�EI#1�o��8uŔ�߂�S�d�-�3atNJ�EA��)��{O��N������S�Ze-�U��;�wÖS��WI��Ov���E���� ����b�N]�Y���/O��-`�q��K7i�M	 �Mڢ��+)��m	2�˼'Ϋ>.�L��<�i��ex�?a6�S���@��4���9H+A�7@���o��x�V����g��&k��#�ߛ=&}~�Z��On�}p� �86,�Ep�����q���_�"�ć��C{��lUm�OmǙ�l�AS����Nz|�T��O5�ٯ6���H��� #��ٕ��N�N^)��G���#��55��B��B5�^U�\����,ߕ�[|$||�D�M�i�X\`��ە�g�\��?����CGrS� ��qC$�E��V�#��r���je�?�u��oڒ�&^�\it�� ����a,�ǊJ�b��h�.?���8^�!�����/�n�m��.^�����(��F������fv]��Ie�WR��ࢩ��18���P�t��'�}��s�Y���i!��w��8��������b�&Y���!�m6��`<P��4�-�A�Pc�	�	�1CӁ ��@�	2`��>���;���5�;�8iX�>{]Flx�N����p�r1�I^Z"��:D�ذȿR�|/�`��٩�����u§��1�E��6��k��e�{(&|�� �Z����b�����\

=�5 J�k�����P>�?q��]�="��|�f�w����������
ɑm�m�-���|:L��r����HϤ8�������^�	�����L�������,��`@n/ (����]�x)�!A���;] ��w�-�}��E�t(Ŀt��u���k���-x`j����}�Zr/�A�7e�E����.cA��f�06Dn��qp�%����Ӹ�bw��q�0����NaHp'Bvl6�Q�łw��M-:<�����"3�t�� �����>$ק�`��M�E����� ��	.�W2q ���jFlt��fq�-��?<nx�sU�g�ڥ��\��-��EN�!E������
��p%��R��:J�_l�_�~2�7<;v0sK�ZM�#�'L�zfݱs��p>�9r��� ���0":�6]����KlA����=F��P"b{��&�k�M�O���Hl�2�s���-��"Cһ�� �c�p�|JU�Ǽ0i�Gk{G���?���SF}	j�?5�C���[*�-��?]���N�0VD2B�0.��B�z���C�[��˭�7��!�x�ㆰ�r��0v��@��a���Z,�n��p ��f�U�'��F���&L����E��R�E&�ʀ.A�k��?��ݢEQ�^Ϭ��� 1""���[����b6�E���fq߲쎿98�E������<�2�`J^6�}S���w.�����b�������P>|�퐦���M�ė8O��e��]�z����x��"8\X
��p��
��V�M�
��3`B��]tI3�wW��]-��!����pg[�d�9���5�;��c2c#a�����+�8"Z-�Օ�P��Z)���%�����S�sGq�g�8���"�,�g�������u�w����OP��*#����i$�-��w��}@w�r����5aL���2��N�lX���B*< �)d�8��3	� ���Y���Pӎ	AAq���RP��+r�T٪I��ǋJX��aA����M�B�=xO�(���@ϭ�/���}����2�Y�����7uOci��PQk����&�w'/)�E�<[Z	3>�5��&���0xw�H�1�a��Y)�
����v���^���b��s��ά����kK��Dw0���j�����.ʂ�����v�M�0���:3<��Z��H��u�X�{8RSp�Ӆ��&����Y~�Bt�3mhlر����gB��-��/������Y79_�:������k��	�
�>܁ ���l�j��G�]x�p'���Z�!�����I���	�C\Z.n��^b��iK?'5q'KW��B������=�]���;����d��"�ms��R";�&N��l�jy+�aW���S��YJ�
���0е�bנ�!��Ć�<�ǖ#͊�"gJ*�������������7���i�ܳ�]}��>r~��*�F��$�@���c>���7���W�E�ԕ��	�����Sl��oo���g�� �;�[tW$�g���fq���`��	t�6��2�qh=����8��(J_,�dJ/�V4�5�M�\DÔD�~���E��n��Rn�~��FVv��8/
�#�}��HpW�	��v����b1	��[�N'�z�n��1A~�M� a�FPq�<���֞�zD$<�Upw�`��w��Em�#}��`dv
���F���P`(����:3T��1��\�;5��G��5W^[Ǭ6��ԧ�_ ��9�%7�w���D���`fd�����4��}���!��W�+��D�gbd�=Y�J1�[�&�h�޵�������Zu��SpW������.69��j/熸�����x߅+,��q/<1z <;n0[����9S-J���T�؆B3����=pK�,����(*�E{�;�G��������_xn�P��� c[�%&�#����n/qQႩ��m�
�����w�4x��_C�p���q.�a��#����x��{�����|?��݊D���Q�o�v�O����f�m�Z����@���X;Y���z�d��QK���Z��X��d)(6�-�HBx�,����1��n)L��x�a���C��k�f�&�`��R�Ps��%���d���|�77�V���R�[�^��v�m�.������>`�SA�$W����{�W��9�w���mO�qY(�r��~��R�<�~tmw}������3Xq�!�ú�����-������i(��anaN������C��}jn���B׸&�g$²#癘��B�qL_x|d/�kj欮��wG����9�.���_ϖ��<w�W"(ZcL��'����&� מ��Wթ�[�ĕf..����sX��l-��N�5�{[�l^s�w��.]�����Ĭ�������������Ò�D.����9����}w���W*]�Ԯc�	�A��Ͷ�b��j@V�m����:g���w�Y&�8A���-�Z��0gD{�P[�����]�����~P�s@�D���롸��TT���q:xz�0(�����Zf%���vr9��t0mp.�'D�ղ*X�� Xl�/<�o6������Ȋݝ�e���`>,�
�j[v�%p!�_�پ��c\��Hpw{���ܼ�=���q�ŧs�1om��3�U�}WaE%K;/\�m�	���Gw�
y]@�`^W�;	?���v�?zfσ�v���h�����Vתj���c#rᧃ��������+p��ΛĠ��}TVL�M��`W1t�ū�6��wܷ�:�.h�3�d���T�פ;��`��+���4��R�����X_?2��"����p�~8u��G�#�לZ
�Z�޺k�ך���\>��Rf׹B�
h�>�/���y�����؞���qCX [\D��w��x��;!�t5��?��1����G%eJ�	�A���~�b��<?�� ��;Y���Y,�_��b;���i6�� j}����Of
�D����D<�0�����&�/��'�_�?	�� ���f�<�nK�q@�����?sS�����9�_)����.���c�uG��S�>)�v��SLd�y�Pu���g_.���9تc\.�w��������p��>�%�կ�t1⣝��7wqK ���dn�G�\�S�J	6{/��7?��Ά�]]C-�h��:�;|{0�V���N��]��� �Ji�:�o��u�Iy��yk|�����x~5n�� #s#��ihm�f�T��/���Ő���J�S��=��g6?K���V��}��m;��˞���w�|iL~�+X��4�T��*�����]�7�8���绎�|��ۖ.4�u���]?�68�D#�v�,����y<Vk�{p+��b����B%�Tk��o��0��<���
��c���V�E�/
�Y@ty-܁'w� ��d{�9��پN��t5���,&HM����@!�o��"G.U_�ƸZ"�u�}�K��N���b�'P�Yv�,Z�x1������!�����^9���
JLp�������`i��U@��\�	޺m��릚�~�ry%��V
��vnH�'��f�b��ݮ�?o��Vϗ���\��?>G��e]�
��l3ۑO���o�i1�c����&�i��-
��5#����Լ,���ŕ?2Ky���������ٓ���Z�LqE<��;x㾛�A���m���;��sF�C�m�w���â����4Ǯ�B�5�8j�Jh��1Jh�V�z�R��1P��^�]on�W*Zc���u~���Ůc�ǩ#!/9��1Zs)��1g���x���X?�A,�P�	�h��~�l6c��!B�Bs�v^�Y>A���U9_,� _-���`|p�$��\�]����J�s�e�Ait��@N]s��ŉ�ы�.�,~x�����s� V:{/����x�����("�z�H�jX	��I	,5ES����������e��~������!�^�]~K�l�<
?]�j�w񠋙�������*_�:�|���OK7�~6�=��˦����8������g��>��D����=Z���b+|��h����'�BߴD8WҲ��l=u~�d=�q�MLt�j��jeL}{	�w�D�/��Ar6E�p����%,x*��h���P�F,/{\�o���Rf�lB�l8y����ַ�t�H�+QĢ1�}s�E��볢�?���o��,$��N��f�o�Xpy�r�S1Y���� ����A�ٞ����_�~?yL�׭E�������߭آ�0j'ǎ��Zu��v���kp�?@tX0�VB�E�m�ώ��QA��������m�f�ѓ�'���>=]���Ҕ)�����{����N!�=��ɫ%�>�|���ݑ���+�����=�i�ݝuB�Z���ܓ��͹��R^W�
돞B~.�U��7����,!u��] �?�x�gB�}��(\0ik����.� O���M��k����w�͸��/6����٩P�ʀ���w���?�Z�GK����zw��^���i�&,�[�9t1�0֙3�<y� HќK����y|j��l��Pܕ�7z���"�!�ժ�y���� d�У�)y�������`�o?;
.���b��|�]�D��2�!7)����ُ����/���'Ak[�W�;��2��ʪkAm�zzXf2��i�?q��_d�r��%�]����ݳ]��n�5f����.��G��~���:7�	�X�4�6�����lp�g�x�,��z#�I���ʖ]��p"�Y<BP�\�?�%$#6R"� 5*�:�^���G��Aa���+�T��������m:~nkX�껔�n`ө������J蟦��ʟ�<���Qh�﫱AP��{��[�݃sap�.�/<�`�MAx�	�s��N�l��B
c�@������wWV��?�g֑�ȥ�J6��D-�'��t6^qyޜۘ�I�����1���o���Vo�)�r Xx�]`oNLj�=\$��%��s��A��u.A�Z����ep�����}�2Y�{�3��Y�U,���~�\�!�i��n�B{ts��/������/���]Hp'��A��f+R9��!B��E���E�v��>� �i�*��q0�����&�]u�JM�İ�F��%�'n�W�vxກ�޶=�Ke�����ؑ��܂���-�MRk	<���֧w����X�����߸ׯ\2ADk �]aP\��<����|^�$�P!��(�wƵG�P��T"$�k�&JH��ct�����A�$F�B���6o閛�1p�������w:A��"�w9�	�F�	���0����iᡡ�ή����&A���9#���'���R��?����������`^�&��Z��('>�R������TS������خM��rcNL�׍���r�q�U���-}�`j^7x��5�s���:��aR�L��	�_.� �JLHL�����k��b�E|���@�=�����{�*�^&�΂)y���U[� ��R܉c�Z�m6ۍު�OU���<o���B��*���1��霣]�5N�\�����<�'|fџ���5�/�K{��=�&¹脤���x�p��V�;,/����g�($����`"��PL��O�v�=h*���AD@���n�02;Fd%C��h���ej�<?a(��l3\.k{�:����p�{��C�Q��A�]�KD�����b�Vղ?g}�P�F��v�was���AJy]�c6���[�-�blP���� ��ڡH��ߧ��Y~�^G�/��ú��|w��y���^l�kP��KM����w�gA�w�-�5G���cg���	�#�^ ���	�s�BH�c�j͑3�k�D��Լl��+���⎓2CZGsG�1!Q�Wo_�e|�&L���,��|�{y��q=����z�A@�}�}'��h�\0�-���N(Ix}rr�+>��E�ٴ�D���;�����
@D�'(H�&D8)B�0�m��kw�w��H�5&�3~�dc�?{]F�09�
�3��G���gH.�q�H�mQ��q�2�<t��s���a�0qŲ���ϕV�܅�@<=f0;��j=��jj�>֩[��O����H�/.c�z?��sB�KD(�N���@#\*�j��/�mO�7tKe�y�в���ǘ��K�J�w	6�Ix�3>��q����y��S0w��k:I���u V;\�5�̜�ڻ;,?���@�k��ť����A,i\D�x�axpd_�a���,�(�o8y��,@h���v�iL4Lg�����_g����;��ˁ�]��}\k�5r��Up��$!/s3�̤F.��h�o*o�\i_�e҅�L���Ut2�+�:�)��t7�x�4��	�	� ��� � �ݠ�Z����U��Ē�'���hâ*92���77mt3<+���}`M��;�5z-֥��qۄ�헚 ��!#6�y��sEl��b��=8~7y8{���{�������v9E�4��ca�P�DpB>*'^\���A����؄爬8��}�XpO��U�͂Ԩ_���־���M���+�x;�����$���=���6:��M�9g*sy.Sj��*����e|w� ��1y��S.��u�J����|��\{.5���쮠e~�r+�͂�E�����a	�ʖ�a��|��pR�����E���AM��RJ5,����,�'�ʀ���G.m�.+5�Ϭ�1�H�i�X\�.�VZ�-傘4,Rc^&�f�4rh	r�U�Z.ud�*;/�������w� /��@f�2<�d�N�߃b�Pa4�_7�ٿ;��n��G���?_�	A�E\(xf�`x���[�9���wa��[<-�A$��Ĭ'�=Ђ�LZ
�|�B�����^z����0k@w���l4�뷏a����:��[��C��U�t���$��k�d���.%36�~d:����P\�m�J��~�`ަ��-g���#'`Z��.Ǖָ�ƭ�a���"���/b������5�<�Cs�M	�W*�྅�]\)M���.8���xa�0xpd^#K\��c������Ѱ�\q��ӎBPdG�m���l���l��.iǇ3�7.���t�d��%�ڤ��;� :s@�jo�f�݊͠%�>����rA���pU����� T֙A+�y����Ǽ-ul�փ���~��傻��Ka-����K_}��ܕG#S=� �]�hr��	��[����7�����MTѲ����h&P�SAFǐ{��^�Ɔ�Ltn}�� <(�=�I
[jn�Gq���?���]J�����<B��(������{�����{���vq�$Ɏ���Oot<.����_`���/����A8Â;�p�N�����YX��)��������,.k�!��0 ��T�|�'���g�дd�k�V�5n�I���Z����������#p���g9.*E�����mw�����'��U��li��*��w��ZŲ�Y���M�������������2��@���E�Y���Y���b��W�j�O8��#�R�`���m���n�76����\/�'Y^�dAR�b�ۙ������w�M��-���ma��"���m��X.�s҄2i_^��of;զ��18f��|9���n�Ӧys_��H�;�a�v	�h�k�iD"��0Yq�����`��\&����U��K|�"4N6P E�>�-X��@�R-�_�5�?�rLy��n��.��	N�Ω8	���v�`E<O��ܜ�>2ã58��ی�,Ք�	�-!r�+�ٓ\�i)�Y���� N�>c���^��������/�9��H�����x�Ǽ��������,�0r砞LP���P��&�|�qq���w?�?��!Fc#ww���E��N	m�;S޽s
�}���7����]Y��9�,.�#W����C��Lic��W��w��p��[X��w`Z"}�&0�QA.��&�݃��s��-�랼��c�*� <$t��~�W
�җ5�v-4  ��|f�ǔ��Cxx���e�����v����e��h�������� ��-����oX\-K����&�	
Y^"#]��q���WiBlG�����.RYY	�/_����FyAp���i�\��\�t��%&��u�߱���.+6�cz������ ���0d�N�w!�k�H�� ?dჷ:Et���*����F.
���G8��, $�ג؎��Z}�U����0'�9��d��#���C��fZw=d��0������b�t�uIU-���RX��Y�����z�Y"�m=��1��WM�]�����u�!%����e�Y~lSO-����^&ԣ�>�1Z���g�����X�`�_Qg�gV��߭�#��+�\�\Y����p���ӁE�C�W���}�dxp�r��w�vD�� ��>�&�w<{�0��o/�U�
��!�?�2���^�,@����{_Ht�����`���p��,�uI����e1]�<�x�O�88}�4���[p���ѣ���+���Q�ŀ�Z�Ks��,X �1sf0��;�ٳg;�G�]+b;�7sQ���k�?>X�VV��v���?u����i\Y+4g!�z�jx���l6��̚5��~��x���7?�/�f�x��7�b�����3g9s���D��aZ��W�.��&	�
��h�p'��a�����J^��<��!��@pw����x��"hp����\��$h	�^raWYQ����u����(|��(D*�b��W��'�#]-�v*��`���o������-]��/��������t{2wtC Qؗt��mꢩ�UE�-�;|>��Ô����Q���PX�P.�f3�>��|�CR�`r�n.�������s�U33S ��x�<=�T[,���5�.�<�E�Vx��z£��^�q�O`����0�p�-~Hw��bk�~p��U&�#�����%�NKq���p?-��ඥ��LlG�?�N�b»���Sh���+V8El�?��S�<y2DG�����⁵~׏�fc�Ǎ))�zvV�_��E���aҤIХ�c���?쇪:��}���0>^�h�r�-����^#�]Vj8�f������Hp'��� � ���Ñ�;A�Ǻ�g���}]^�@�(���R�����VmՔK9�F��fK�ol?s��1_���&A��ߛ�3W,v^{�*w7�cA E�;�[����vM`]�d�a��\?[�r08��E���l
�M��ґ{�{l��@<�*��:�M��w���矁=/C���\%��A��蛔I��(w���%s�+U`ʱ{\���=�@nB<��7,��;Srs`hZ
D2�y�c�8�`���p�c!-J;�3r��]9v�� ����\����ʙ���w����#//������󐓓F��N�E{����5�ߡ���'�8E���d��K�Bs�hю��1XF��D$=F[}]s!(Hc��deeA||������+L�2���HFF��5,���`�镹�;�w���t:�fӖ�Ah��n�y�r� ��t���>�o7�����;~}/|��8l;s�	�(f�����<3�����ڙ�K-|����k�{<E�����3�*EP\A7 j"�߾�Lcw�^Z][�/2�$Z*w�Er�x�~���h,~x�?~�V�.tD��<�Ҷ�����w����=���X����ڱm��喞�Xj	�,�Ā�.�剟�������;�i\�trDVr��Z��2��H�a�7�� �������JH�i���գ���O����K�u���.E�}�����0�fZ��]=w�}7�5�Y���A�\����n��a��@�+Æ�Ç��2�e1D�Y�;)��>|8=z��	���\��q�X�Ւ�l�����,�C�AXXX��L��d����!L:N7���[�3D���F�	�A���b�G?_����K���}S��.���g{��n�=�<��Q���ES|������쀿�p�x(d�m)n�����g�0a�Ĩӹ����;�D8o\@�x�<|w��f݂�2v=��/��w�p��矯�i,jE7��6[��SAMZ��돧]	�Ņ9�_qA貆�
^�	=��3��9���s�\�<�}��`��\�
���k���|
�����^lw�� �ѣ؎�F�ÒGg�����{� �jPe6Ø��Լl��'r\���{�<v����w���W@mPȼ���Y>0?��b]�G�vL��]UK�r���e��6�U50�Y^P@w/t#��q'$��7	�z���H�Ƽ�ױn�n333Y������;��OWk����P�&��L��E��ڵ+K���ڻ�'�@�(�0�P2����9�w�Ðw�hB[1��N�zp���C,�OM`����vk֚'��N^)��R�k��~<�ȃ�1L0U�@�+��n��cz�n,!X&�O��9��j~QqQ'���	(�{�;/�w<+�I��/�}���jb��X@ڐ C#W9"(xr'�\HY���'r��Y�[�|���	옴bq��/,��n������hr^��&BK�������p����e��/�����Gvϛ�'�	�x�o)/("~1g*T������1�U(�WN��\���b^p���{'��׾P��>���sE,��>�_��;�:l)/�3�a�3w���w�G��j4����[Ypt���~)�-~>H��w�D���%M���x,���o�of�:�{;��~)-���7=}���~6�4����rYg׍/y����JHp'�w�h(���v�	� ���WXzi�6���+Z�y
X��&�\�>�y�D:񩵴mR�a#L�=x�&w�X�(8a��\Μ(*��:��}s� Λ*X�ަ��Ի9:s���M�;�cH�c�CwKH�p�(�4��?�>.�T8�&w�f$��B�)�.�������C��Ȏ�;��
���w������̀��2��.���`\��n7��%h�$�P�^���.���B^&	y�L^�M��{�
��J�Yߊ)92���:Fd�4�K����Q�ӏW����׾���;���
���u,���^��:�&Xq0��{65�]�^Y������`�3�����;�j0���	�"m/͕KFl$�u�����6�!Z���q%�o�ܕG;-Q9Hp'�V`��� ��R+%��A+�I��0�w����~�}`�w�0��bm��;v�ȇ ��&����n]�r�"�&w(�i���Wli��p�c��B��ɷ�e���6���o`�b���h{9������).b;֓�'�úcg`��?������ES%|��K��E���Ddp�.ps�,Xu�4h̋���]FQ|w_��G�1fZ�}�g�~�0/�s���=��g���ӻ��s���^\Y_�:�RT0��IcyA+ki�u\dג�.傩�Y�ą���EI\�!hM�;�k4𰴽H�-��=,���`H��C�c�uܵyϴ��	���N���� �=�P�#��#Z)�c�n�&Jc�-�p��'9��\i9���qSV�-�?K7�3c���j�F�u�@��f	V�=*�11�	\���ܶ����t�I����c'h�"����vtà����xi��s[(��Å���E����{�%�Y���|�O���v|��!��ܥ�=�cBKw�/��o������Ⱦ�ܥ`^D���Gf'Ä�L!/i�#1��=PsV��^�O�	]ϡ+4���/�Y�#�nµV�.$����x&X�8	��Zn铭Y�]JS傮q1AWtD�쵙abٿ�iW ��
�q�߻l�Z�PUU��n�w��J�V:L����=z;�3���R�^�G&r��e�r˫��p��%�2�3����v�MH����_�N�cR���0�}PPP��z�/���N!rU2QB�7�R��.����
�#�U���� �A����Sl3��B��k�w�c�i�}�~���#L��/R�����Ne�/-�๢�.��( �B�ĝ;5��Q�xO�]#����0&���Ja��j�:i8�� �	����E������w�3D�i��l�Ƞ�D�5��w�b�Xh�9v���I��z�ݾ�Hp':��j0�LÁ ����3�x{�l6�Ơ� ����V��H��`Dq�Z���,"K�j�]{�<	� Z\Š���\�D; � ��d�kp�m��c,�:��H�~�up��g;���ˠ`�é,��d�փ0�/��"]%�d�A_sk��:��w����zr�D^D+�fp���RaXF������[���T���nɿ;��j�JAAAD�fe��z��y�u�B�w��pG� 	�����0�"�>;��}l�	�zLZ��8t��{6�� �u� � � � o�,(�����'d��D�����j���Hp'����������C`F��d����(����R~�	�޴>�u�;㳐 � � � ��?)+��{I� $���  B-]�K�
�_���e���Av\�2s4<?�:xy��h�!
�BAAA�����UV:^zIVсw���t:�	��ʋ�z�� �O��E{k����_��[�֟8AAAA���eӫO>��w��0v���8�{�*:��uQ	��E;t��caDV
h���hX��t�z�)xz��`��� _���[
�xKi0Xj�f� �Av�0��8��6��兿VN_c��N��WqA��\`w���AA�L�<o����J}?	�D��w)c�:f�A��]�{«�n�`��n��u����p���b ��"Av�H�:f��yk��,���M~��1��>X���C0X#+��������_��u=� � � �� ��'�^y�_J����W�R(�d�p�q�����ԘA�e��~���������'� mPWy1�܁Sz�g5���f�� ������`�؏�lV��Y]��x�m��͋���8Z��-���s� ��vc@���&|� zC0�	�o�>Xx���`���G6[g�T�6{��n�ۭ�j�h�qz#( ���R���35�]o�y�ޯ��_���AF�	 Tð��%�l=��=�ڻ�Cu�`�e�#/�Ӷ6��v�A�����б���/��z;�c����U�'䁟X[	1�� A���������.(|;��/�^}��J�	�ʣh@CQ$����p�cB���{�Ô>������$H�o�Ah������兣�3#�zՊ��BO^�����D�	�����Q�����֯;����?|�����G�&��\]
���E�o"�ɾ*�ۀ�*�7�o�	�,����,k�؈�$��B۪�<G5z��"�@���P�^�Э0<3|	�.���!4��~���z�f�-	=y����!����j�i��A���;� 6�a�i�܏���$�+�0�j48(//��(P��n�7z����#�߆��&sz}�6X��FEEAXXX�c����A!��[�T���V%��'{2�#W�v���p'�s���\j�(�j�d��+�	���/�L�9�]
���6[���ҝ ���n%�� � ��`�� _����L��"�/}��O���$��@ee%���x�7E!�)Z+�[�V�6���7!��q��W#��4���k�۪ �>�3n�
��_n�.�*a��| Beld�NAȌlA���B�;A>�oم����*}��%��a�	� � ��Y㆕���rd��U���	p���Xa	�:�էF�A�mȥA��;����0�{b�?N�;�&�O;A����Z�0P_����t��ǜ������{�F����f��D�g�0�ޯ�h���}7�M�X 5���!�n��AA4��\����|��j^����]��)��<�&���I��p�&�_1h�`�xc��	g��q6Zm�
�� �g`��S({�7��XcP��ݭ=6t�Vk7�q:]��~L`0�:C�@y,y�Y��/��Gb�q�H�Ւ�@�:p���A���ս�h5A�Ϣ}��R�kL){�	U�܉6є�^���ju�7A��,��1|xͯE�ȃ/v��犀 ��R�-;�n� ͋#�N�K�q�F��B��*O�p���r�F��'�	_Ǽx����TZ�ݨ�.���5O���Fێ#v��5[�8�}�2i���p���ho�WHpo��|������?Z�[-��|g�"�Ї5Д�V��)M��D<��Pyy�xB�s�-���x~r�kOnU�DHpW���FmF^�\Z�]zxw�6�w�����>c4���B�Ӧ��:�6�;�����@IP\�N�p�|}!Ɖ���fq�u�v[�A�ۃ8�Dq+::�zy���a�*��]�E���(���RVV���5o�y����-/X�L����Spp��G��}�y����`��m��K���������"��PW�>�9�)�o5E@@ �KK��OC:�}���_���
������W�z�S��f4ٽR��R[[��U,b���$r祮�N�K%4x��§���t�z���_��K��\xg� rֱ�qK�=?44���e�����2o�1O8Ό���u\�P.�K�A:�OF��|�X������'��}�i�S�A���UE��o�h�ɚ��xZ���5�I_�ؑ�'�aQ݁ ���-#!/9:�`J^,;�Ax���.ep<�b�٬�/[�q��rN�O�H�d>���Ĉ���v']8i,))VT�q��JI�K���y���by��������XoKK�<((HV�qX.׼*�;�)�wb^�b�x3/���IHH(뿔^ls����h�l�mh��r�			�/x�1����F�(���f&��x�݈�9�:����V����x�7/AB^j�ܔ�U,�����-'XoQ(Fo �	�O�ǕJ��{��q��[��Z��_>墳�HpW���Xž���VJ`�O�$�!�� 4Jߔxx��~Йxz�`�	B8{�QP�8)�ӚJ
NR������;�7���¡���Ehh�"�"
�ee&���E���h��P<�[��E",���2�((��n,s���x�pQL��� �.�vR(^;9��}	��u�c4��
��b���E��c�BKdo��ϓ�aGAỴ�����bn��ж~��d�Z����5�ZڃXǼ5��]`����u�amʋ�;��6`��ܤ���jFlGHp�3�pWS�=�s����2�O�_�m�D����{�?q����ަ��D{��BF�d��	��"��'D�[)p�U]]��*C)��
�J�e��hY�4�x���R�u����}9]�x�Z!J]�(���`{����J{Q2/���
o�
q�K�*�V-�o��&��hʭ��(Y��o-��=-���!/%�}�Ҡ���b."�w)�q'��m�!T+_�pl��R��t^p�i[w��@S>ePl_���]�1HpWa��Q��ݡ�o�<�˶͵� �F3 Kj��B;	�U��ف��u�+���t���|�C7�V[^�u:�96e0�Yn�	���Cz��N^FmjpB���:�8����'P<VZpǼ(9�C�LP�W���,������٬�;Bpׁ�8�%L��X.�&����+	��ro�wG,��rewR`���_I��ъ��q���y�2:[� qAEJ�,\�Ep%��1%v�S��X�Q.�,�������"��BqW����;��uLI�e��]5�;J��ؿ�5/�vk��:���y��B������5�� | �o���Iq���'����{[W	������N����(�XR�P����%�R�$<�|�+Wl��"�7A���)e�,.�x�\P���TT�BK}o�(�����;�����J�v�8��N)(��X����ȋw�VѵÊ�Lt������))�L��8�+Dz���,1/�@��)�M��8�Xˋ�uL�u�)�����J�1o�ELv�O*�����	� ��A�]���؅`�&�Ʉ���A^�z��[�q"��5����-Z�ykR��N)9�5�7'x�ﾺZ~����a��Q.�̅�`~�%�8v�*��ۛu��I��b����sX�ʿ��v�ɜ��t];�v��(
or���^���J���8�����y���c�V[ؕ�6����r������yJ�r��q���Ѽ��[����>�|�S;AÐ�N����:3�z��Nޤ=�B�K��WU5LZ��~��+�8��Z�&&&z}R��򡲲ڹ��~~�x�S�'�K�$U�"ܥ�b��B~<�/����'^���t���ZSK'�Ҽ �k��䱩���5��a(���;^��ʎO�џ6�_)�M��"�T���˥=��D``�b�����Qf�E�];h	n0���]rw�{��͙o�1-�뀟l�~Fc���o1Ľ�g�(5�#�C�L����_���t��mP�|����3,,��A5���׮����뛿�q�ߚ�a�j�p��]N��&�>������H��ր�RVV&ۂ{LL�jy��2a�3��5m��	�A~L^r�t'#2�{:���Ŧ|�9� ��Y���#��8�>{��,g�F���s���K\���ӻ�E�rIMMo#͋�u,--���ǲ�b�.v�;ssØ����pw�y���r�%11��b��^��ڡ r��gFFW��{mׁ;(���V0/FcH��g]4Bg��n��:�l�ңGN�������ҝ�C�`���ט *99�^_d����v�,ߕ�� IIɠ���PTT$�wy{!W
�k\<��"�H�w�f�^/�?�| �;5��l�#�3Y����Ddp N�?t|�KD��]3]�|�Z-Zآ�!P��Z��28��	�������ǝ��:���\^a�ہ,��[�*�,ko�n�l3��_N0/j�ו�r����:�@�k�������HD����hm�+��BZE������'����O��	�A~
Zv�G���OK�M�'�� �D{��}��P��UC���ȋc;�N���j��#/���i������]� (���f�̀��Z����w\��x?�K���ZZ��U�������p �����/��ڋlr�����x�Z8��W��>���AD#�"Ø����Ax	��.et���Ɍc�o�}��v����b����o%�q�D���F=�]�r�"�f �ƿ/��qG���kH��P^�oW��ɍΏ����O�2�-�u<L2��-��ޕ �p!>L=?sZ�w��"|�|\`�-�Q[�a-RQ�5-���+N�Q5��Qԕ��]��4,��}�{���u	�Z�h���:����o\���!�^� �SK^}j� $�wf��N�	����:�?�
Ax���5��������".��~T.�`�� �ȓD�X�j�E�_,_��*�w�җ�{��I-�PƑ�vvm���aoS�R�x�ue����^��<�=P��S��G!�� ������ޡ�� �
� �D�g6�Z��I�Ů�gF	�B���_y�[ S_ԕ�*�Wm�@�:����)�]����NS�_-����w��Տ��/��p'�V��?>	�A~HBXD�Ќ��A�����V�ک�)a����y�wZQ��Y-QD�rQ7ؠ�אΏ\d�) j	�'�]	x�����/y�x��{�0$�A�!4Fk�mɦB������dF����K�r���ǟw��Ұ�cy}�QOG�����B��y�J�m�я!$�+�w���$�>
G3��W�*��l7�l@�v'�r�����w�}���x_�:&�=��͇z[i(y~�D=ѝu�C�:F4�?�	�W������Q�L8����/Pu�\� C@5�0$�A�!�3��85f+��v*M-}�/N�l6��ą9�Hm��~k�y �U8��X.�,�kAt�!�rh�D��/z�#/�!R��0��lN8�}��$w� B[�-)����B^r<tvL5u@����d�H�)�����n���5���f��kI�.��-��nW}G�\uL����F�E�5$�9v�h�|:�?���'�K^�·�1=�)/�Kע� �,�	� m�o~��'���τ���b���*8��1��/�����)/r ���ZYi�E!���ڐ��gxZ�p���v�?���k}��
�GmUN����QG�_��/��i��;3����R� ܨ�5��{�:2��[pWs��ȋO����ܰ�Dٱ����hT��s�u���KyB��.5�l�C i9��UP���8���-�ƒ�Dj��T'�p.�/��;�w� ?��w��+�@�w�8}�����b(����F�v�����1/8�Z���!r-P�␚�y�l�Vy��5Q[��C9qG�����V�-�2���)���Ý�r)���$��ٷ�_s���MP8�0�h7��\� �CG(�����`���6�)��-���܋:j��K���!5Mt�#�஦�.���-��O3Os)�/"���O�q�ǥ��"5�Ga]'�yG�;��а� ��:��TTAbD(tV��,p�b1���q���QV�c5'�����������b4��W`�4�f{1����r�}x?r)ӡ:��ϼ�^O���) b]US�����=!�d��q�̥�W��C�{']�i��� gJ�;���c�%�Ҡ� �H�G�"�"�%R�Q�e-�'�r	���UoV�� )EM���\�j/<��Z��d�ΰs4U	�v�p�"��a�t��y����N�.6 ŝ ��×�Ẍ$�,=p�+��q��.���	��?h��=�����,u�0�)���kU5p���U۱��&������ڠV8�:�q��*|W5U�@����J��/-:"�!"8 "�`��"8[R��؜�hH�r,�j1�]��r�^����IhhY`�	�p�7E
˪`י�.��9��6c�*.��G�ûێ�!�M1�G*X%y?~�.�7�c1*8��Hg��c��f�m���U����!'!�!&$��k�����^�6�<ߦ��ct�4�Ϯ���^�
�)`�����D">>bbb�������L6���@-��#""�=�!�D�in���U3/(R����񯴬|�)�5Q\<

��� v�x�b�X���Xf��0�����-������@!/�s�F���׌���=\t�Iĩp�~՚kA-�������'O��55��k`0�;�ϳK�.�^�s�s�>�r@��b�0����V�K`` ��ݻC߁�y	�^0�5�w��b[q/�;R�{^��u�9傟��PM���<�1l���:\��E-�kj�%;;�e�M���`���c���}JM����l�'���$22��>YD����-��vYb=�J�f��X\\,�;�Q�G�G����?��8��\��a�3������N�4��L�G��/�9���W:���`�x������CϿ|ŕM��H��P���I-�F�0�'��G��绎Õ�j���L��n��w� ��5��
,�w��+j�؉����	.���d�G�����0w� ���{�]�?6��7�	�(ࣨ����##z�C70����7������[ࣝ�=`�?O�f�
�{^ �]/.��ښZ�����F�5�����V�+�����m�zB�������_�=���\�,U�v��D�� a�b�ŷ����'P���`c�K�2��u�$���NUk欬,�	�3@���`]/L�/���������ib�,B{�&Gj����޷o?�X(�G������g�"'��2�Y�`	��cy���#����=&.���~�y	����`d僋|�Ei��w��6̋��W�:���1Q��}_��^J��T	և�ҠA��c�$������b�/�/[L�z�AVV7Yb0�%%%��_m�?.�b��v�h3�El/:7�u��g��m���m���K;V�����$�lX.Xxo1�i�/��/�Iq�����cQGh'B{�6�ֺ�}LX��^������4꓅d�5�/v��~�ncu��lQ��]4���h+���~�>Ҽ���v���_!/v+�,�����_ay�'�P@Z.�9�m���iǶoU%/�.���	\n�,߇y���R����('3SV+{�M��h;^��%���a�1���VQT��G�Bi��{	�!00-���(ߜ����,�����d���i���
�u��]�(��'���y���#𻥛\����� O=��8(�I��܁�����&��AF��ޱ���Ͱ`o�:��jSW��_�󙐗��9����n�g��Ovo�y��c��=[<�wRl��sZ�n��;�����wfO������\����#80�Y�{��i�d��I��#2,*kj����A���A��&ݭE/����U	�YY��'yAB]FQ$���U�;���9!'�m�����(R*L�-��B�KpPP����@�9A�<X�U��
y)�j����@Tx��߉m&>&�KM^w!�B��(��v��[D����R[[&�ɫ傻7�����D!�\�c����MZۏI��@M�5�u`*�t�a����ܱ\>���."wm��'����RRV���K�po�:�bnk��:�u�T��fu��닇8~		v�5�"�ul�L�O�Џy�\���*����Qż���?�󯬮��*�-��y�EG�*P�wE���q�5S���:���(1.J��T׶m���:<���o�>��(�����U�z���ܫL3��.�`j��Sȍ)7$B1�Mȓ�}_r	_��mB �u����)68�����{�m�K�,��zߝ;�V�2�;+ό����GX;���w����y!�!�᎜����4 %,n3ԫ���}n���uΨ��;.���7Ӥ�W��T�mnT��@��'��>��f�����D�4����pP��Qr��jZZm�y/�s:>g���UA_�?��)h�݅3��9��Up��R��һg�
���iɢ������/���N�8H�����̳��q  =9Y�"�B%���Xa���1����$��0#�MbB?q�Wi���-�^)I	~4=�m�y��LW/�ꨥ���]�&%�ꄂ܉Ya��d��lw�e�����2�9��A�X=�l!��=gi�y۷�-\6��C�ͤ����l�}�&%vЌ����`�5�~o��w�KMN���3/�������n����_l&�������X�fA[��K�*�e��㨿��������3^.F�
g���N"���kz�Q���S�	��U>VV�X����lQ&��5[�Md��&�"!��G�Aw�H��ҏ��}׌����o=vƒ��e�0��]7r%��P}Kh�'�j��#�4,3�F�?�R�|�\_��k/��6|t~o�9NK?�Eߚ4F��<��썃�N�&u}	�_�Z�T�VgĦ�Em���(����	w�5�ϝ���ʇJ+u.��������v׫�
$kM��ʱ�L��m'�����py�x�׾9�Fg���8���y���W�%+\;b��v���5���Q���)��;�s��L������c����6Ս-�[Ew^u]5�y��ܕ	�͞�H2_�d��Q_�x������E]��j[��k���D�yh�Ό�x��J3�HIJ�f��q��t�n3��	gP�lw� E��t���P'��^.t���2��L||��ma�9�e(������&%��V3I]�~um=55�̪���2�
�t�rI4}�p�0"rF�i�dn�z|I0���c¨���sے�n�f+y?����+���03p[��%.���S7#Ut������8:r݉c%/�j�(�g�d�Xiv[X������;�C�;�1�$�E� ,�σ'�\�}�ݖ�g�O�PZ��;���	m���s5��-ۜ����K����<^7m�%����0}i�^Z��-�s�8.��u�Ͻ�'�;����;ݦ1�{��y<�����_?�1������w
&:@Ψ�zp�8��;?��];���K�x{{�qz��<J����l��Ab��b�����<�g���:���>�w��ghz
�7h�D��/�=ۧs�����[�̊��H��"V�]��(���v�)�j�H� ���_�VT���53=U�m�F�;�k��O��2�5��	������[M�������d󃺌��,nK�9Aw(�_?k��ݮ��u�9���ϭ��3:���������`](��� �dR@������]e1�Z.���Q��K�=�,��bƝF��G��X���}7���b� ��x��NU����0����bf�;W�[��Δ@5��hr'��c�걲��Ɣ��'Y��Aw�ï�#Ԋ8�"#�S����;@��g�I��x	M1���no�QK��k�r=ӬhheU8���	�C�7x]�v8�hy���2�,��nC�4��1�a��?a���.�MR�lMC�4���6�5ܵ2��Tr�7xz������T�Ү�m�=i���?�c�O���S������k�۵a5ʨ�4��5Ho��\WmۯY����_Z�w~߾f<�${�B����� �`;S�P�|agU��Ed便Q��Aw�����:)�f���@��0��D�j�����Q�uL�u����*:v���� ����ѹ�t��	bA����D48�#�c5�s�`��"]�`�K:�T[/�B��/��!��y��w��z�D�d�*����!�M����v>[�Pߗ�m7����Ī`�����0F߁ ��Y|�d�>�^[��ǌ��ɩ֞'w����d$�ֱ��;�1Iq��@���E���x�[�k�I�����o�l�D������St���/&�޾>]��q��^`4�P�A#P�ܭ�y���50!�B�ݭ4c�%"��ݔ�л�
����e���^�Acq�=��2���Xzh�xZ��^]�~�`�i�!{��w]��L��M���܀������%�z�����>Ӿ:uV��*�����	������X�N��UO{�_��n�7����rmUI����:/Zd�/�����b�ؓ�n�<�w18��<�!wd��M0�-�Mş�K���>#S�@/�^&����.��:��P��$��W߿ΐ���䄄���xW:?���ܷ^��rQ�r	�]1h�+���]$�ebp�`.�ҽ\x��z�����F��?3g�;��1����pq}~�v�F��UF�kKr��k���q��;ױ�6��D���5��ȹh�[R�������O2~�W��[�����//1ت��O�:���ptm��Xdل�Xw{x�9����ƴ�K{��۾kY��Ovv��to+���--��!�>�)��� ���Kd��9��a�����[��._(^&b`Q2�ӽ-��F�����ü���i�RxR<ֳ���1�擄zeN��0��{_�HB��O8]]G?[���c6E�7w�l��8��j��A�w>y�����g�Z��&�����#��R_�����y7��ܫ5��{K|k�kѺ�����i����ց����Zu�c�d�j�e�O�.֎V�Ҩ��.��ͣ?l+�t�ۥ��<��no��_b� ŗ������{ �I�70�gzO�#�Ϋ�:����L"��Z����k�r�;�߭�H�����z�~���p ��<��"ͽ	F\��̣-������
ܺs=�j�����������*�'����V煴'H�с-j��Ui_szl+D>���Gū-�v0+�/���"~���Ȼ�Y��}9X�~��
����g�&�����p���,S�u�w&yN�
��?v�ƪ�����w�6��������˥��Gk��Ύ ז��3��8�<P���1�����}��C+Â���/�Y��V�����.�}��9����;��bp�_�����oǂ�q��������
��"���NU�Y�E����PQ]�1M������������+�&2���Z�.nz��4�I�sw �F�A�bp6}oJE�����ڭ����у)��6ߊ�&:[{>xXx�N�*jhTvg��[�po��p��Q�it��ܦ�׾����a�3�]�W��L��Q�&>F��A��{�#�%�����{�r�W��w�v?N������?m?t~S}�uځa�;�'�_kqD���e~>c0�q�q+�1�F��Q|�ʸ�c�e^��mq�W[\����{-�|�/�7����H	�Z��g�@똥{f�"���E��\߯G��[��H���#��d�3�)�9#���鱽X��iE�Á�;�3I��� ���������f� �$����ꏨ�ٺ����s��qkw�����\�Iܮ3(u��A4e� �|P%�j�z̵�7:�k~�2��42ս�Z�p���E�*)��޳C�ި�V�ŶSe��p1�{�<̣3&Қ='���V�~[��rk��n�����[����guVy��z��j{�-)�l�   �:�b(��7�H 蝢:��p���N���� f�����>���4~@E���~�e�d:o���\��!�)�tY���2�g!����)C���%��Ր���y#�@,O��W�%���^Y�Z�m���]R��ڝ��r���I�G�΀�,���peп�����;=�Z�=բ1�Vg���r���&�,��Á���;  @ ��q�\G  �Ȃ8b[��G��p��{��R� }���������Ewy���k�:@+6��=���Sz�;gЭ���﷯KY���m\��{0~��}�_�o�R���j��$�4ʦ��);��m������hE-���(}��1���b��뼏�gj���A�5�s���I�����l��h�������Uh|�!=��lé  +,Q� �L�)�sI
s��aQ������k��~���y����t�x�=��f���F��v�	9t�gߡ����9~������t͟KӬ�v��>Q��u�����^6�2'���4s�o]�c垃��6��/I�@Gy��Kjt}>���zK�(9�)�m�Mw_6��־�Y���[�FxL���15��ϴ�g�/7���]��y��镭{{4�V������Ow�</�M�Y�=  @��  a��Nа���p��$rj� �Yt���5���o�)r�v��������qĹq|��t��lg�2�iTV*�>eeC3�t��4.']R��-�ػ�vJ�Xz��Y>Y���mTPZ�1�x����IN�|�h��7���w
�����^�� -�}���x�7+��p�Ǵ1]�ߺ�2=3G�n7;�΅�9�~_I�G��`��,���2�i7�JR��Nw{ϔ�M�{L�9r0��NG�USH$�  `��JqG�; �7s�ɒ��;�;�M��� 2zǫ��s�Ϥ�S�(\���(=���!5��D�?�G{�\]w�^玄��H�~�� �������iw���d\%e���&��Gf^J�5��:�Ӂ�%r�s���9)�4c�@�_R�1P�w��"��w�8�����ee�����x�`�1u��:d��Aq8=�2<3�NU�Ҷ����y��'󮡗��g�n��w���u���`�+�1���m?<[I�!|�o�<BO�0�c�q?��{�Э/�	i;sH2�   t� � �EV�~�T��{_���v ��7�\��(*��~�����<�!��|������5j�ϴ��V�{�zjS�K����;f��R��3�^���GIM����w�i��wRr\��kNɣ�ş����y��;�NGi��y���\�^�|~���bT�c�����w�ߋ�����*|���u�U^e`j-[0����w�#��x��F�~�}�����3{��Ѣ�y�.�j���A��l������{y��ݖݴ�Y�Ӹ����累�S��L&�d��y�|��_����T�N]�\��?�y9}r�4}ZX��oy���m�C���Z��s����YAY,���g�iW�9:Zn'��p���2|]���O��c�������5klk��w����w�^޼�{Zs|jVmr��u� �X��8�b/�J!�^���ho"c�L_�)tkHʺ�!�z��&���,:�zV���@�1>���&��#��)�z'�$�b��k���$2�S����{_&I(( ������}�9�eL.���f���t%�r��A�9����>�^�D����C��23.S��8�qK�o�lw%5�˂pM��WD[x3E�%�Q����0�g���/�8���Mt��V���������5�g�� ���*u�:��zO���I��dH��8����U�ݻ��k�G�)�h�Fi-o�T���4m���K=0y�߿����/�d����<j�?���hڒպ��_ݺ�n�NS����s�����N�s�EG��g�ui܀�:�s�wϢ����o}�9-.9��i� �R�NZX��ѓM�����#�5Z����� �ZJ1E ��6� \��Wޡ�Mɣ��8��{GB��xf�VQ��b� �{��-z�S�G�i��~y��n��{��}�D�vƙ�Srshӱ3ߧ�γ�'������sE�^�K�w�Uc蕭���Z��Uӳ�>���K���'�n�g�O�U��,���P�=᭺�YtR�R艓5M->��$�s��_o�I�{��sZ��������i��_�	2�Ο��/��:��j�xI�(	�K��7y�ڶ_�<�M�\��M����
�E��`;kn�o��:Zr�,���1A��'���1��  `-E�=�  >$�E ��6�Y �������Bzr�U���ydi[�kQ�|���h�����ɤ̮N�O
��n��2����矵r==�Jz`�$�~Ԡ����L�����Uu���Dw�p�z��}!���N�bu>�'KE�MGN�����vӧG��7M�9c�h�������ͻ���]s>�M��N���	Įp�k�Ӕ��&�f��^7��zv�4��<�Y⭡�����!���|�&�n�8�g���i�/�"����m��K�f^A?�y�OI�������؞y����on����?1�*�2l i���8]Fϼ��v�8@,     @ �S�����>M�^� ����6�?��K�w�}׌��g\�9Ц�V�:ڜ��Tz�~jXf-ߴ�>8xҧ��?����饭{�+F���d��OV���_�AQ6�l�$ʨpƴ�}%t��5tݨ�tk�HQ"e\N�(g��H�P��}��;�r��f����]d��w�ܳ�J���kG^B��)�3�R���j�q���`�ז�M����K!d�W6��W��w�yV+hn�������������W7��>8��'�o��l��f�B�2R�Q���Q,�]��A�i������b��tt��ЃKм��NZ�y]5$��g��T�����v��Dz}VX$~�&�չDɠu�<�@���T��v     0�Sn=E �>L"*�=a, 譸�3�~�u�=��4VԎ��{�g����}��?UJJ/�A��R��DY]�ؼ�g:w(���h��_�Y���X�]���Z]Vk����ߗ���`j��ď\��U��F��0^7��.$��1��.|� ���(�/�9J      h�a1M�0')�� zq��'�OFB?�~�`�3f�9Xd���V�'G��S�g��R��    Ɛ���   B�e9]d��a�ǎ��Ͽ0� ����9�ו��%F.�E���h@JHN��S�Ŋ�\2��������4��1��U]P)    �I�QS  ,��#!p��*_|�l�S+��N$ ��%Fx`��2�)     �  Dt�"�}���C���;         \�� ��Aq8ߐd�/ee         �z�6g�v���q�˞8��Ԋu꯷         ��$�~\�tQ�ԨE��)9�SV�[	Y�         `Ez׾���=J�w��%��>��5"i!         ��`TTӿE�����t:�r����      aO�]�  �{KQ����ROw�=Y������c�         �$�p�����"�Э���H]�b.)�w         �Xv�����G(B!�n$�&����׏���      �3�� ����$�u�}bE0��ӳ[�O-��F��D�p         �0�伡n���(�!�>�_X\���K7�$e��0�       )  p���2ќ�%�P��;h�_�Ha��˦v�l�'      ��� ��J۝���e��`;C���|񉳉���C��&          }�Y�S��#G�A�jX�X=�bFj��<��!C       �g7q�uD�ü�+���M��:o����U'Id�w���*)r��YC�dZ�-��fEVZ̚�gW�`"��F�"�6�hg~��?*�>wn�c����x���(
�R�d     xkT�H��P=IR��N}Ã(�2�\T
)K��&�g�$E�%�HTCNٔ �Mq�;l�l76��Ô��洵8��ٔyK1�ɔ���؜��o޺ &p��K[����_��c �r�z��O�Hm�lR�$i&/K�6�²ڝΨ'�yOoq(	N�d�"E�*J"X�/�Lʼ�8+Ť ���A��i�,Ӳ��TC�IY:�bJ�SR�3���cZPHR���כ2o��I1%�!)�6�s7�1oY�V��iJ&Z�B��q���j;�8�� ���~�   K!�!i\��9���R�\�I�T�}v�$��HJ�������q2�D˲�@�M"G���H�Im2�ߠC�,9b$���dE��-���~����$EI��W���l�:*b%)6@s<�+K6uc�!�d��Ԗ\��o�������?�ϳ�S�u��֨�"��R�(�ڡ(-�N:U֪�*l���j��NE	�R8I��	6I�C��w^\мIR��4%��n��N�9��(RZ;b�L	6%����Y��)�M       `���d��MV    IEND�B`�PK
     ^�[�AWv�'  �'  /   images/97fe1122-b934-4e82-b9ff-450ac31bc7af.png�PNG

   IHDR   d   G   ����   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  'IDATx��}�\g���^���:���V��%c9��f`{�a�s`=g��93òs��viI;,qI�����%[�[�[ju���9�7��W��:Jm���:�~�7������4�G������M�XUU��:4��U�z&1�隦�����Q���I���eK�p���ͦ���5�5EA�R���k�	�|��o��]�����~���Տ=��i�`9���&�3�ejE����}D���G��p��\�yV<��k����o6�2��^, Z�N���͊��T-��#��ό��F�&��I�V�۶���ݵ&B�?=�~��)=����+�F</����77��u��yI;�%���ȉS�pjDz�9D�]Q�}h:�^�֦��_i4��OVT����M*�Û�:��T_�ޟ���C�P��1X3Y�Aw�l {^���͚�+�[C�uEX{��.]-���j�*�jEM_� g(WG�JE&��#���.�??|H���5Ժp �z�=p���ڻ�Fo�y/<�&b�JSS�PLD'd�p�l�D�--x��9��FF�r�
M��
�ZZZQ�q'&��}8�n"B	���f3H&�hnn���en���G<>�r1Ϫn���a��y��F�e,�C2iF.�C|rR�2�����N'� 4�B>/�V�C��	.�K�Ô�5�r2n{kz���_0Y>F�XB�&k��x�o�t�_�{���LH"^�����&u�{߇��p���!���g��U!�jMǪ&�2��-&��\�EB���<>�قX<��	�ha�t/�� ��b��L�*����Z�;Q+�184���#��j�J�rCã�s���8�;,4�����1x�l��MC#h��d&�H
�7���kr/L!�B�	9�h
E���D'&��ց�^����^���'�S�i%��!�ji��t��/���Hw�a1�����.3��e��C!3pf��j��s?�)�o�k�Wg[}j M���N���M�������.�O{��[�*��cmںM��R�7c/}�o�I�]w�!}���X�Z>�����x�ͷ�Q��o穓���D�u3���w��'�*�s+׬�B}dMf~\e�c!�޷�fy����[D�p��P{o
�84,v��'��h�.�k�*�H|[p#�G���k��5EhMa�ҟKE�̒P[.��ua��M�dab=� -=ҿ�RIDKezG�>��X��?��C�wG7M���|��E�wߦ��X`��q�V�����hJ����6�3����z]��{��Kg�_}��y]د��&�+�"�֓���ᰚ�����T���)d�[:�p"�Êf�S�ϊ^/[8�}:|N�ѻ�*�a������(��D�^�TA��%b���y�V����hJ�"�F<_B�P��j����"�2���(+�b_<B�I^,�c���U�|�VU#�퍈9,��+�$굓��JW�bQ����\�����3+dMJ��1�_߉YRϞ���6��݅ÿ9��ہ��و�>�G�s�+Ф��A��5��W<O�V�r�JL�H��hcCK~}�.��n߄_��q�ukQ���=r�&�nz�@'��r�lw�����b�$�t�aGg3���Qx���n��N�c�쏴���'ӏ�ߏ�k;p��+����H�I<E��=��a?�9؝v�a�&A&S\n�-�!��2L����[-&¾вw/�|�=z�6����A���FE1k�=r^��������Vu�l�mf�
d�鰒x�TI�)ܝ~�O�V�FO+dM��*�
���%�;s^�dt�tϑ�a9M��\F�w�w� 4�F�89<AT��(d��{��� ��F��1�bI��!�O�3���Ne�`�����Qy��}�D����`	Q��>E��=˖��+ۼa��b���gq��V�mY��hp]�qΎ�Ѿk�p�N@�k<')l�լc�ٻ��%qU&��˄\�n�!���]l"��B��=G@��ʦ�&xm&�u�*1��z��mD�^�_�Ӂ�޿U8�a�����e�����"�YL2';�^�8��Ob-G ��Pd�rYj4l�x��s�<�n�6�`n$�A���1�{���-	!�e���0�9�{)]}9Qi>�b���3�L4� jb�U�e�w�U�*e����_=�L�,��qb�(Y,^+�<]��3�ݱn�,��G��3�&�aR�L4L�<V!p"Gq����c�J\G�P�R`�l|�����8q���������8���pL�3eIH¸��T0��f�'FR��1"uQ�&��c��3�L!����%ƃd7��lZ��'���n�(�V�ɜ�O���~?�������"}`pY�P���6H
���I%H,ؘ�9��#<J�:],��Q=�vV�×�B�YT��lY��9Gt@� @&2�
Rt����H�a���X��N���l*��� *��P<GH��+gp�\M_���D����N�W�U6ҭ����������.�Y�.AH�V�����oF���V7�8E��E&��K1i�H�^���J!j�����0P&�P���3����f�̍t�\���,�>�#�ٌf�È���iQ�p��6�(�}���d���!Dq�<�ѧ"!ǤNQ��,��fo�%�����y��!��G���ԥ�{��/4�����5�}�Oa{��6s����EM�����Ѳ28Q�ua��Ѧ/�RG'�k��Z��5��K,�9��M-�>�K��QIٯz�G�V���ͩ�8K�G�*����>F�Y̰�O�DW���01�C��OE��	����ǘM��Qu�:̡P�~]R�D"0�3yr11����##8% \=u��1$�w��^X)rI��cN[K��v�����⢧>z�N����b�D��}���#ŝ �÷��??u?���h�p\D�l��|	T�\N��&b�-���N�+� ���u���D+�����7�
@��|O��؛NyW,�b�U4����!�Ә!�c�7|
�ɡ9#�J��rd���>��={_|�p����{�(Nۧ9����֐C��?��x�xN@��]��^��A�cQ�+C>2(�!�P!�!M�p��v���y���Ȫ��H*�Ⱥ!�������8���"K3��5KcQ�!�{�����x���h���G^�+d(l$S�k�?����6�����;N;y�q�D�kAAħ��x۹*��H@��H��0�ʂu��<��tG�c��1�d��4!3�����P6��Tw���bV V�"V�u�V|�g����}[GXD�g�v>��+��{wn�k��i���.#���D�,� ~WWI���A'�����R��	�|��?fJ�������F��OW�Q���18F����n� 
Ԥ.�k&��{�i|�/���?��HV����c�0���܃���e�\�>E⥄�Hg�����?;���,R�%M.�̛����֐8{�hqM��C��g-}z��%+�׼q#��7=�o9�*׮xl��1Ό'p����5F��qAS�ۿ�K�^�"~_ϗ�2�r ��?߻EB����N'7U���q�����~]�v;y������Ⱥ��_w�K�����+s���5�f�pfk*ݫ)ߺ�[">4�.I��$��%:"��e�y��DA#�'� P��Y�(�a�3��w�ڀO�y�8���Y##i����x��(9�W�!��?�\����M#�X�V��gmJj�m_Cr�C׺%2?U�r��T��Zd�l��s�%dd	�0�3��xʖJ"nJU���{��HU����leUmN���R_~���v�Y���K���p6�n�X?�7z~���׽��x��9��c� ?�r^�e�G$j�K�P��[`�t���$u6�	"٬'�
�|l>�����a'-�rb"W�w�D���d��ݳ�Du�P&F�B�*��n܂�dB���836IĠ���������,	����fEy5u�\m.濲����oߋw��GPLV<��cx�C	����[�B�g�P	��87ï�����7V����}�n��X;�[���C#r��v�'A�u�a�HN�oN�OE{�����3��0c"�������D��_ہ?��/�לC�zf�|�`����'Ǔ(W��eD���aj���by�O������3�|�T/�����Ș�
߲�U�!��ק�	B��k%��\�XK#˅ƹaU�2��Yъ��\n�����<���4��F��M&�b�RV=��|��ĉ��%�\e�M�u��#
�8��%���:XAN�?��bSsH����;�W���\��0���&E<6�Tyw1�1��_�6���UM~���Z��;��O�$>���N7)E�o�J��л��h"ϻ��m���L�In�f�/��lf3ƲY������QBF�\���ްG�cN��ȓNI8e�s���(>���𡛷#Cz�3���^3Ǳ�KISq�k��/�ǌ���p2m���nx�@���D�4�����q|��$>V+�C�
^��g�H�a�TI��+�X��Ȧ�/�������U5�&��ryO$S������1��������}W���x��riN�S5 ���h6�l� �Pkd�X�+6��[͜�+�մ+��׺����w���r��t����l�J��� �y=bO���ux��lz���W�Aj}�������&�A=�W��	܍TJ�M�W#_,#b7�b��AR�f���O���X����v��,����̍���.����0?�O��<<���ۗ)�̸��x|p+}�R��D��� ���y���18^x��P�Úm�3�cɑ!_�p�۠8=D�ڦ�Ρ�Z�#��x�''A�	"���+Dg�T*�05	S�.m@��l_=>��yӶ=>����ڗ������+#żPPN�d�
�#~�)۹��ۘ�4����Q�j&�d} �*�)\{���\:���Oa���d��B�
��ƞ/��л�ʎ�e/*S2��g��0���c�jՋ�2o<-��,��V�	X��2������<��h�/W��j��JF�^*`I�л�������R��<���!�{�(�k��]�la ���̷�z�}�>�EI��~�0S�x��ev$�Z"dp���n$p:MW�'��fy{��P���[<7C7]�^���Վ�͏W���(U��z�Sr/�b�<�`�<��*�'�N>3B��)k#ߠ�s�z��l�Z��HLo$��f���|�`�� �]�,J��3=(��M�*R�ڴ�q�<�-���2�ym�f�,,�nk1��\;�oEϙ��6l�+�� �\ Q�~脓�'�	�ˍ���زj�+�w��p���A�Vy�i��eR=����k�&��)I�0?�,|`�<��!�.�t��}}*��q:I��/]g	�����gr@��nF@��iB��[|��p��0�"��Z�H�ZQ�@��,�i�P�]�dS�ڼa����aE�<铣1������E�nQ9���b��9&D(�,T�s�3��l�	������Uzn��H�.��Y��ײ���dq����]�gДź�A�d�#8u���KkIE����!��ɤ29�mf|�ݸ��%[�����#,:g<����$��{W��/�Ð����J�3BdC�j-�k���x�7��۹�۷YR����+͕H4'a�M6��gxq���4�������|^d��!|Z��+b�����yZ��r+�o�Il�X�w��R�o��S�NUU��~Z' j����$�)>�������hB6������?yN��.��b?/���)���+Y"�'��&�x��E�	m���W6:�C��2�����s����	���3E�ϧ�O%7�a������u������Sק�#m�T	�JY��M�O_c1Ϣ�3��7�Ğ�frzݢW��W��(�{�5�1���8��a���ȧ$ZT�d�Cn���;���e���K�kπ��F�Tuz��z�׺
3�����=�pR�z�N9
ᲨS��\bc�n^�02�$��9���bW�����{*i�1��)��^sRֵ6�� �?��{I�R��72d�<v�}�$W���^q��6�RW�C;UR܃���ŏ޾���Νh���x^�x��m��j(��I\,;J�Kv6]dŸ}�R�wx5#�59GrL����ᧇ�Q&+t<��}�Ŵ=u�H�
����;ФTH
�(�Z��o>��[�*��[�Fb�|��m�w�ݏ���8K-C���k�H�]ы�?��;1��Sݲ�l�s�l)�	�y�����B��U�\>��U��d����;�~��LW-�����V���ǥ/��+��-17_�6�I�%��K�8��D\�d><�;��d�^��k,6Ik���̥$Lf�;��%�9Z��h�@+�%�l���S��%� �!�,�T\R�a(v��1�l׼
e2m9A�hA�׿�nYl1�iU��@lyr2;uO��e3�>���2
f�SL�������[5a9N�հ��:��l6�ݙ,���b+)hC.؁�dǯ�XJ[�:+���#�/,8�3w��
Ӳ�=z9�+�YZ�dߓ�K��,{���){^����'Y_�93?B��K����W�1Gi5#������kژR`*蓟�6Q����mX�x׵@iQ�!����@o�T��W���T�P���#Y?rU��{��:���LO�3�~ǯۏt[w=s~���eE�Q���U��p��.R¦Ji*
��*sz��7��m̫�n��5��R`ͧ�V�s�VD_����\����u�]�=_٥Rg øn�!##�u��]D�Z])F^�,O-d��'��'�CtB�
���|
w��3�YC7N�KEPn^����;7��� ��ֈ�Ҍ�>7��9'��;/�V�鮭4Y> s��9��m�&��M�3�K7������!& ���J���Gsz����x^jʢ�TE*@(HFV֚ި"��֕�
[&�P��Er�,d=�vs��5��_�_ɽe2x�@s!�+<g�D���YSVw�YY�2y��vh�D�g����,�a�wKN�䦛1�fuÃ��h^4#��K��*��W���kծ@�OR,�t:Dp���c5�jm��iZv��l4N��H��F��J>�B��������"��:2'�?m�y�N���]-W�Kd��u��/�4el2��|zZo#��ԓ�/�x�N�I��<{�]s�G`.�ꈁ�g���R��-JTp2�ŊLSjN�F�,�@y^ʰΓ�+��)�(+��V*��V.����f��f2IXs�9�J앢��U��s����{�|��N�Cz2�o�pS�,D[�p�q�s!@���ݸ��[�"z&��7j�)d���$}!�U�g�wk6ǒ��Ջ�q��Y&ܥ��s�"s�B#�&�R���p���M*�RVO�}�Ej��F��0�6ü�gV���7�i@5����e�éI���8�0
��! .*�00.%p��F&�ܻ�8_�t�ɍ7#JK��r�����r.9HDb��ѥ�q���b��ܹm���\Ɏ����(�Zm��z�%i�sZ�+�h.��e�U_O_<Sa�e-�-k$%SJ��{�l7��DJ*�m�j�ٱ�T�2���"j*o����u�5���N�ry��\&_���7�5�p��u(T�S�f�s���tFb~|v������(lԧ�jE4�t�*�a!�f��o�3��~x�>���͉�k��3&L���_#����c��P�Z��v�c4�Y� T��4�.;���	�9�:.��%Y�S9Y4ƙ-�����Z�f������XmS�	��cؽ���$�Z%M>3�i�X�����ˉݝa�/HI���ܷ}����K�W�^c/���1d�x�5S��v���ӯ̋���R\~]-^V�sGt�>��w�VΑ��͗f=��Z��)bi0�����%�_�Z��_�ӻ&Ԅ�!?~{��C'��F�2����2��� �j��O��a�������Õ{�'�(�,.���h)���z�ń$N]��Z>�ӣ)�vZ���Ta�]���K����Ӆ�,.�5�+��F*�V�i����^���D�{�źA-��4^�V�ɱ��i���u9�Z[�,����\S�Sr�z��IJ�irp�Az�g$��ÓS��a|x����q>�����\A��="�:��?��V�JԠ�<�Q�?Nf��{�z��/�J��_ݴM�<|��焈��C���əd���]�U�)�ͭ�f6*����=��H��!"��NQ_�QOי����!�@oٲ���}�:�o�ح��TY_\��m�����/eߕ��.�)��x����W�HQ��D\L�S�.��-x�� �$�zFcx��v�j�Z\�9؃�ˎwl_�GN�㓿~�|�p�$�Wց�5{k�9n�)^��.?N(�.��jE1+�rqJ��W�\��X�!�qт'��̴�I1��X�a �϶��ƚ���<�{���l���.eEЫ�26�$���M�06���Ef����4,�^	��9[�<n��ph�ϴ���q9�e7)��F�����>�Q>�@��%�lV&����m�wY�z<��?���6y�'��Ғ�l��ہ�Z�x�h�T	��i�JA������G1Q�K=�{U��(���S����摈��xb��N�A9�An2����.���Q��J�p�nΧq�l^If��&�aP��������)�*%����z*y��U<�S�����D��g��7�'Ŀ��wH��9~%)3n���>@���!|*�b�����Rɪz+m]�u�oX�͢dg�9
��ɴ4U��3o��q���b+o��?�SgT�����;�U��U�l���|�R	��F���g��:]d
�%��u{�(����X���S�+�|�ӼN8��B��uY~%(@:$�J��aױ�Z"�nf�Γ����I��rh��:���$4���n��#�j���G�4\dFo�y��{���瓹�g�h���|'�v8?����>�+���l��w���8��}���B]:I3��'n4��wt�$��Q�Ei<kB��?�Q�Z�Wf�G�R�3gΨ����$cQaϞ=�3L��9��I�802xUI���#����عs4Z�ѣ��Xy�ahh###س{��L?�s��7���KL�="3qH)�¹�'�k�n�`��S��!a��c��#.�G��~��Ql޼I������[��>zz�s�ކ@dG�0$ݕ:�plժUH6���i�W�'��������v������H�rE�,g��d�3պ�F]�\U��_8��;Z�q�ļc����?���҂�p�8�Mblﮝr�V)�{�Cx� ��G �{l��رCt
Ssgg'�ڌ�a�o�N.z�Ĵ5s� Q��a����s�Vy������m-�p�uw�]������{��O��@%D�%�}JU΂������~��I���|�����q��]{�����r\�mo�MB(1��H�'��G�]�h&ഋ#���R����6~�ͣ�Ik��U�ں�����T�E~�JWl���׏�FQ5ۙ�1v�EK�l�ѶM_TLf?��Y�0�$����[�_b[2��z_����zm^����Z�S�@c������C@z�����`�l>Dc�*��֧m�ζC"V�����2��h������D!G3y��A2>�� %��ۺ�_��$LO��K7�Z�'����B��j~�D�c-#��"�ʹ�	/��;v�s��O�����m^!�:��b�+�&i�_�%x�� �48��4    IEND�B`�PK
     ^�[x^��_� _� /   images/d5d3b89f-59ab-4c38-95f7-2948dd30f8f5.png�PNG

   IHDR  �  �   �Zd   	pHYs  ��  ��"篻   tEXtSoftware www.inkscape.org��<    IDATx���wxTU�?����LH�$X%B4���4E�"(*(�O���,�����HY��
X@A��6��,Xhb �d`���"�������8��I$7Sޯ��qιg�O�p9�{�0�LDDDDDDD>�h4��; P�; """""""b�NDDDDDD����&�DDDDDDDn�	:�`�NDDDDDD����&�DDDDDDDn�	:�`�NDDDDDD����&�DDDDDDDn�	:�`�NDDDDDD����&�DDDDDDDn�	:�`�NDDDDDD����&�DDDDDDDn�	:�`�NDDDDDD����&�DDDDDDDn�	:�`�NDDDDDD����&�DDDDDDDn�	:�`�NDDDDDD����&�DDDDDDDn�	:�`�NDDDDDD����&�DDDDDDDn����� 44M�4A�z�P�Nԭ[!!!P��� "?? ������t��s����ٳ��ή������ȭ��� 44�7FHHBBBP�n] �����w5���Ɂ�jEqq1�\�b�_�x�Νùs�P\\\�?y&�n$   ��~;Z�j���DDD�y��hذa�~����:u
�Fjj*RSSq��&�DDDD�S�ի�֭[���-[�D�f�P�f�J����8v옽�m���j���C�A�L&Y�A���� �o�w�ubbbp�w�h4VK,����ѣHLLDbb"v�څ˗/WK,DDDDDU!44;vD\\bbbмy�j�%77����HHH��}�PTTTm��2��hLHHp���L�u��ݻ�K�.�������<�����رc�n݊�����uQmڴA׮]ѥK�v�m��K������_�}�vlݺ�.]��|tӸqc<����ի����;�r��Il޼7nđ#G�;"""""�bccѫW/��ٳҗ��AUU$$$`ӦM�����Q�!y5&�>@Q�{�x���q�=�@Q�f����<��0���7��
)))X�v-6mڄ���*�>DDDDD��}����ǭ��Ze�'33ө.   U��


�e��]�{�L�*t/V�V-0 O>�$7n|S_+--���8u�Μ9�3g���]��{�V�fMԩS���C���ѴiS����iӦhٲ%��� ���������W_aժU8{��""""���C��w��7�|�j��ĉ8z�(Μ9�ӧO�ܹsHKK���m�%iQu�Ա��~�-� ,,aaa��ߎ:u��p| ���c�ʕX�~=


n�kџ��{�F��o���뇠���~ff&���`6�����C�!==�
"�S͚5ѲeKDEE!66���7�P�j��~���C�UA�DDDDD%�o�#F�@ǎoh���ɓHJJBRR��ߏ�G�����
"�S�ƍѪU+DGG#66&��~\���|�2>��s�Z�
YYYU�oa��E�ׯ��#G�'���i-���l6c���ؾ};<��U�5k�.]���{�A�v��g�R�~��ￏ�G�Va�DDDD������Ϣ}�������,�ڵ;v����ۑ��VEV��`@ll,�t�Ν;�U�V���!33+V���U����S��z7&�^ 00#F���a�P�F�
�Ƕ���͛��?�ʕ+y[.�C �8.�<.��$��d�Z/�Q��\)�B�!BTUm �h�������H �+�3v���z�B�.]*�����u����w�u�y����/x饗p��V�=YYYضm���{�ڵ���y�%)����B�pAU�K��dJ)���
!� ԔR֗Rֿ��n!�l!��@�r�߇���W�^�ի��
�����X�x1�����~��{0!z��	& 44�B�p�֯_�իW��V;_J� ��!�HB$�~��GW�^]�����ZG	!���n�����ĀY����˗cٲe\#CDDDD7�V�Zx����SOUx����f��_���u� Ҥ����`�Z-8W	a�жm[����� ���� ��s���͛�_�~�ׯ�֭[��s��q����_~���}tռysL�6w�uW�����X�r%�o�UU��H!��wR�M���X,U��Ņ�8�FQ�^ z����6**
O=�z��	??����'ObڴiHHH�ܠ����ȫ=���x��WQ�^�r�����o���U�p��	W��?	!6+��}RR��J�:����p�ު��BDh�3��ѣ��֭[W�koڴ	s���Y����>�G�.w����شi�/_��j5� � X-��"%%�T�|�ڴiӰ����' ��d�I�&<x0X�4)%֮]����#;;�j�&""""�иqcL�<]�v-�mzz:V�\�/����&�� �B|QPP�����n����d�0P1���v��x�:u*��edd >>�~�m%G�}��{���P̞=qqqe��R��ƢE�\%� ��`0,MLLL��X�J�6mB����	!F hY�zݺu1l�0<���ϟ�믿��~����%""""֣GL�2��#�rrr���K�.u5 ��c ����\�͟�Ett�] ��$4���������w�]��ڹs'&O���/V~�^�	���ׯ^y�r�Mۻw/�Ν����Z�B̷Z�_V����"�111=�V�x!DO %����[��/�w��e�>��*���cѢEݨ������\pp0^{�5��۷�v��������"33��b-�f��ת�U/1115UU`���N�:a�ĉ�����:/^��ɓ�s�Ϊ
գ1Aws5j��o�Q���ܹs�7o6oެuy�����?WE��-66�NUU_��Pj�{LL^}�U�y�e~���$���K�靈���ǵl�������l��/� >>Ǐ/})_񑪪o��қ!�PL&S_ ��u�f00p�@<�쳨]��AMRJ,]��-r�?��b��ƚ4i���痙\��Sϛ7��A!�6�����b�Qձ������ ��j�n6W�����/�\��+W�`ҤI��W��IDDDD7��ěo����@�m._��y��aݺu�/����o��}��<.�!��dz�t ю��ׯ�	&�;���o�a�ĉ�|�rF�Y����v��a���e�w9q�&O���\�^J�*�x=99�����]['3@��)�����o�}��.�[\\�Y�fa�ڵU%�!ƍ���~��v7n�[o����UU_�X,�,H7%����C��s ��x�����o�����|��ӧ��s������P=t7ԫW/̜9��M�֭[�Y�f!77ױ:GJ95  �]w��V'���W!�;p�Q!0h� �?�̳+W�Z���xN�!"""�rF�ӧOG�>}\������ٳ�F���:�b�l�� =@DDD��)R��p�zݺu1}��2w����Ą	�g�=BukL���ȑ#���ϻ��,;;�'O�֭[K_��`0<�i��W��m��)**�.�|�b������o��f͚�|�M���믣��-�~Q%�U�.\X�)I��ɘ4iΞ-1k������iǎ˯�8=ITTT��(K �����&L� ��a�������
�-1Aw#cǎ��ѣ]^?v�Ə_z�G����?���<Ytttw ���ꂃ�1s�L���.���/�`	(((�� ����H7�k��|���(�m֬Y�ٳg��ٯ��S�%�ʃ�Pݺu�t�� ��a���;�����ѤI��I)��[o��>�)R���!��+�`РA.�lٲ�'O.=����r`JJJr������)����:EQ���b�ȑ.g-�ٳ�?�<����
������P��d��G�c�̙���/��������W9j^1��>��VנA,X� 111��Rb�ܹX�j�NQ�&�n`	>|���.�C�1�#2�:>o=
�{ ��y�L�:�唛��D�=�I:���[�.�-[�29�����/��;J��%�a6�������i$�\	����h4bƌ�ݻ���͛7�|�!�wJЕ�x�^x�er��*fΜ�9s�8&�yRʑ�����ߘ��䏤�� �}��3f���5����~�eODDDD�v�����]&��ϟ�SO=U:9߯(J[&�7�l6_hݺu!ě T (,,�k��Vf>a����O�0I�ύ��9�ƍӼf�Z1y�dlذ�^'��(�|�W�5�jmڴ	-..^���.**
������6oތI�&qww""""S�F|���0�L��O�:�g�y��fp[�F��111J)W�e�5j�{�9����bҤIؼy�^!V;��W�>}����׼VTT��'�H����k����۷�laa�} 6��,F��K�.i��gϞ?~�NQePs��q��;v���J$�Rʥ���������M��> ༭>B||<�t�U�f�*s�}�:>���i�ӧO�ܔLUU����زe�c�>���511�^1���f�n��a)�
[]jj*�y����k�gذax��'u������n�ĉѭ[7�k'O��ȑ#q����9)))�l۶�X� }��b��`0t`?�j�ʕ�;w�f��� ��_�B����
���=44���F��5[r�i�}@B�F�������z��KV�^m���!�\j�;r�H�k�_y�t��A�������<��<x�浳g��g�AZZ�c�����Wu	�G%&&WU���2�V�j�*������CBB��{�!88X��� ,X� !!!��gϞ]z����� ��T�իW[-�( Klu���Ǹq�PXX��^Q̝;���DDDDT�L&^}U;�NOOǨQ�p��9{���L��a�XN�n �����}�ǫ�h�3f�py42U>�O��x�DFFj^��O���Ǳꈢ(}-��.U:)�LII��lu			�2e�暘��̛7z�IDDDDP�^=̟?_s�jAA^x��<yұzfJJ�l�$$%%�QU��?lu���ضm�f�x #F��+<���	z߾}��#�h^۲e,X�Xu������l����2RJ�~��Ä�mu7nĢE�4�GEE��_�->""""*��f�B�ƍ��I)��o 11ѱ�����7t��,�UU���.�}�W��~���=�bcc��gym���^{M�����1e��c�2TU}���'t�Jضm[����_��{luK�,qy�àA�p����mРA�ܹ�浏?��ĞO 6�nݚ��T#����Q  ��������ʕ+NmfϞ���:��]Q����l�7�q#�|UU�X,f]�$'			����� ��>i�6m�;��V�iӦ�nݺz�IDDDD��v�m.g8�޽.t��+����ի��G.��� F � p��yL�4�q Ӯ�P�<^��2����S��������r<�9w���;���# �T&L������4p�	�CQ̘1Cs������	�%�����l��5Hr)99�� ��V���_�x�bͶ}��E׮]�
�'y]��1c�h^�ꫯ��?8V}����.�Q�Y,�$ /��G�����5������w�N�QiC�ATT�S��S�NEzz���*����x\���|F�q�]��ҥK��o�i��2e
��W!�KЧM���� ���'ObΜ9�UG���F�]����% >��?��s���O�m_{�5ԬYS�Ј���蚰�0�;V�ڧ�~��۷��B��)))�Q�JHH(B�\�4�7�@VV�Sۆbܸqz��3�*A�ի:t��T/����ӑ��k�*B�5555S� 麨����2��;|��7����+kҤ	F��""""�M�4	���N�'N����k/!v�j��-=c��c6��	!���z��g�b޼y�m�;�C��|��$�?^{#�/��{��q�z�l6��%0�a�%[J�7 V �x�b������p=�#"""�i�۷G�nݜ꥔�1c��B� �pS8�g6����u��W_a���N�E�+��!�����IЇ���P��.��w�q��)%%E��mr;�e������/�������ߟg��Ė�iY�fM���If���XrKF�� G��[fΜ��as\\�w�wx^�+����1B�ڂ�T+ 0ZJ)���n���� �Wo�f͂��� �{���;<""""�ӷo_DDD8�gff���s�ڝ���D���%$$䪪��Mu?y�$V�X����^��`�3<��	����5wLNN�ƍ�e!�����z�F7/!!!���ѣG�v�ZͶ�>��^a�$???���׼�x�b�]���#��·j�[�X,� ����,Y����;���?�gh^���z����'�Լ���c����gu��KNN�`���h�"Ǚv;v�]wݥghDDDD>��CӦM��?�իW;V-LII��n�Q�RUu"�, ����5ۍ=~~~z���<>A2d��Α?���f��,�|�رc�z�F�K��" �r�
V�\��nԨQz�EDDD�3E��O?�ym���(..����:K����Y,�� ����ׯ�����.,,���ȣ���@<���N�RJ,ZTb�])))_�U	��|HJi_ôr�Jddd8��ر#Z�n�klDDDD��G�s�?z�(6o��s!�t��rY�ب��p�z6�|��n�С�ѽ�xt�ޯ_?���8�oݺ���\�qQձZ�3�@vv��+��gXDDDD>a�С���/��ڗ���Y�懺EUf�Νy f�ʛ7oƑ#G�ڵl��:u�34��	��Ҽ��'�82����%(�r8`���z�j���:��ݻ76l�ghDDDD^-::&�ɩ�ԩS��Kt��y-�#/�����I��(����5�q��rxl�~��w#<<ܩ>))	III���(���GSe�B ����W_}������<�ޡy�h֯X��q��|VV�R͆�RSS��Ͷ7n܈?��é]ǎѬY3]c�F�����_���O?u,Z�f�f͆䱒���!�c+�Z�������s-Q%FϞ=��333���:V-���^i)�K P\\����?N�x��G����xd��x���ҥKغu�c�|�p�y�wl/N�>�ݻw;5h֬ڵk�kPDDDDިO�>�''mذyy����B�=�Bf�9�L���k���{�1(�G��n�#��������N��|�M�����?�50ҍ�l�'��a+�]�V�]�>}t������[=��C���K����f��b"}]{���ŋ��O?9�iԨڶm�wh^�c�Ҥ����?ORB����MU�e��?��#�\���������qy�F�!&&Ʃ�b��89IQ�=�bf�� �n�����^�z��W��A��Oe��ߏ�'O�˪�~�g\�?)�j Y PTT�~���M�:uСC�C#"""�={�Ԝ��a��������E�e���Ν;5�z�����kP������O��ys���,)))ɺE��b�dK)����{�vݻw�-&""""os���;թ�Zzpd%�~�~����qm��j����������.�C���w��ũNJY:Aw�V����(kl���݋�/:��ԩ��1y���`���:՛�f\�Pb���F�u�-!�o��j��s��z��u<*A���C����>��g���B�/􌋪Onn�f ��'����S�[n���v�ޡy��;j����?:S���:5"�$�Xm{������l�6L�o�G%�qqqv�߱þ�7���f����qQ�IMM-Bl���o�^��5󂈈����*�*���F�`�-���o�\=��_uj����W��Ֆ��FM7��)�}nͮ]�4�d�:"""��Շ��?p��{YU�MN��k%$$���Vv,�B��}�<*A�:ޡ�� ����(
o>FQ�� $ dgg�8��&66B�C#"s���    IDAT""�X!!!w����_�\zÆ��P���s.�t �{P�<&AW���N��EEE�������y����3 �Y��}��ڄ���E�:FEDDD�����48����?o۶�y�"y5!�O�קN�BZZ�S���8]c����h�Bs�y������Y�EnC�����g��d2������Ҭ7�͎E���V�Z�d�ʥ> ��o�z��<&A����5�SRR�;5��SUu�����YU�V�)''G��������[�z��}n��c�����n��'��ذ}�.���Q�~�HKKÕ+W�ڸ��3��Sjj*TU�������(!D����Ç5�p���yL���	^��ϝݐO���?��VNMMuj�Q��I�&N���XG���M��>�Y����}#<&A��A�ȑ#�;Hgff�5(r			E ��)�n4@͚5������#���knW����Ԁ|���hZZ��ӝ�4o�\ט��G$�B�'x'O����R;v�X��q�{�R>}��f���P��!"""�T��L�N�r,rṗ���`��K}6 ��}#<"AoРjԨ�T_jz�qC"7�(�1��3g�h��M�����|M�6լw�8�و|µ��N�V�;,,Lϐ��G$��r�f��s���A�8)�	�kW	:oDDDD���K)K$�R��:�D���V�;((!!!z���<"A�W��f���Xt�SA>EQ���.\�l��DDDDD��3edd����^B�tjD>Ea c��rxt�^�(�4]�!wf�+dff�j�:5�<"""��խ[ש��&`B�?��O�R�s0�c�����G$�~��7	!�E��!�T\\|��ZJ���L�6�A�O��T*+0��9�DnIa�gddh��z�C�yD��YY���z�C��`0\r,k�P�V-��!"""�TZ}�R��{�����V�`��zyD����Y��`0�����������B�6F�Q�x����<�V�۱����)������\�r��ct)%����e!��'�|��R(��������ADDDT>�>S���� ��6�t�]�MЋ��q5��M��rn�A�����c B{�[kp� ���]Qn���bYn#���E�8DDDDDT������wEr9��G$�ZOc���JW��@���h��'{DDDD�'ǥ�6��o)%��)e�}o���w��	��t�ι�8|*�v�����4T`/&�������^��@@���E	�+rO�:u
`�C���O�����ʧ�gr�{�-r[B{�j�	���=;;[��v����R��z�C�)''��g $$ĩMVV�n�y*���c� ��)e��:u�h�a���xD����{�LQ�$|��j�������DDDDD��3���6{�|�����[��f�+W���7����/��&��jC��!�d0�O�����6d�NDDDTZ}��	Xff&��>�"#��_�H�]�R6,qOh�K0�TUmn{]�a�'xDDDD���3թS��F`�S�텫�7���	��s�4����쯅�5��B���v�l8r�Y""""�?�?ީNQ4i�ı�Bǐ�=���B��]PP�˗/������;I:� ��� �T��̙3:ECDDD�\��BCC��^�{�u�������ٰ9s���z���<"AWUU�)^�f%f�DDDD85"�!�����iӦ�mΞ=�[<DDDD����Ӛ���o)�z�C���ŋ �k����{_?�H��ԩSNu-[�t,�ըQ��n�[B( "m�R� W׿dff��Gr����c�t	�ܒ"��:$$Ds�ɓ'u��xL�����TW�N4n�ر*Z��ȭ���� �V���۝�>|Xϐ����<Vzz:��Ҝ�K��ZEEEu�܍=A��{�9�ͣt��AQ�vz�C��n��u�A�Nm�9�kLDDDD�Lkp#""B[����/Vנȝ�������l���yL��j��d�sf����^�۱��'R�ADDDTqZ}�ڵk#<�~���>J\}Jc s��lTU� ���ȑ#���u���-��.�S�N��EnCa�ǡ�g�.%%E�x����<��bѬ/��b��bbb� P�V���sjs��1�����1	��j�����꣣�a0lE����.�F�.22�>�[�M�6Nm���������:$&&j�;&�R���Üw�V��~��F��>� �o�>]c���@RR�S]PP"#�wCQ�^z�D��h4����r`` ���6f������JKK�<&�]��>5����:t#���\w�}�f�܍��Q	�޽{5����k)%t#��i{ݮ];8�q��!""""״�P���%֡�������sW[�s�Κ�8�~c<.A���w��ҥĬ����(�C��+8� �![��g�n�Νz�DDDD�5\��J���%r��t|�5:t����ĉ8s�ޡy�J�

4���y睨_����(��z�E��СC]4 !D��6�/_�����������ܹSs�����X��Ԉ�����ѨW��S��۷��7���e+��=z8V=�Ԉ������uTT����ر��ω���n��+Wp�������11�����Q�h۶�?�Gm�^��W7�رC�����%����!�t�/��hk2�"��W���2
!�	��Ķm�t�������lݺթ�`0����yCJ���1Q�(,,���9H
���I����ޡy�K�ϟ?�y�u\\7n�X�7݂�j�(ʣ ^{��={:�����/���whDDDD^���׬���wEEEq7w�gϱڴi�F�95ضm


tʛx\�h�$E����g[@1���^�Dǎq�-�85���y� """�	�N�Ҝ�ޮ]���+�2BϸH_&��1�>�r�~�4�mڴI����G&�7o�\Sܿ(��Gj\TTĵ�^*...�}N��k��������x����EDD��-(ҕ�� ��V�Z��W��ӱ{�n�C�*�������Ņ���cǎ����%=�"�X��p��۠A�w�}Nm��Ҹ�$Q%X�n�����}�Q���'�֮Q��p=�"}DDD c+?���pj�~�z��	U�G&� ��_j�2ıxWTTTg]"�DEE�0�V~��'������믿��j�12""""�t��e���N�6,�]1n���C#ԨQc0�[��K���n�ڵz��<6A�駟����T߱cGDDD�ˊ���g\T�Ey@M ����ڨ�����J�Ј����֚5k4��X������% ����B�I�����_b��ٌ�G���7���j����?w�B`ذa�U�cbb:�U���� �l�����N�:N�~��'�>}Z�Ј������ݻ5�V�Z�^f:�[�n���#:th0�V�����5ۭZ�J�����&� �z�j���:�?���hѢ��,�|Sǰ�
Y�֗ � @@@������������H)�r�J�kc�ؗ'Cq���'����N۶m�UU�l+w�����N�Ξ=�~�A�ؼ�G'����o��E��Q��z����rjH%666�x[y���hܸ�S;�ł��D=C#"""�	�ׯ�\f�Ν���I�϶m��U�����B���c�j�[�b�~�$��WGJ�v
�ӧn��6{YU��j��TU}�֞׬Y#Fh������(,,t9�����;yܴ��h�fC����uL����~�L&�v�.]r��7]?�O�Ϟ=����(x��W�"/_�<ʩ!y�������G�����;�ۿ?~��g=C#"""�)�}���(�w܁�z�^�R�rm$y !�4!D ��������[�.]���|]c�f��WGL

����nt���^�R��M��t���OJ�>�}^�6m���zJ��{�)�������,[�L�ڄ	l+֒R~�[`TiL&S[)島�SO=��͛;�KKKs��?��H������g�i^�8q"l��V��_�F��ҥK/���'M���;�۳gv�ܩghDDDD>i͚58s�S}���1r�H{YJ���d�glts���! p���g�yF��E�4J��yE�\E�x�S}xxx����L&���!L&S$���r���q�}�9�SUs���12""""�UPP�y��i^6l"##�e!Ģ�m�6�+6�9�z@[���^s�aw��A|���z���&A�����E�4��1�[����DEE��ݘ�m��!> ������[�f>�gxDDDD>m˖-ؽ{�S��`��o�	??���M
��ݐ���6RJ��p��{/�w��v�ܹPUU��|��$� ��W_�b�8��n�����EQ�	!����6���3���_y�4j�ȩ]zz:.\�ghDDDD >>���N��[������3�L�G�[����)��? F 		�ԩS5�nܸ			z��3�*AUUӦMӼIDFF��g�u�z�d2i�ڙL���l+w���>��f���x����]�����˗k^{��gK�%�X�F�1U;UUhe+O�<6tj������x=C�)^����Ç]�$�����;VM����G\Tqqqq-��q��٤IL�6M��Ν;�n�:��#"""�>��C?~ܩ�`0`���

�UՐR����t>+����d'�j+0 ={��l�K�.�����z�8z��S��(x뭷�) V��ĴrjLբu�ֵ�V�7 ���h��o��ڵk;��������������`�ԩ�����K�����_1p�@�^�Q�L&�}B��xdd$&M���v����b^��`�ĉ�[�7h� ,p\�^OJ�]LL���f�������� D��&M�Tbj��Y�f��ٳz�GDT��F#a4������`0���(^�O6y���D,]�T�ڃ>�!C�8V�9x����Fe���n-���֝׮]����<��ʕ+�2e
��z��S��d����Æ�K/��ym��՘9s�c������;w���%8r��������w9�}Æx��t����� +�R"!VB��u|�^�@! �p�^ßF~~~�m*BJi� ��j/;�QUV���ŰZ��Z�(**Bqq1�����*�����"�Jc0�b�
�����b�={���I)_NII�>���\LLL#)�. �W�-B�N���J)�������;L]�FcBBBQu�xy��(
�}�]�{ｚ��~�m�X�±ꇼ�������C�T�bbb�)��g�:t��ŋ��;q��|�Idgg�#�?!���`0��k{mK�m���$�f�L�^�lI~餾��EEE(,,���:DT��M����?�\������C�����UI ����?�3Fڶm[���p+�;�2e
�x�	��+W���ᘠ�v�����ЬY3�k����_Ɩ-[���_���m۶9oOU"::z<���r˖-�b�
;��������q��=C$�jfK�������???{�1	��i�_/UU�#�EEE�$>??(**��<���{��{�iޓϞ=���;n2�
!�2�͟��k۶mPAA��B�.��#F��_�l�w�^<��3�'ey&�:kժV�\�5j8]+((���?�ݻw;V���7�#�U/::� o��M�6�'�|�y�puM��M��
��tb0����Ѩ��kͦ�t���W���>_\\������#77L�����ѣ1v�X�k���O?���L[�U��l�D� }T۶m�m�Rv�����S�N��7)--��_q��E]���jеkW��_��|�����1c�`�޽���?�5�U'&&f���~}�F���'� ,,L��G}���U.[��� ؓrO��,ޞ��ǖ��F�

������|�E��n����?��Ci^OII��Q����c�R�7���;��M����'��Na?w�{��/�G�MAA�~�i$''�gu`�^M��4.;;cǎERR�c�O����X,�u	�Gt����ҥK�!\�ƍ�d��h�B�=7n�k���"7�(
�F#jԨ�+�/'�Z|=A/�-y�M����Evv6w"��>�qqq����ۇ�{�q_!	����9z��+bbb�"��  �VףG̙3Gs����?~<�mۦg�Ն	z5��?����������\�7��� �(��PRR�a]�rQQQ���3)�ö�f͚ᣏ>r9r����ѣG���P�8��l�S�m��q�&��϶���{vv�汪D�BBB�駟"<<\��b��1c����X��h4�v������ƶWU�[ �mu�<��O��rۜ9s�j�*�B�vLЫ��(�1c���y�v���?��X�&�����曨BL&�m��Y��s�>���s�łQ�Fq�v�j"�@@@�}T<   5j�М
Gׇ	z�Z�(((@^^rrr�����y�&M�����7BCC5�>|cƌAZZ�c����dBB�w/~�b��у ,h�<x0&M���ߠ����[��3A�f��୷�>�y]UU��Ǘ~jdB�LNN~Sr��u3�L	!V�k��С�ϟ��[; 9r#F�@zz�^a�4��`�%䁁�L"�����*��������v�j֬Y3,_���LZZ�}�Y<xб��b��lޭ�&r�ڒҙ ^��	!0z�h�3���V�Z�9s|o�t7��s��p���O?��o�]��ׯ�F�3|�W1QQQFEQf ���}�����믻ܙ955�F�r<���*��(D�5�8=]_LЫ��Ҿ�=++����Z���O���[�d��Izvv6^~�e�ܹӱ�@J9�b�,� Y�\[o�
@G[]PPf͚Un��{>1Aw��`���x�G\�ٻw/&N�X�h�?��O���l�� =Xtttk � ����F�?�v��`���9'�D��5j ((L�t��8Ҟ�������牨����bɒ%h֬��u)%�����w�-��p��(Ó��������� �# !����p,X� .߷l�2���;:D螘��EQ���c��.ۜ?/��RRR�%���x%99�J��Qڶm�_XX8�T8�wiҤ	�͛���(��MHH��q���&���#00��9A��ݽY�V���#''��ϯ��-�܂?���_\�ٺu+�x�dee9V_B��������%�L�fB�� J�<>���1c��%�RJ,X� ˗/�!J���<'Nt����j�G}�?���Ӽ�R�SRR��K�n.&&����C8l\=cq�ԩ�S����n޼���:�]'[B��5kr���`��YlS�sssq�������4P��R�vm,X� �ڵs�������?�����җ�*�2��,4���{V1@-[}@@ ^|�E4��5����:u*6l�`&�n�w�ޘ1c�F��6�����ɓq���җv������*ctW���a��N0��)G�Z�0i�$<��e�ɒ%X�p!;;D`4��xPPwT�PL�=��EEE��͵�e�x��c41}�t����eUU�l�2|�����-�o�������r>J��y睘5kn��V������/��}��Uu��	����Ă\\=�mٲeX�dI�#\T)� ������X�ATTT=!�KB�9^�ڵ+&O��ƍ�x�ճ�M��M�6Uu�D+((AAA�i�f��ga��}
����+W����KD.!0h� ���K.7��'Ob���سgO�K� ��h4~����[�������6R� J<���1c0|��2�
�	p�ԩ��c0Awsu��E||<ڷo_f�`���0�ͥ/X)��孉zddd}��P��ZӦM1q�Dt�̯֭q��	�?G���H�<���?j֬i�Ä�;1A�n����\�r999��[k߾=���Q�n]�mTUŗ_~���{W�8mu^1����#oMԣ���0@_8�� ݺuäI�V��X�n�O��%��0A� �����;F�U��Q)%���;,X� ��G���b2    IDAT�b���_���[�4`��L��E'�|@M�k5k��ȑ#1dȐ2�	 ��0k�,nG���Z``�=!�r��ݷH)QPP���l\�t��T]"ШQ#���,w�,++|�>��ҳY C񉪪o���x��B�L��/H)B�ļe˖�4i:t�P�����Ü9s��_Ve��	�����[o�����2��o���ŋK�f�`�U���{DDD@�5B� �ḱ��}�>�(Ǝ�������1{�l�[��
#&ro�� ((���

*��y'&�ͶK��+W������D�ئ�O�0���gϞ�ҥK��W_�j���\�[ �Z�n�y���N�Ylll��r���o Z����#G�_�~��E��~���8q�DU���{���`�?O<�D�����\|������O]%�� �K)�Pe��lv�9oݺu�x�b7!� � P�t���@���#F�@Æ���;w�����q���*��Ƚ٦�ےrN['&�䨰���ٸx�"��hݺ5�|�MDFF������X�d	���;�u 8`�����_��������~~~� ���)�ǈ#��#���f�z_��㏵�͢R��{�6m�`ڴihѢE�m�a��X�G��\���!����~_���cbbI){!z���[�9ްaC<��0`@�Ǧ٤��c�ܹX�~}��L����5k�F���&�䊪����222x�	�,����C�b�ر(����U�Va͚5e-�<%�ؠ����������fVj���d2E�)���> �Yw\\��nݺU�!bb"�|�M������b���0d��9AAA�W���Y��7o.��q ; �R�Z�V��;w�̻���u���/--�v���VJ�	@g w���uEQйsg���]�v-��p���f�,\������!???�(97w��0A����������/jM�%�zM�6ń	н{�
������͛�v�Z$&&�մXJ��. ;�X,Ǥ�U��$""�v@@�I�A�@G ��j_�vm������GDDD���ŋ��{��o��ҙ���4l�/��~��
w³���u�V|���صkWE��X���!, �I)�8�(�EEQ.]ڿ��M�m۶u�Vk����B�� �	!Z���!D$�H e.|B ::�z�BϞ=ѨQ�
�� �g�̙3���~�'���Gpp�=)'�(&�t#������ũ��ڷo��'�U�V~ω'�i�&lڴ��Y��r B�Rp\JyZJ�&��TTT�~��A�s�u�旑�Q�j��SU�>��B�B�Rʖ�:֢�o��]��W�^�ҥK�f Wg�Z�
K�,�&�7�	�����رcq���_WG+##;w����۱c�\�|�fC)`pS�h���p��w�s�θ�{ФI��zrr2-Z�]�v�LDn�h4�V�Z�Y�f�g����n��jEVV��Ґ��_���BQ���cƌ�вSG���;~���ر����rq��}SS�BCCѥKt��:t��eq�����믱d��;w�f��iLнPdd$F�U�u!�TU�ѣG������$��f�>}Z�5g6DTT����;��xJJJ�ҥK������;���,�|�sj_O�K��3=3����(�"|�B 1�D��̦��(���DB
Q	EA�BD�%A��D�(`p@�oc�3�����3�/�Wu���~�:t��z���S�}I-�]g���t�}��}��B�D�F�6���]ש#Щ������8��}�{DGE<��#��G>����c��b��W^yW�^ŵk�p��d2�S�t/I�099���o~�q���:-��J��o~����Glll�B�Å}������ ~�w~��[RZ���}�6������lnn"� �N�Z=�׏(�p:���|�����Ν;����C�廮��h�?���_�׮]���!�E� �l6�n��n����q0��ii4����b��{rXQ���_��_�>���-o9�sE�Qܺu�n������;�+��F8�N��a��������q������d2����O<���&F�]`@N��<�ȱ�:G.�C&�A�\޷��`0�d2�f��(���D��o|_���92���`����鼫�$DGŀN���H����%����x�{ރw���p8}�F��t:�B��|>��a��j��`�,�0��}m��M������H�)`@2�.]�o��o��xǑ���\.���������˗/�+� ����g>����	�H���*�_�λ��5��mz�SSS��_�U��7������/~�WF�YF�?�0���wᡇ�ۣi���xꩧ��o~KKKZ�3�Ї�(�x�ߌ_��_������:o�M�x�<�~���駟f�����_���eh&��ʕ+�я~�z�	tҒ�b����Y���}N�r�N��f��?�����~��v�]��R���x�����~7o�Ժ����N ���1<��Cx���7��Xc�N����]���^z	�/_���|WՑ6�1�g�Y\�|?�я�:j���0�S��V�H�R��b�!GM�$�w�}x���7�	�.]:���Ǳ���k׮�ʕ+�|�2w�i��Z
����_��?��Ә��F(:�7p�dRm�q��-���+�s�0�a	�F7n���~�#<��s��B���kEA�TB<G:�ֺ�S'Ifff033����i��7���c~~��������/��@�#�����2��v��r��tB�e�t:H���
 (�J�T*P�L�T
�t�LF�D���ɮ�4�}mm?������+cS����zY��@.�C$aC*:��###�e.�.�K�&�I=۞�f�(
*�ʞ���x\}ｽ��Z���o��K�s�z\�R���2����.����r9<��s��w��s�DD' �"j���4�����D�(�� ���8i����Z���K/���}�{�v��<u�N������E�P@$A.�Ӻ,"��ĀND})�J��?�1�����XL�r�����b��3gP�ױ�����-�%"� t"�����W_����=���|SHD�I��3��R	�X��刈:������k�ԤR� �#��\.kZ�e2�066�p8�Uu"�b@'�}�k_Ӭ���j����f�������v��
loosj�11�QOivv����""�/�SSS��jH$�F�Z�DD�Љ�'8�NȲI��.���:@��!�����߫՞5LDԓЉHSV��,�n�k]
�A�t:�t:Q,������DD-0�Q�5���\.�F��!"�.2�����d2�H$�uIDD=����F����rA�e���u9DD�!�N���χT*���mv'��ǀND��h4��v��p@��!"�"�n7�n7r����yN���:������1iDDt$6�/^D�X���&
���%u:u� �Z��z�0�LZ�CDD}�l6��ٳ�T*�����Ύ�%u:uD����^�׺"" ��V������Z�DDt�Љ�DDQ�������r"":z��P�@ �x��߉h`1��]�$	.�n��ى��+DQ�����E2���֖�%u:�9iMEx�^x<�R)lmm��hh]щ1�ё�t:5�sT���6Y��N����	EQ�.���1�сt:�~?dY�9����P�A�+�DԏЉ��x<��������W̉��/� ��Y��J�����z��uYDDGƀND{��������O�Z�2�Q�in}w�\H�R��ND}���  �\������o~�bQ�r���Nl��fP'"�e�DC�T*ᩧ��7����y��!""�8Q��x�r����F��ND=��hH)��'�|_��ב�d�.�����5�{<�b1�b1�K""�C�t�oA �2�� W�4�����Hc�Z[[[H��Z�BD2�_|��u WЉ���fC �^�g8'"�����066�`0���5�""�1��Ʉ@  �٬u)DDD=G��cjj
�Bkkk�T*Z�DDC��h��|>��v�K!""�y�.\@6����g�Q�1� I��v��v�yƕ����v;fff�L&9������h�4�z<���u9DDD}Ku4[4e�w"�
t��p8������5Q����`0�ǃ��u�r9�K"��w�D}�d2����b�h]
�����8s�
�VVVP�մ.��:Q��$	�n�[�R������bQϧollh]t�>#dY����9s"""���n8�Nlnn"�Nk]t�>b�Z`0�.���h�I����1����T*i]�9t�>������9Ϝ���LOO#��buu�FC뒈�O1��0A��z9Ϝ���4�ooo#�Hh]�!t�e�����.�����HE��ax�^n{'�cc@'�1:�>�N�S�R����.�;w;;;X[[��(Z�DD}�����\.vg'""� ��t�n�cmm;;;Z�DD=����L&�A�L&�K!""�E(�XYYA�Zպ$"�Q�D�$	�.��M������l�ŋ�H$����u9DԃЉ4�t:���!I�֥Qy<8����X,j]�t�.��t�iNDD4��z=Ν;�L&���U��!���N�E��@���DDD��u���X[[C6�պ����#��w�w�.�����Kx��ǵ.c�1�u�^�G(��bѺ"""�1�$arr�\����vJB�x����k�\N�g9�"A �2Μ9�pNDDD��l������Ժ"�WЉN��hD(��4""":2Q1>>�B����e��u�K"�.�
:Q�	� �׋��I�s"""�+�333p�\Z�BD]�t�2���DDDtb� `ttn����DC�+�D \.Μ9�pNDDD�\M��t���t�b�v""":m� `||�\+++h4Z�DD��+�D'��DDD�M6�333p8Z�BD��+�DwA��!�f�i]
Q111�L&���U��9��{*���� (�����������x<�������k���������Ѻ��ǀNtLv��`�$i]
1�Ӊ��Y,//�P(h]Α������|'����ŋ��ZG�Z���7o�ʕ+��w�����S�-������O�uzQswi���$IB0��n׺"""" ��?���B"���֖�����������?��:��.]¥K��|׮]×��%<��s�\)�vx���f3&''Ή����� �׋.@��k]�>6�������/��ἕ��_��W���~��h`q��^�^�W�2����d0p��ylnn"�J����o�6}��=�k4x���w�5�B!|��_����]?�=��#�x�"����X�c�K�Љ������j�"""�^'�"FGG�t:���EQ��k=fgg�|�$��|>��կ"��s�s��9��?�3>�� �Nw�����-�D-��vLNN2�Q_���x�f[���S	�M������>Qd����t�]DQ���,�Z�BDDDt":�gϞE4E$��k�c�=��s�5�B�=��y�D"$�I� �˅��<��Cx�[�����9|�A������?��ӿ������!t��Njss�<��e�1����d���HO6W!"""�[~�v�KKK]�+>66�}�Cm/�J��׾���A.�k{�O<Y��я~�}�{۾G���?�'�|����$���WM���A���A� ��nLLL0��@2�͸x�"l6۩��G?�Ѷ��c�}�Q<���G
��t�����mϚ;�N������j&��4�$I����~?Aк"""�S#�"Μ9�P(tj�a����w���c�D�>�(�����/��2>��"�Ͷ|�=�yϱ���1���2�����ls"""*^��Ν�$I��-�T+����˿����]?���>��O�|lbb333w��D����������$�֥u��lƅ`�Z;��=�P���;���˗O��O=��~�閏=���'~~"�1��PE�p�p�[ډ��h�I��3g�t�#�����������ޱ����������:�DZaw����\5'"""�A�.�F�Dϥ��066��󋋋x��WO�ܻ=������F0�����鎽�V��NC��trK;Qf����
��9dY�(�W�^=Ii�(���^zi���؉�:4Q
�Z�� """��5��_�5���o�կw8-?���/���#?�N���l��ku,�N���qȲ�u)DDDD}AQ<�����?EQ��k�Ng�����N��G"�h��v7	��:$�ٌ��ɖc>�����`sss���?�L&s�_�.����t�,U��Щ�1����e�����������n�R)<��cG��nU�V�u�, @�Ri��Ә�N�ML040A@ ��v"�k�F�z�F�F�Z���Z�BQ��u ��l
� A�Ǜc%IR�,����Ծ�$AEH�A ������!E�s���j���(�>��Oڙ���W�Zř3g�D�����Vv����l6[���Ŏ�Q71��@��t�v"���J�RA�ZE�TB�RA�VS?�ժ������u:t:���?߉�5�����R3�7k�]w�F�(���t�� A�͏�M��?�h�	��`0�͆������E���`bbb���v{�kj�����Щ��f���pK;�(��(��(�J�G�s�P^�T I�F��O�^���� �N��N�f��V�G�5� @���	����E�i���z]���j�?���fÅ�����z�+W��裣���UC:EQ�uf��1�P_s�\����&�hX�J%�E

���A��a�h4�d2A�e5��U<EQ�i�00{nvX,�FH���fh�����<������Yx<�}��jw��َ���9���r�_���Щo�\.�� �c*�J���j/
j(���z=�f3L&�v;�F������h4��
�H���$i�w����	�N���W��}�މ�O2�ć>�!�������^�x���}�������u:�I�022r*G��s�A<��!�ˡX,"���[���t0���x<�X,0��0��-Wf�w��u���5û�dRo�X�V�F P�5{��w"�M���_�*������^;;;Y��N�;�ڒ$�ܹs�>���ܑ�'�:�������Mi�^�cgg�l�l;;;����VEEQ��b�,˰Z��X,�X,�3څwI��2f���C�!�<O_�V�4�k7k����?������O���&Q�ַ�O>�dG^��a6��}�ƍy~"-1�S�0���y"��e5�7��j�T����t�j��a�d2�_�Q���M� �h4��)�7rv�T��j{{�R�6y"-//�O��O���~���w��]�������jG��HK��dYF ��{�.j�������A��l��f��nW9��PE�п�^�W���M�z]�ͳ�\i'�L&��{���'155����m�D"'zI������|�\��������0�S���|�x<Z�A4��,2������Z�f�6������gt�ժ��	���Ps���fS������zsϴ��J��O~�x�߼o� ����8���������k׮��;t�Y�("���HD��(
��,R����j��WǝN'��QOPE=��� �~����v;,��s��h�R��c�*�
WىN�իW��SOa{{��������y晎��Щ'��z����Q�4�=a<�N�3�wEQ7��}�~Q�����K��ժ��Z�0�L0�L ~���2J�;Q�|>�F���t�9� ^}�ՖgͿ���w�u��ĀN=�h4bttz�^�R��Vs�<�H �H �����    IDATN�m�՜U-�2�N'9��}��o@Y�V8u��؝N'E���x�����p�ܹs�}�vGn~E"|�S��@eD���z��b���h�1D�^�XD"�@<G2�l{޶��W�eȲ�-�44��:x}K���"F�Q�p8{��7W؉�x�f3.\����E�j5��!�y��3�N'�� �MQ�^G<W?ڭ�������Y�yt��gj��z���n����Q�l����(�(�(�J�OtDz��ϟ��۷�ȍ���\.�~?�9�!����h�D��9r��։�F�\F4E4U��7�H��N/hn�ovv�':�$I8w�������.��g1���� dYֺ���h4�L&����Q(Z^'�v��m�sȉNf�v���u��f88�N�l6��n��e�j�RI]]'��DQ������՝+D�:iFE�B!��v�K!�)�z�D�H�h��=Qa���r��v�y���5W�#�t:�zl��p@��z��z��v45�
n�'z���Q��D'D�	I�022�U>���V���b�F����m;�����	����ͭ�D��jH&�H&�{n�5���������۽'��;�B4l�~?�z=���;�|>��(2�S�c@������5z�J��ۈD"H�RmW�$I�����������h4���º 0��0��jX/
�Dx��^����҉��� ������c@��ǀN]e4166��_z4�j���(���l��\)��|�e������ ���w7jlv�w��(������4�l6Ν;�;w���A3���}�S'-�$��Ʉ��1nɥ��<S����X,vh(w���x<�D}LQ�}+�n��,�K�M�\.���^,�i��f�;w����~�˲�}�C�4�Щ+�V+FFF8hh(��x<���MD�Ѷo8���}>ϔ��+�$��m6 ���l0��������h����q�֭�}XdY�����GU��"t:u6��p�ᜆB.����&677Q.��^g0��z`4�X!i�^�#�#��`0��r�����v7����(
���T*WNt��z=.\����E�k����:�*�Áp8�uD��Z�"�`ss�����$��v�����tv�B"�E�J�H�HD����xԝ4�$�n��n��Z�"��#��q<4I�0==�h4�����x�{�˩?4T��Ը�n��~�� :�� �bss�x��-��~�.��;I���fg���MȲ�Nmh����eN�S�_,5���􈢈p8�����G竫����8�ʈN:�
���ϧuDW*��������χ��z�|>na'�ci4�u�����ǣN?�}^�^����ZM�ʉ:��h�3��{�1<��m�[]]ŗ��e<��-Ϯ�t�(A ˲֥u��(H&�X[[C4m;���Z�r��N�DDw�\.cccC]U�z������$��p��p�YUo�=���(�������?�<��C{c0�AŀN#�� ����8�j�����"�8EQ�J��J�Z��?���UuD����J���~+++��W��o}�[��@��:��E"����*b�؁+Q6��`n��gˉ�+v���\.���=gtw���Ed�Y�k���(
���	��������'�4�Щ#B��9��z��H$���ed�ٶ׉�Y�
��l5%"��ћd2	���׻�fa�z�VC6�E.���w�k�dn��x\�R�N:�� ��*Է��"��ְ���j�������`0����
��V(������-u��^�W��tp�\p:�����f���N}+ C:,t�k����VVV����
��v���zZ�ZE$A4m��]Eu�z�P@6�E�\ְb���P�("�jR�͛7�����kߍ�vR�a@��"FFF`�ٴ.���EA,Ý;w��d���t"��ru�:"��ؽ��f�!�;�f�X`�XP�T��fQ(����J   MB���Z�_��:� ��jպ�#���������
�B��DQ���A(ڳ�DDԯr�r��f3|>߾s���N���ԩ���H$�u)DÀN�"�"FGG^�/T*���buu����$���!�|9�b����Ulnn�c!%IR�}N=��!��r�4��� �40��Ț+�����"�ܹ�����`�A�=oT��U�V�����(�^/���y�(��p�n��A�����~�����-�K!:1t:��s�s�e�`���q�M���p8��@'"6�ђ�hT=ڳ�� jC�|>�L&àN=�����hp%��:����r9,--akk��`n4
�̉�~FQ��q$	�\.�B!��=�X�VX�V
d2��i���CQͺ�u:��z�q����|>G������J��r�a2��\���^,��dP�T4����@ �F��9�Է��@�p��z�������l6ctt�3̉���A�U�L���ٌb��t:�u�9�`�� �Hh]
ѱ1�S[�pv�]�2�T�\�����/3�9�]zcPo�������4ϨS��PH�:&�'贏 �p8Z�B (�J�}������z=B��� Ϙu��ު������KA@8F��@:�ֺ�#c@�}� �N��e�\.cii	kkkh4m���t���DD���L.�L���"���<��r9d2�Q'�	����1 `H����N{�AȲ�u4�*�
�ܹ������I��P(�P(�9�DD]�h4�F�L&�������l�Z��f����9�+Q7���rg�tR�|>�s�T�^���*�ܹs�RA���0::��y��Z����-�b1��}=?A����fS��AG��N� �����Ύ֥��  .��G�2hH5g���ϣX,x������,K��#"�vj��������r��<.�"�N'l62�r��F�Ұ7o����
&&&�.��-�$8�N�ˠ!�H$����ڵk�s�͆��Y���0���fϐ����!\�$��n�B!��f*$z}A����C�%�!g��
��.��P.��իW��/"�Ͷ��h4��ٳ���{9Y������y,,,`ii	�Je��z�>�~�_7x�n��j��'>���ԳЇ��jE8ֺ2�r7n��3�<�X,��:I�0>>���>����I�R)ܸq-�}�L&�B!��nNߠ�+����?�3
�K!ڇ����l���(R�4����駟�����͂|>��~���=M����(��H$��^{�x��56��p���恵��<������ݩ�0�!�����Q�s�d2�g�}sss� ��l��{p��Yn}$"�j������C>����(��e�P&�I�
iX��i|��к�=�І�^����gFSW
\�vW�\9�s��`��������.VHDD�R(0??����7ku:�~?|>t:����������h]��}�H����1�Lҩ���XXX��˗�*�"��0��~��~no$"�d7n�@4my��l6#
��t��u������/h] �A� `dd�A�Rh�E�Qܼy�R���&''92��h��u���#�ctttߔA���T�ͼ��]�rO<����7i]
9�! ��0���R�����Cg��t:������w�2""�U�R	���p��ݷ�]�$x�^�E�R)6��S��o}����nb@~���z��4����֭[��P��|�����B""�#�L"�� 
���k6�a2��������'���w���l�{��&�Kpn�.�K�2h@�R)ܼy�l���,Μ9�EDD�Vs�{:�����f�Ǜ���f3R���F�Ҡ�����۷=�Gt������Ӻ@�j������8�:Q166�`0�F?DDt$�\sss����B����r9��i4�*�A%�"Ξ=���y���c@P��P���:�8Mদ�8Ӗ���MQD"�R)LLL�܁e����t6��NE�Ν��ܜ֥Аa@@F�###��Q�r7o�<�	\s�_ �� �H�R��[���z122I��<���\2�d�/�(�^���iܺuK�Rh�0��N����}?��N"���^C�R9�:Y�155�q~DD�Q�x�Lccc�ey������t�ͽ��L&&''����u)4$�Hsֹ^�׺�R	7o�D4=�:�N#"��V�Vq���\.����"�"�n7�f3Wө��v;�� ����.�� � 	�B�:�ݭ��5��������̙3�FDD]�J���f1>>��t��χR��t:���q�l6�K:�\.���U�ˠ#�;�����p8�.�@�\ƍ7���N�$LNNrR u]�VSW������k��[,$	��SG����\.��BZ�sd����}�} 8x<�ˠ�Dp��T���s:�8{�,Ϛ�����p:��7�L\M������:U�}�9N��$*�
nܸq�YsI�011���DD�3j�n߾ݶ�{s5�d2!�Lrn:��(�H$��EQ�rh 1��1�^�qjtb�X7n�@�\>�:�ݎ�g�r�9��x<����:l�X`2��H$P,5��E�����.^��u)4�xۧO���qjt"�Z���
�^�z`8E���e8'"��V.�������(���qQ����v���I'R,9z�NW��T8��hԺ�S�L/��2
�י�fLOO�b�t�2""���D"�f����lys�f����� #j'�J�b���uo�!���W��������^84��|>\�t�ᜈ��R�P���\��*:�~��es9�����@6�պ �}F�e��n�ˠ>T.�q������ G�$LOO��ٳ��GDD}��h`}}w��i�y[8�N��~��v���C'��}��Ʉ@ �uԇ"�._��d2y�u���w���@I�Ӹy�f�Qk�qlf��˕� P7o�� ��>���0::ʎ�t,�zsss�v�ځwvA���(fff8ۜ��R�R��[�������f9����[tl�z�o�ֺ l�A@8�N��]tt�|׮]k�Z�d00==��ޥʈ����(
������099	�^����
�^�x<�Z��A�ԯr����
��.��W��@ `�.:�H$��{��p�p8p��2��P�f��y�f��^��P���ض������u���{���,�Z�A}��h�[����������V�V;p˻ �z�p����N�r��6���ƀ��L&����eP�(�Jx����r�uz�333�""z[[[X\\l�l6� �ґ)�r���v�{���qD�Q<��3�d2^�p8p��%�|%""�eggsss���-7���NGV��p���ˠ>Āރ���JQ���㥗^:t+���W�V����h4��qQ��zy���,��bssS�2��0� ���;�t�j���ׯ#�Hx�(�8w��nw�*#""�O��`}}�B�����kY�F��x�z]�*��D"��v6�#�
z����Rt�l6�g�}��pn2�p���k������$P.�[>n4�+�����ۼ�CGƀ�C�#=������{�b���N'��^�� ""��B���mG�I��@  ����ʨ�(�����ˠ>���#DQ���H˭TD�Ͽ�_�~�Ю��p/^d""�h�b�D"-�����P�R	kkkZ�A}���{D ��hԺ�Q<oNDD�����Ŷ��m6t:��8GkQ[�xN��C�R��q��8�����z��h4�9�)i�Ko75�d2!B��w�2�'w��A�VӺ�a�k��$j%��^8����f�ys""�SV(077�B���q�N�@  ����ʨ_(����9�ˠƀ�!�;�������ի��e�x<����{""�.h�KO&�-E>��ۘ��j����U�ˠ�d��`0�s紏�(�y�&���(ʁ׎��bzz�7y������h`yym��e��Ψ�D"�T*�uԃ�$N#�,��*�S�Vq�ڵ�w�DQ����^o�*#""�7�D"(�˘��d�8:���e��vNݡ=���ш@ �u�c
����Cù�`���,�9QH�Ӹu�V�#ilG���׺�1�]&B�ge��T
�>�,�����Y,�{ｰ�l]��������177�R����f�8m�7�T*<�N{0�w����dҺ�!�H?��Om�p8p�=��`0t�2""":�J����yd�ٖ�����ω+�O"�@.�Ӻ��]d�Z�r��.�z���
�_��z�~�u>�333�$�K��q��u,..�=�&�^/��>����S@ лF��!
i]�����#uj�8{�,�E�EQ���������Ȳ�E�CQ,..j]� �.h�;g�F^�r��u,--x� 8s�&''�Su�������>n�����x�T�|�hT�2Hc�]�r�`�Z�.�z@�Zŋ/������E�ϟg�""�>�Fq�Ν�[��f3�@�m4�666P�T�.�4����d2���i]��R����T���t:fgg�����h ��i,..�mk0�ӒT�6��O�(���ܺD���x����֜q�1jDDD�#��aaa�j���z��!�T�Z���Z�Aa@?E~��#�;;;x���Fm2������""�T*�����v��$I�|�H �T*�vd6�Sb�� ˲�e�ƒ�$�\�r�Y"�ł{�&��K�Q���e��ϣX,�|�9+�����hp1����Pn�hW�^m{��f�avv�w̉���@�Z���B�co�(���qG��h�Ν;Z�A]ƀ~
x��677q��u����s8���������u�vvvZ>.�^/{�����i�0�w�����к����
^y�C�$y<���p�
�j4�}�6��t�k�n7�v{��^���̭�C��v���8�z�---aaa���|>�����h@(�EQ��FcϿ���5�k4�.�浍F�F�$A(��NA IDQ�(��$I������(XZZ���d��.�� �]m��p��-\�pA�2��;(B�$�� �ܾ}����^���q����&�A� ���`0�����������^��Z��Z��V��V���o�{���Q��4����5_�Z����Z�k���{~/��C�[�!]Q����43��B��x<�׫u)t��;D�e�b�n�:R�@ �3g�t�""jE�$�F��z�F5���z��e��e�J�=��T*�T*�
�ij�����#]�(
�ժZc�ZE�X��Ύ��i4A�=�=&�	&���n�4����.�ɲA��d�\����u8��#�l��Ā�z�~�_�2H#XZZ:��`0�����/�hȉ���M�Ѹ磹�].�Q(P,�J��^.�5������v�����������34�L0���D]���
 mC��� �[���(
nݺ���Y�K�SĀ~B�  
�Mː�������ׅ�a����~ADCD58��f�FX,�=!�\.#��#�N�X,�T*�X,e����7��RE��bQ�s���{�� ꟱�d��b��b��l�y�Z]]E��h���p8 ;{�r�������!Z)
�Xu�	ɲ�9�Cjnn+++�^�pNtrͭ黃��b�ss�P( �ɠP(��ZMê�� �Jy�+�zp/�J{�<�J�Ҿ_o6�a�Z�|��5��[__G��@0l�x��;C�p���|�2�(������|Z�Ax�װ��v�u###�BED�十�d2�y�\.#�N#��!��!����ijo�����硽�g������X,����l6��+�Dǳ��	A�NbH^�(brr�H͉��0��@0�
����;R8���DG I�V+�v;,˾�WEQ����f����\.�j��a��kwhoޠ�������n�4C{4����6��v���O���.J��    IDAT�A�nwgH^f�n��dR�R����,˰Z�Z�A]���p�m��`��ډڐ$	��C]!߽��(�Ƴ�,r��:/�z�$Ip8p8 ^��W,�������������Ύ�2�\e�e���c舆���:Ah�k�n�CQ6�B�P�t�;���Nǭ�C�֭[G��ح�hQa��`���p8`6��]S.���d���%��#��������(
Eٳ���uN�S]�]jD�[[[� m��7o�1�Q111q����?��B ඼!s���#�9����sN�b��n��n��Z�j�L�t�L��n� �9�P(�F������Q��5�|>����&DQ��nW;�Ұ[]]� jO�7r8��/�cC��>8Џ�yn������p�|>�sZ�(�j���t��rA��ﻦ9s���y�/�(B�e�c|�\F6�E:�F6�U�j6uG���*�z=dY���,�\]�����Aڎ�j��bX.cccx���su@0��$Im�t�`Z^^������y�^LMM�C1�^�vdEQ����d2�T*��nԒ�h��h���Uϩ7wV�>�P�V�������v7��U3��\���˲���� �"��Ǐ�'�z�1��~6�"G
�.�gϞe8��`0 �2�N'l6۾���g3��,9�$Ip�\p�\��T*��O��@2�D2�T�л\.���}#����(X^^�(�p:�-�i���r]���b���K��K0w��`����b�<���M��۸q�ơ�9LOO3��@3��Je�s��z�t�D�L��d�#v�]m֛+��l�����lp���x<0���N��(XZZ���t۩Bn�[yH���^�_�"� �9�#�w��H"��+��r�9�ł.� $�NY��v�a���=��Õr�va=�L�k0�ﶺ�
��
�����m�4p�1==ݶ����QG��+���W���}�cZ�B'��~^��?؇D:��K/�t�
��l������@�$I��a��� �#�L2��&v�����H���ξ��ͮ�+++p:��z�p�ݼ�J�^����۸p�B˭�ͮ�X�rY�
��~����~7FFF�.���!C�N�4X��,�^�zh�0�x�"o���hn	n\*�
��8��(��QOEQ=�^�בJ��H$���m��H��j��@ ��k4��*p����!]E�|>D"6��w����Z�Aw���`�狇@�X�O��Cp�t:����\#�=�^�������^�#�H ��0�I���z��zQ*�ԝo�������`���E ��u�k�J����p�B��}�(���#��;B�'�੧��o��oj]
��8�ζgzhp��e\�r�ЕAI�033��ܥʈ:K8�N�|��[���<��(���S�2�L�����z�鍽E*�
677�����������ԗJ��z&��n���H$���C��'�����vN��C�mp��p�����Ozh�Ap�����R�zYs�������h4�N��F��d4���t4gE�\.��e�b1$�}+��� �� ��pU��Z>�������Z�h��t��|�F���1�j��q��_��֥�11������ l�5\�v�H�w���xV�������k��[*�����x<��xF������H�ӈ�b-gD�^Uw�\<�N}'��`mm���-7�x<���N���v��u�?���f3��^{�x����������P��I������v[[&����6��t��#Ҟ(�jS�b��h4�d2�o5QQ����dB0���gx��x���`���˅d2��ʨ۾��/�K_���e�1�.]⭳78s������Eܾ}����~?����P����zx�^�������:b�"�J����j��d2�h4�J���:I����
��>�����<O�ǛG;h�E"D�Q���i����/�Ę�����������~�p�r�p�̙.TDt��V+� dYn�x�ZE$a�^���z�|>$�ɶ7���:����D�v��ٛ�z���*C�ƠN��z��q��m|��w��t�z�Z�A�(���^;�:�Պ��iv�e��<[*��;�lDt4�(������ �� ��.�� �H �H�n�#��riP1��E��۷q�������n7j�wW0Q166���%�K�#`@�����l� �����k�m�b4q��E~-P�iv�m���r9lll�|9�	� Y�!�2r����������l6���yX�V�����r��.��F��;w�����-'y �����F��;|�X�VX�V��y�K�C��ϘL&LLL���*�Jx����;,I�瞶w��� <ρc���,677̉NI�X���R�ԁיL&�������=��ł��Ϸ]�h��T��U�T0??�u=��Π3�����dێ����?{w��v���Y{��*��z���X���B1�pl���X�L1��#�(O����`>�U�<�&����`��H�䥸_v��F7�{c-�Z3�Ь��}QyШ�s����{;��:d-������i�Z���~W��}�9e�0E;cԐ�R����J����urr"������X���ddrrRFGG	�a�b�(7n��x�^����&ǯ������)F�� �0�bQ&&&�����ߖ���k׮u<�S;0�|�r�r���}YYY�T��Y���	�h�1���err�����c��<O�߿�"�KL
�{~�뺜qc�?�
����	�a���a��������2s b�\N�]�&����Kj��,..����LOO���0uDjssS��l�������E�_�)�uerrRVVV��
:�� }ddD�ɞ��!�666daaA9n``@�^������ejj�c󷣣#YYYa�9`�\.'7nܐ��#Y]]�J�r�Z�&sss���&SSS244�L��s�Z�ѐ���g�0�J%��ڒZ��Tp��.qO��r��uV�c���@���(��r9y��7Y�Ad���err�cc�YYY���ݐg�<�}!T�M�P�+W����@H3�+�Lʝ;w:�8�}_�={FS'''277�4�aR�{O�SSSR(��.X�Z�o���J2��|�4D$���LNNv�^4YYY���-����ۓ������J��\�r��C�l6+w�ܑD"q��V�%����l6C�°��Ė��0)@�ٴa__�y�Z-����Ǒ�7o�#t�TJ&&&ddd������Ɔ���q�`���A)�����}��ߗr�,###2==ݱ���jU;vvO$222Bg�����$@7P��cccQO]�������i)�J!�x�ݐrbb�c'�gϞ��ʊ4F,�xE����ؘ��Ɔlmm��y����lmm��Ύ\�|Y._�L�w��\.���z�������N�3C�%�I�gϞE=��'�R��q�쵴�$����q���r���f<��̥R�S�����<3 aH&�255%###��0x�'+++���3�z�j�.��E[__�{�i����^�wl�{������0=�<�n��R�kooO=z����;�q-����۷��ի���z]����޽{�@�f�r��-�q�F`��^���Ǐ����t�Fh�<y"�j���R����j�s�\�>44D�V����Բ�%�I�}�6e��D"!SSS��k������<Y]]���~[���#�!�(�J%y�7dzz:�tpp w�ޕ���t��<ϓ�����Ǒ����`�R�Ա���H%�Hp�h̴�©��:�#�n�b�]722"��:��888�{����ʊrQ	@|������288�q\�����~�}��Z�&KKK�'	��qG�����~�������1s��}�p��U!��˝;w�ʕ+�f��<~�X<x '''���������͛7;�7YXX��]���/��������E%ة���D�!z&ZM��t펙��eY[[S��)��u]����;w�H__ߩc�ٯ��ݐg��bQ�|����D���}qq�*t���z`�P(p\q�8�#���QO�C����81R�TdvvV9.�N�]300 o��LLL���rtt$��ݓ'O�p�9 %�u������k�u\�y^����!o������g�^�����ppp�}�1��f���?�i����s��|1�l6�?��2�q]W�ܹCS@\�d2)ׯ_�X��>*�wޑ���f�f�\N�ܹ�l"W�����2??O9\�f�)�����rGFGG�>3tt�^O|�:5k���޽�����ի��<�7������P�ݻ'����)
���y���*�����6t���a�~�d2I�I�R2<<�4zZ����~��rQOdqqQ����𰌏��0#�T*%333r���S�2<ϓ��ey�wh�¤�i�}��\�z50S�h4�ѣG���#i4!�q���!������yʢcf||����}����H�S���ߗǏ+�e�Y���	aF�CCC2==������C����j��� 􊑑������]���R�T�ڵkd�pa���$��w<i`ppP����j��g�nH$266&���QO�'�:�>00 �L&�i�4����X뺮ܾ}�c �E2�����v�ک����� �-�N˭[����?�G��7��j���B�֭��a���I����[�8���w~��5���!�qW,���_�x<c�C��Q p�FFF���_W�Y��ݕ���tzǅ8>>���Վד�$U1�>F�m�^,;���.KKK����744DC@�2�uejjJnܸq��1��ۡ��� ���f�Ν;255��������YXX��t��gϞ.��r9������U����벂�JE=z��N��w�W���'���zǅ���Fth`�qd||\n߾������3�{�.G?�---n�(�J$�b�u]�t�R���9��K�ҩ�/إ�j�ݻw�+����͛79��dll,�!wggG�ݻ'�J%�@���>y�7�ɉ���w���Ȉsk��މ�82<<L��Y�t�u9�1&>|�MNN���@3B%�I�y�LMM�zj�Z�������� c��+׮]�����F��m:>�z��'��ަR��=\`�qdjj*�i���胃�dRc`ssSVVV��
��LNN�0#�Q�����xڍ��B �$�����o(ȕ�e�{�n���@���U9>>�x���_r�\�3B��E��*@'{�jU�y��D"!�nݢ�g�8�LNNʭ[�:n���ޖ���s| ��i�}���qj�ѐ��YY^^��g���,..nE���h?7!�
������r��]i4ʱ333�s�3K�Rr��-?�z�Ւ��9�����1 k��+���233؅��}Y]]��j�{�U����G7�G?Y���&@w]W��^������*Ǎ�����3����^{M
�©�ONN�wޑ����g �188(�����Ը]�N#L����v�V�l6��k1�8�\�|9�i����g���C���W�K��r�ڵ�O�266&7o��XҾ��%����ls ���f��^�����q�z]�߿/kkk!�q�����
NX������C��6�H�=���yr��]i�Zʱ333��@["��7nt�����,//���%� b�u]�z��\�r%�w������Sy������l6eyy�����k�Y�p�"@/�J��XnaaA�����8��2��ܹsG���כͦ<|��l��1::*�o�Vf3www��ݻTA���~�6�t:��~{�E�.�>@w���;88�'O�(�e2�z�j3Bȝ;w$�͞z�}���� �I�P��^{My[�/G�\if���������$�N�8#\4�qdbb"�iĚ���� �8�<O�ݻ�,�sGnܸ�{-���r��͎[!�������R��B� ��}�j_:�F8�V�%O�>�x�]���v+�J��]du�N��~�?��;11!!�6s]W�_�xV���
��@�i_z�m�}�sss�vB���@���:^O�R��[����eu�^*�hf���=YZZR���r255`�T*%�o���0��jɣG�duu5�����Ǖ祋<?N����������*����d2!�mpp������Wɞ���<�����8�q����\.'w�ܑ|>��z�.<�����g v(�J��k�)�W*�w��43����Rw���r��ȥK���F,Y��E�S���ܜ*Ǎ��K3������*�޽{rtt�� �.�\N�y\�V�w�y�EO�T*�����z2�d���Yd�kt���:88���E�L&#W�\���`���1�y�f�恻���c�����4moz��YH3�������$��溮���E=�ر2@�{��/�󎲴]D(mG�˗/�&��ܔǏ�� ��u]�qㆲ|��}YXX�ZtGoj6��Rw�I0���Y�fe�C��^O�<�:wzll��8��8r����Ǖ��MNN������{ccC�����{�����w��J�(u����f̺ =��K6��z8���#YXXP�K�Ӕ��T�dRn޼ٱS���277G�v � cccZm[[[���i�Z!�6y���4�͎�)u����h�S��tVh����ܻwO��}��5�����R)�u�VǦ��VK>|(;;;!� �T*��h;88����K�^if�E�ٔ�����9��nTA\,���t:��,
3����7��J%~��>�LFnݺձ�D;8�9  pv���r��m���l�utt$�����T<�=vwwehh�c ��d�P(p/�����������Z��/����Cy�(X�A�D;�j5y���r��r���f��r��c����ܻw�: tY>��=n��jr��}�J��,//6o-�J�J�issS���Cy�_��_��|�#��V�	�9+�^�=�:�jjjJ2�L3�-
��ܾ}�㾴�����T�Րg �)��ʝ;w���z�.��ߗJ���`�Z�&������K�`K9�#���������\�z5���5����s�����ښr\>�����f[���=�GGG�����j!� z[:��;w�(�6�My������flll޻��#,���Z/�\.'���#���_亮�J����3�<O�߿�5�ڵk,��]����]�+��<x�@�2 p�ɤܺuK
�B�8��dvvV���B�L���,//��tZ��'�'���O��O�o��o��za�"@���H�-..��ёr�����R��`S�Tdvv��|  b�D"�t�6���ѣG�����`�����E������u��>�)�q�Fh�+�^����V�Zg�'�I���aF���А\�~�� ,ẮܼyS���/�?����f�-//�ϋ�"��Z��}������^/�N�g?��X%s��_���߱A�u��}� �ʕ+����4e���<|��� ��UO��e~~� "�G���z���P�n������~h���?���я~4���6�t���y��lmm)�������h3��FFF;q���ˣG��f D�u]�qㆲw;H�yN@�mmm���I��\��q����}-���ԧ>%��㡾f��g2���QOg��g���ի4��˕+W:^/�����c�s 0��233��/,,�C|ߗ����1��d��}�s��^__�|�3�	�5��� }hh(�)������Í����2<<�9/��d��"g�)wG�R�����דɤ��̳��%������>�!��_��P_����_F��j5��p��fL�J�R��R��9 ��t��q��󡝛s�����Ţ$�g�W�8��ٟ�Y���������B݋dl�^,cՍ�<z�H�ͦr��Ԕ���fSvk?<<�[; X�,�����8����j5y��Y���(�2`������011!���'B}͋flLs8���eY[[S��d2r�ҥfS��9?<<�[; �@�q\___�v�T����ؐz���z�P���    IDAT �c���/��/Cݏ��233��^#t�V�σ��]�z�ʈ��������9�I$r��Me�i�����AH3�i<ϓ����1$����k"������^��y����J�R�S����J�\V�+�4��a�|^nܸ�q��Z��Ç��I  �L&��͛���y2;;+���!�����l6�	O�����կ~5������9k��g2e)��j�dnnN9�q���l6+7o���7���,m �+�N��۷���VK<x��U�Cu���� ǮY����#y��|�3Vn�0.@'{n���%�V��q###,���t:-7oޔd2y��V�%���Z�# ��2��ܺu������hȃ�V��43����H���:^�'�loo���z�;==-��k���*�t�q8�"�z]�<y�纮LOO�0#�&�Lʭ[�:�^�����  ���dffFُ�^����,۞z���Z�偁zY�����#y�O~�2::�k�W��+J$2<<�=>��pơE���n��.]�����ݽ7��t3??/�J%�Y ����/ׯ_����� ���X=z$����X���j���%ccc�^w]W��b`�fy����п�}}}�[��[���~6��}]Ч���o��o������<~���3�E999Q�y�A�|�r3�i�]���aii�so�G�J%�����O��;88���9�u���{����wL�
�T*TYX��jɗ��%���?�k�ʯ����_��<|�0��>c�#����-2;;+��)�MMM)��!~����I������F�3 �fttT.]�����+���ݟ��j��ǡw�e>���G�������D���aL���/9�)@S�\���M�L&ӱ4	�511��gggG���C� �T���Z�!777#i2�hmmm�������,Q5�����y��?�k��z�^�o|�QO�fgg��]�r�=c=fhhH&&&:^�T*2??�  ��r�
帧O����N3�)<�Std��U�8�O��Vl�1"z��7�IgKlmmi5����244`���>�z�j���jU?~� �{t������/���rxx��`������X3���r�g�W�n�7�|S>��E��gaD���/})�)@�n�szzڊ*\�t:-7n�����Z-y���4��g �A2���7o*O��<O=zX���Qeы�bH3��j7���o��o�+� }iiI��梞4lnnJ�\V�+
288`�v�#��nnnN���C� �6�lVfff���z]>|Y����|�H��d�-U�8��[j>�D��:"�ig���R�\����������L�MqqqQ���C� �V2==�w||,sssl��!kkk��ًn���-������O~���H�f�)��ַ��4���k������fLNN�ߛ����  �3::xH�����0#���� �gU*��|>�p^���_��_E��������둽�J��w��]�T*QN<�;��s􆡡��c�*��,--�8# @\LOOK�r���*��{�NGwz ��?�a��������&#п���E��д����xppP�f
�������F��C ��9�#ׯ_�T*�;??O��qpp��K&�����p^�z]~��D���B��,zdz�\���~;����V������yoH&�233��{��dvv�� �W�J��ƍ�7m����f3��!J���d�-��}.�����>fdr1� ��_���Z��^�VWW�V�)����3�t������=b  ���듫W�*�U�Uy��1�[=���,zL<y�$҄N�P��~����~'��0��y������/_��l`���������M���
qF ���jW.�i�#t��0����/|!�9|�c3nA'� �ɓ'4����ښT�U�R�$�B!�!J�R)�)����k @WLOOk=k������n3B����O"�n��|�+��~�X�_��_�t/�$@�9��|��ΞONNvy6�Z&�	,1l6�� ��q����d2������=vSut/��E�����looG:���������dC�[��|���eqF���ZQ�l���㺮\�~]�D�1< �-�JɵkהAW�ٔ��Y�</��!
�JE�E�?����/��~�T�~����t/=@��~ �r9���%{>55��� j��Ӂ7���5���qF �^U,�ҥK�q���l����ًn��~��QOA����&"F�����|����+�m���������w�^�Th� ��ĄV�������0#D��� ��3�J�E�@�Z�w�y'�i���Y�P����H�����y�qd��-���m�l6enn�}� �P9�#׮]c?:D�,z\����M�S��E$�$B����Q�F�/�3z��V�<��K�XaF�B��s�������ٕ �ޕN��ڵk�q�VK?~�~����<u(�NK.�qF8���Y�>�E�ע�D�:��̷���5����655X���ɾs @���b��m���lǊ�gϞ^�����ͦ|�{ߋz""�QD"m�Z�^�T�޽{a�Ρ\.k]�LF���B��P,ett�����y��i�3 �t���Z����u�����N`�n6��L&��e(|��z
""�E9�����zKZ�VX/�s���>11���1�J��;�<O���( �u]���	ܒ%������yi6�!�a�}_���ǐE7����)Ϙ�1�-@���l'''�� ��gJꔓ�NW�\	l������n�  �-��jm���벰������d`.��j,��Z-��7��4DD>,"?Ջ������Ç�x)�ӓ'O�3���+W�a�������rY677C�  z��ƴ�����*3��S��
<V�q�������~;�%���7�iBW>tP��emmM9�u]aF[:��˗/w��j��:  ���k[\\�赘����9
��&�---��-��Ed"�-@���>}��E�t:���j�D����E�T -�N˕+W��Z����͑<��F���,��|ߗ�|�+QOC��y��!��z����I��`�VK�����NLD���.���������d{{;� p>���Z'�T*Y__aF���R�P�ٱ���/G=��� "���������-V(�����-�Zǘ�.�\.p��hhw� ���ӒJ���VVVh|C���rxx��z"��|>�pV������hHD>��v=@�������+�͞_�t��3A�Ǒ�W��"/--��	 ��d2�U��y�,,,�H�!�\��Ae�"Ϗ\�qAW_�qY\\��K��������r\6��R������佽��n�  ��T*���r���lll�0#�i?�B4�NK&�	qF8��}�kQO��<?v-4]�]�eU�`KKKZ����٫3�l6�*��j�� �ڕ+W�Jݗ���Z��0#���}e���f�mb�O��b]Ѓ�B#Z�jU�P�uell,�!LW�\	<f��ӧtm X-�L��Ԕr\��񲽽-��u����U������[QO��߉�dX/ֵ =�HpΠ������FGG�񊙱�1)
�(;� `���!)��q����l*�\zB�����.�)�%E�	�źAS6b.��duuUk���x�g�0������d  q��k[ZZ�z,ft�ű��\���&m��������Z�Ί��666�V�)��E������������U��  �P-N��Z-y��i3BXTG���˳��Z�����?�zm�"�o�x���|�ͦ{���x)�J�e~�jU���C�  ��\.����-���!�aQ5�#�h�/|�QO�E��E��
���R�h�xR����$����F9O�<1�� ��8�\�zU��yqqQ�O찷�'�f���L&���ј���z
/�e	�Y\W�h���keeEk���({rb���˒N�;^��ޖ���g @����dddD9�Z�j���|ߗ����1d��U��enn.�i�%E�7��"�;�#}}}����Z-�f�V��l6+�����Z-�m  �lrrR�ɤr���:g�ǈ�̽���Ĕ�>���G=�����fq���y�����.�FC9�X,J6�aF���t�Mgyy��� ���H$drR]��y�<y�$�!�j�fq�w�^�SxѴ�|��/p�4%"��-o'{����[NNNN8� �S�����=��r�9ڰ���uttdZ��Ot�/�� ��v3J�\V�K��244�m��*����4� ��q�ʕ+Z%�KKK4��	����K_�R�Sxѿ�+���/4@O�R����s=i��ǝ�� zR>��JHT�U���aF�6������n�SxQBD>֭��Bt>�f:Ks��fb�G:�ܪ�y��  =mrrR�o���
�Zb�fq�Z[[3���7�����gϞ����.&���o0���R��B�  fI�R211�Ǣv|T�U9>>�x�u]��r!��|ߗ���QO�E�E�g��_X���\kkkZ�t�������T*u��l6�+*  ����1�����rtt�m;;;���e��|�+QO�e])s�� ����T�V�?D"�X���C��mjj*����Z��f ��t��<��---�0#t���^`��l6+�DW���9=z�(�)��"r��.,����L���Z]�����1�������ߓ����
qF  �Mu�l;88�صh6��'9�C�P�jմ��a����^X���L4������˗�<}��c�  x������h<���ט�_�b�Sxم��_H�ι�f:88�J���N�e`` ���T��*�����8#  �P(������ȳg�B���\.6P��hs�(ND���E�����d���U�q###)a�D"!���c�; @g�/_�zZ]]5�'��Ι��7f���2��RFD~�"�B���<O666��R�n���1I&������} � �\N������3̥
���|H3�Y��/?�я���������^9@w������-�z]9������r�dR�=׭�  ��MNNj�J���X"�K�Z�x=�H��l����z
/�%y�0�B�r���jf�]��h5�]�t)�;���#���!�  ;��i�g�V��݈�Ru�'�n���٨�𲔈|���	�a�V����� �n�tZ�Eaee%��  `���	������4�f�n�	���d�����ꇈ\X�;z�6O���L&�-�.]
�q<{���0  ��J����x�'kkk!��R�V���k�o}�[QO�e�("��kz� �u]>��-�"{n7U����= ���ǵ�蛛�Z=`.�����[oE=���rA��_)@�k�V�%;;;�q�����P3B����[[[<4  pgɢ���n� =���o�@QO�4��"��W��q��y677�����t3B7�4��y  秛E���`/����z�Q���H6�qF�qrr�\\��/��+g@ɠǌnP622�噠���Ǖ�s�� p~�TJ�y��<�-�
�HJ��q��W��4^��_~տ��z2����a�����*�Q�n�t:�|`�i  �Nu�iYt���l6K�������G=�Ӽ�>�s�XI2��֖x�����/�d2�������;;;d� � �TJ��.{���h4�e�4�6���r�S8Ϳ�W*3?w�Ny�y8�<���s  B��V֦�f����N�n�f�)���QO�ey�Ы��������<����;88��٠[���K������  g��d�T*)�5�M�d	̣��,� \���7���i^�����D"Ap�lmmi��
�;K���<�&5  \���	�q���Z�a�Z�&'''����Lo��v�S8�/�H���t��ͣ�bKs8{�8::����g @o��r200�W�׵+a�r�x��<+++QO�4#"�3���	�c��<����Ky�������� ��t��8���E��}�ժT*���q������t���eooO�h�|>�{g�����c�ժ�  p~���Z�Q'''�@f:>>�Z����3m���z+�)�&� �u]�_F�{!�s{���onn���!� �ޤ�fk#�n/U�;�.�|�{ߋz
���"r�<��t>����N�n�|>/�B���V����  ���А�R)�r�̩*�RU?���<���QO�4�<?�����4K�R	,�iK�R���p�T���� ��q]WFFF��nllty6膣�#i6��'	�E����H+�����ɠ[N�Sh�T�����ɤ��Aw�  xu�����G�����@f�}_�t�x�<���HD�|���t�q�@F���T*uy&膱�����r�,�j5� ��R��ֶA��!�,�ck�����|'�)�f@D>x����ʧ�f�da�h4���:�#�b1��"9�#��ÁchB @�FGGeggG9nccC&&&x~���Q\:��u��f������?��]}�����t��	�-"_?�p� ��"�looku����d�Lo5P*��8�j5�  \���>����Fp�z]���i�k�f�)���{o9�#�l�F���k�����Űs.�����g��T���jf9��s�GՄ��9  ��:�����8n�>�����~V���k;S�������X&�������}�� @����$�H(�����aT��I\��r`deiRD~�,��v�Αf)��R�ו���4G�YH�=��ۣ3,  r]W�����XT���qk�؏�.:>:�z
�����Y%2�Nc��6�9c���  ��n���֖V� �Eu��Yj5cO6�����)o7����8��ۧT*���j5e�  �\.'}}}�q�z]���B�.�]<�3����"2�;���Z����j"��fR��Q& �9TG��mmmuy&�h��H&��=�8�#'�Ɩ�k�C'@���ޞ��P>�go�e��7z�m  �ohhH\W�H�����?�����8��dB�T*�V��K݁Zz*��m���?���>�Uxn�  �%�Hh��9�	<0���R��D=�N.6@g��Y��K�S �y(s�/��ۥ�06����hu��
�)�0G�^���C�8�q�n�����-	g�=   £������h=��� =�Nkmq@8<ϓV��4N����$�n���]�c:���;��<��p;;;�v� ��9��u&�Yt�4�M9>>C���|�V�;t�薷���,��*��qC �\��n��`�]*�r�S��_�R�T�L�At�?'@�K�XT�}NI  ���rZU��FC�ec�B�F2�,+�Oev�a��8�?�de����ZMYb#򼴣P(�0#\�����뺕   :�����n��7	M��r9������o����F��t^���)tJ6̡� �P(Ь�"�DBY�@� ������q���]��X��l��I��]:M�v������j%8C��:ts���i��{�]TNNNL�a  �H�RZU���i?���2w���p�����������j�������!@�'�� ��}����]؇n����w�yssC>���?�4g�9Հ� �u]�5�l6��0���#�L*Wڹ� `�R��U澿�o�y�8ő��T*�S���bv����ߊh6�1*"ׂ~�X	2����֪O>��d2p��b�M���ؤ�  ��J����O9��<��B�^�^�Z����8$6rZ���ʗ�G�$0�������Ǔ���i  اT*i��=>fPe�In��#k��|���l��g�.�[Bw�� ��DB�~q� �>��������n����u]������|�{ʎ�!8��|ߗr��5� �����j���  X(�NS�Cd��r�ҥ��Y�ٔ{w�l��_�H���� �}f8::�j"�L&�a������v  �[����'''���H*�1�B�FGGO��Ǐ�<��ɉ��.vГ�$�Ay{�8�#�b1p��  �Ku�o���3��'hPU7��4G������s�U�#p2���-o�)�������ͦr�  0W.��z��o��+{��    IDAT���(�Z�&�J����Ӆ��?��͠��ӆ9T�ꔻ `��d�aU�Ne������� �"2�j�Z��6t{�n�4� �~�:�}{��AM��qN=nMD�V�|�}H�����A!�n�r���G"��J2�aFxU�l6�����D^v  ^Q�P���t||,�Z�44���c����8N�Fq	7�lާ$"ӧ] �n8��Ǐ��k�R�f��l  @���K�{�(�ccc��y&kD�{�>�S�D"!�D�
�ΤR�nU�}�E  `����q���A�8{tJ��<�S���� ��9tt2�vp]W���>4  ��,z��0���I�u�B7�i1R�4(�l6�ټ�~��3�Z-�@[>���lp
�B`�F��,�  �H��Z�/��8n��g�T*��{ �wZ���33��T�:t3h5��d24���j��6  �2�xi6��~Ad�������o����f�>�E�}��St>Pf�T*Z�(o���M�v  �G��� �:Yt�app��.K2s�f��y����z�)q7�n�Ny��ɤr�:  �300�u6���'�XB��x���������ʴ�����8��� =^T��j���  �P"��z^�}�,�%Ƞۣ��}ttL�����#�������/@O&�Z+|�.����P�nU�vn�  ėn��n��"�n�B� �DB����Wg��0����PZ��r\"����%T7f�� �/�B}�v�V����Q�l�|>/�����LMMG=���e�=���J��)�� _��V�NNN؇n�j�x� ��lV~��M���䎼��A7�n�~��~0�jռZ�J��i6   l�DB�,V��6G��*s'@7��8��ˉ���� �PGGGZ���*o�F @�鞇�s�T�}	���8�������=e���� �A7�Nw;��"p#  �؇/d��qr����ȍ����<�S~��tJ��d2��t�F @���:::2�$?A�n�jU/������=z"�0����t||����H$XP���ʡ�hp�9  = �Ji=������ѩ���gv�t34F��ϼ�/��	�̠��Ly�T���  ��2w��J�pB�u��1wΠ�2��EU��
9  �C��]�yѢ���׊z
A:g�	�͠����s;� �6�x���|ߏz
A
"2�����|���k��d�_�  �\.���^��~4D�Z�^'�2���͢�A7����82��S�??99�f��l  @�\��N���|� ������M�O�Y�^�V�VK�G�q�d2!��B��= ���6��M� :�*�u%�H�4�ՂS"�n�82���!N���gt  �2��h�Z�jHb,3��>֘ �T�N�md��@�  ^�[��s�T��Ƞ��� }�����dRǉf:x���#��(�Y ���r9���z�.����7C��n�F������?�'@G���C�:��o   ċ���r,�O��8�-�3�?@ge��%��棼  t����������6""2��!����q  z����T%��Yf0<@wD�t��Z-e�LM�̧*q'@ �w�6�ӭ�Dtt����+z���_!�n݀-�H��p��*Q�� лt�j�*��wy6x�fS�k�Au$^�&E^�	���Z}k#{n>Uٚ�y��J   ��鴸���y��3"��
����P�����:���l�t��3��R��  @7�ζ8�������G�M�P�n��P蔷  �Fq,�O��5C����+"����DO�|� �|�  @���� ��3�#"?	��,hݠ� �|�  @�z|����&q�"/舞�/M�̧ZD�F  t��xn0_���e;�<������=��J��]Y��
  t�f�iz�����kY��^�ٔ��� �l�r�F���^ ��r]W���,��T%��h���j��ϫ�XIDd�����H$x��Z'{  �t��<?���l����c�M�E��tC��b�R�T�g�W��Ѳ  �؇��y�l��}_���a2�P�Ŵ���:  �E��>�\�sG<��2��:�����ͧz��� �6�g;�ͧ
Љ���j�p��)t3�lG0��ً�{  �O�I��#�n�OD"@7�xpG��  ���C�����KJ�A��x�yt�k  �TJ�Q��<�gé��%)jÏ;�#@7�xP��7�M�S  �������,����n�K��(q7]���v  pV�e�<G�� �M�+Q(q7M��q  �t0<G��.�v0����e%'z��k� @7���a�  x�n��s��T��:��}��{�.+9�k�Z����Xt��n��| ���>���M'@'��^�E
��
�R�O�sc  /#�:�dѣ�yFg�	�M��c�{e>�
��]# @����}��f�m�ӭ\�H�e'z�?�����=�  �(q�U� ���|H���U%�n>t  pVd�� �|�gt��&�n �xH&��}E�X ��t3��~DT�#@���z� � ��ǃ���qz  �w����<�~6f�,t��$%���Ƞ�M��pC  �9�I=<O�MU�@r4z�7�#@7�n��{e6t  p^�����Fw��HB��	Ƞǃj7T  Љ�s�f�G�~�Ƞ�@7pc1�l�+:  �D���f#�n>��M.s'�n�2�f��  ��n����؃n�78�·$z�A�U�np)  ���s�fSef����8��ߣ%�����^�M��k�  ��n�F���Ƞۡ�2����	tK��ͦz�� �Nt�2�wB�n�V�ح"�&�ͬ�^�M�sC  ��A�����<<tp�Z<�A  ���ǖ9��2TĚ����'�",���=�  �t��x�0��0�mj�A7�����ltq  �E�x���|1�{D���Ń���  tB����-t�A�t  p^��y<O �7v��&q& @��P @'<��%�v0���:pQȠ ��"��?v�ɠ#t  ��F��?v0�m"�n�x��  �m��������Xi��A  �Ew <���W�:�  @'$l��x�~�j� p�n�  �t�#\��w�U~���� �z�� �NH���������	�  zM����ƾOU����Wf��  �E����t�C�  ΋��xPmi�}6����52��Ľ7� �NȠ�qc��d�M�m<�A  �E��@������d�M@=<���  t�z�h�y�l$d,a��T�nt��n��D"��   ېA��Y�����ɠ@7p�]YE4T�+�  ��V��5� �l4���o�s��p��?܈t  p^���f#@�����A7��-��؃  ΋z<���c�#t��ВA7:  8/���{���&����k��xP-�pC  ��&b(q7���!�2��ߣCt�A����L&C�	  ���s�f#�n�g�A7��-��� �y5�M�qg� �A����# �xP�?�P @'�:�f#@7���fg�)q���t  p^��y,��� ���"�n�����Ƞ ���}�=�1A�8�9�cr��1k&����-}B4t��t  �$ax�0���!��¡KV6z�TJk��Z���GW��  ��,��;Q'ވ���O� ��Ǉ�K�  ^�h4���a>2�60���!���� =>T7�t:�L  �-t3���SU8�=z�n?�}��@��V���R�`i�  ^F=�!@���g���B����}�ԆS�`�� ���A��~<�G����tʦ��H$�?(�_f#@  gE=T����Sk �5<@g���J� ��Ƞ���H�<N�$�����V���g2��f  lQ�׵��l�l�f�ܣ
��Z�A�W�
�P�?�  �e�:�fSU8��A�W@D��"|XL@��l2�Tv�  ���<�
I2�fSe��Zl�K��"?	���DO�Ww��h4ʊ�� �6�g;�u�ec8J��`��hW� ��A��� �.��H��G�n��mJ܍���K���T+ᔧ �6U��6�̧��$)j�K�	�M��� @  �Ƞ�{��J����t>,�#@�U���fC�	  0�n������wq�!�n��P�h�� �6��P~�\��}_\�� ݗ���a���y�_�S�h)Q  m��J��q��1<�G�qS�<.�H]� ��DB����9�Q�V���i�Kk  @H<�czL�4�Sŋ����W���L����q�ٚͦ��7Y  ��tI�R,�N�]���͞����1�n�F�n>��  ���C�A'!j��Ƞ�H�Ǘ �|�C  *�mqm�棃�m'B�n&��899	����C�	  0��y�Mw$��J�o�!���+��x��U����4�3��ˍ  ��t;����S�6��@�n2��ZD�F @o�}_;�B��TM�Ƞ�!�XH��F�����D�z|T����4\�e?  =�^�+O}y�̠
�=2�vH����� �M�t���籠b8�Uqt  z�Y�����l�*���="�2C:c�bt�����[��'��z�(s �w�>�Q�n>�����J�'�0�I��t�)s7���q�un�  �.�sB��S%�Ȟ���s�OD���t��Ǉ�t���/��   �薸�`>U��h4B�	T�.��⿼���1�n�3%���9j�u��1   ~<ϣ�{�p�\����g���A7��0�����rዛ.  ����XkOr&��d��=��	t;$���/�t��ǋ*�N� @���Ny���J{����n���>�[�{v&��>t  �2���,�/�L*���!e���"|xL�N��K�Ȣ�O�BN� @�!��#�<�#�f��@�⿼'@���������Q��|>O�8  z��y��B�����U����t6�)t�9����?���S5�s��q  z��ёV��l6+���{f���T(�#�XL�P�: 3�身���*���8  �C�\���Ƞ���}SODhH�s�E�M�[�N�nt  �F�/�:�ǉz
����{:�S�n �d�#���FL�;  �C��� �|��A������/�t�6�<O��z3«8>>�k��d�@ ����ֳ���f�t:���}���Ʉ���_���D��z]�i��,��(s7�N������f  �rxx�5�P(pʋhg�.g�E� �BwՔ2w;�n��  �_�R��s����c��t5GV�����$S��=^� �n}``��3�EP�$>͑Q�W"@��n�F�n�9��K���  �5�M��6�qX���*@�A�9�Yc3蔸�B7�~ttD� �ܔY-  �t������n�q�{�I|���3�EȠ�C7��y��j�f�WE�;  ����x�f���=�#�i��@?�ݗ�� �Pg)o�Q�T7fn�  ���E�=���ɤ=�EN	��0�C�����3�EPݘ���L.�  ��l6�Z�*�9�Â�%(o�G2e������EN	�)�0��4t;4�M�{�M ��988�����O�XK��D&�i�Lƞq"��"|�LA=~TY�b��L  @Xt��y�t{�t���
��VS�z��{f������ܘ ��r��5�� ;����m����ln�����EH?@�+������i��������y^��L��  pF�jU+X;�s��ʞ7�M�A6H*��z
�̝����d��2�x�}�n�  �U�\[�X4�8(�@���X�������ɠ�C��I�lMDOu�i&  ��t��K�R�g����t @7��G����i:f�)�0z��n�⺧~5 �E<��~F#@��*�N��s��Ήȩw�(��f����:�u���j�g���K�;  1ppp�{��P(H:m�>Y� ��� �"�~z��B�ȏ�3��+�BAk,Yt{���^��  �Q�?:�ϩD6G.�GE����"�V��=~T�йQ `?�q,�ۃ��v1�2� �f�:���qxx(�f���t:�Q+  X���X+X�ot{8�cr_������2�Y2��؃,:  ���������(�4C�#���+� gϠ����B!�E[��
l>�� ���Ї���<\�\.���<�� �L&�)tr,"�.v��y��
�A؇?�ή}}}&��  ��ժ���(�%�INn���vɘ����k"�2��fS+�J�g���y������PH�  E7{>88(��ty6�(����d5K>olo����E:2s���Ba��   ����i��>oU�&���}_�Y�3��|��Q,��V�U*,�*s/
&  ^R�����X9.�HhoaD�2�L�3���<��u]�;��?@'�n�D"��G�}��h�ZʪV� ����ָR�dr ����?�4%s��F�q:�{�ѐV�u����Q�O�28�� `������.�I����c�\�.�*t>l&�='�Fqv)�ˁa�BA��l�3  �Q�մ�ۓ�$������N�Y򊊇��Z� t��v�<>>���"ts  vvv��Q�n�d2�<������}_��?{w��X�݉�q�����L��խReW�Z��eIo�j�!)l�
�#�,G�c(�~�ǖ�c�أ�3#OuWK�*n��	b�w�^�H�S�	�{��.���Q�}H�*� �}�s�O���@o�0bА��n�y8���ݓ��ЭE������̏��I��w��Rl�K��e���ϟL�-G�9t�Y2�r��N�3���QmNBDDDƩ�j�>7;�N�ri2�?��R�����o�N�����jTtv$4���lg-�,�Y��i���Fͼ�G}�MR↦�
$�����/_|nt8?����3��errRӋz�ZUܑ%��R��7t"""�e�N	:Y��nWl�+�2w�M&�z�s�n������	�w?18�/y��@Sw
>���n�k��.�2w�-�Z�*ށu8��JDDdB�b�v[u������!"z,j��y��|nnnn�^�e������kՍk=t�-Ҕ��l�\��:����u�]w"""��ڽ=�9zl�f-�n��fْ$�/���\N����PW[�)A��U��Hk��t���r�="�����v��iS�f����1A��j����7�M�o���[M����:řG(�(�����:�XL��V��"�܉��LD��zO8��n�!"z,n�N�s�u��2�^�ggx��ѼGS������EELLLhZ�2w�Q+�����)"""R���ѥe�����ruu�x������ȟ��%� ��͆��GW�XT����z9�����ժ���.�KS�_2����"�2�ɤ�d2�ˋ�"z�㕸<_a6Z���E�ٳY���d��.<���鴦u����j1� �&���4�N��)g}��u��=�-��nQ�@@q&cO���,��K-A�F�<�FDDd�n��|>��NNa� �ϧ����h�G�)�˚ֽ}s<�H�?,4tpsƟ�h}�/
C��[��R<��N�DDD��d2�>G"�FcdN�PH�:���GkEK:�1�����v�	:�]t�a�>��vѧ��u�����~���p|��&��y���5��%���w{M�;&�Sd.�h6����Z��ǂ�Ţb��ǣz6����_�\֔���n6�� �өx����GK�/��t��2��w��EE��a�u�,sݢ�������	��R)M��>mMj7U��&���L��T����:�7/�S��t�a��hK�ӊo �H.�Kǈ���ƛZ��Q155�CD��X�n=w-��������N�cāzR����P(pܚu�]�r�gd8r���H?�TJ�g�X,����I��~�5L������H    IDATN�u>&z��u�t�OH���|�z���ݮ��d.jet��Ӛz��H��霫 ,o��@ �xc��nߩ���qqq�y���@(41�hޣ��9�}$h�A�2��̧�h�T*�.�"�� �ɠ����<�fQʉs!�i�ۨ�4oPc~aA�ͭ���;GV�V��%4dZt�Ri2/�]�x<�S$DDD�K�e�[ϟ[��FV?��C�d���e�t�u���Ą����f�Nw��<J��b�F�ۭzǗ����P(hj����8Z͢|>����n���L���Z�Z�͆��>b4}7Ax��lA��,���֕L&�����	��Q{�r$4,,o����s�kwv�*WI<���w��{%�܅5���iM똠[W.�S��T���ݕ�eT*�un��pX��h��ۙ�O���<bME|���rD���;������D"����j���[�,˪gѹ�NDD�������B�!GC���x�v�^�$���&���Y�'_�%�UǏ�N���=�f�	I���4$6��e�c ��(�����x<:FDDD4�����:����*���]��J:�|�ln�����M_�$�,s݄���sܚuI���A�݉����͍�u�x\��M��t��������`�����x�I�>I�(�BE�u�JE�,3�[:�V�`�F���JDD��ͦ���ݮy�����r)V ʲ�#�&$I2���p8���?�S�B�L;jxu�/b�>BDQ�TZ%�2��-���(�����DDD����FSYs<״IB��؏���T�T.��+�������䤎Q}�+ wn\p��^���	i-o�f�C���)�L*��MMMq����Z���Q133�CD4,j	:7&�)�H���N����:��?����t��K�\� *į�j�d2�hv�]���n\H��dgQ�N�Tj���.��ɉΑ��D"�i3�����v���%Ib�-�e��Ϲ����/⓯�,9*tzw7����Zum6�e)���R)LMM�P055���k�!""�#�H$�x����Իq27?������am}èFp���>_����j���/�!���є�g2&���t��d6��x����FDDdqw�=7YB@w������x�_�W���a(���}��A� �ͦj)5�orr�Cu]�VcɎũ�E��b<�@DDt�fSS����Ѧ��z�v�^gy�y�A�CPs�p�/|�F��f�<��⬭�� �L�.���t�����ڮ��5�4������q�ܚdYF(�����u�x��O\sb7��J�+Y������;�z]��s��ɳ�#@��97"�I8�N��Pc\��'�9��aŒ��z�Ο��u�]���(�����)"""�Һ{>77�����@~�_1��v�l�kRn�%6����_��W�N��V���oC��� L�t:=�hh�2����a$��"""�j����Q�˅��)"�a��u�!�C��'���G���'�9i�О�f9>��$I�.:�\]]iZ�����s���l���03�1/$� R��b&�#���#T�p�n�5�1&s�d2��FC��j3""�qT(P.�U�y�^LNN���Ąb��f��v��cD�� Vm��C��Q�Z��X�����e�A�����"A�)"""�e��ך�.//�}t��ݺ�>��!hq��v��tI���ݤ��2�B����#�T*�T*���xxn�����鴦YבHDSe"����P�9ʲ̼��B�7WL�A	���T*��qGc�8LMM)����d�d22����x��f��vu�����|��.���:A����CD4ljG��:$I�)����H�l��Hc�		��<b��R󚝝UMЁww���[_�^G&�A4�{�n�cvv:GFDDd.777�*gff4��%�cs8�
�ÈF�X[[Ó'O�g�W �Z(x���V��L*�*�y�V�,��DB�����\.���K��D*��h�n�k��C���z������v�h4t���bii���xP�8�t�]�;���fc��1�n�K�l6K���h�]^^j*�]XX�B�h�`PuaO�Ze�k[]]5:-t�`�>6���N�R<w3"R������lvCDD�T*i1��z��t���ME��v�2��r��R�i��V�1�3)�׫:RxWړ��t���M�e���+��""7�$i�������g�7N42�x<ntZ4 |��o�	:�����uZ�c�5��e�Ł�=���u�����X�tZ�9�h4�J��V���ss���0:-~���o�	:�'���b1M��J�o������ʖ��yM�"""�S���#�"{������;�$I���:FDw!��x<�xp�8�	�X�K�8�V�������EQ�\]ADDde�v������x�z�LMM)^�T*lgb���V9j������N��;P&��Y\:�f?��L&����(B����T*!�ϫ��z�V9�J�9������V�L�>���.��٬��6��ن�@DDd(I�T��w��+++V٭#���,r�$��1��P�:��e�R2��⢦N�T�?�R�T��f��q�݈�㸺��92""��J$��G{b����^�����8�={��711aP4��=�G)?J��j��j�xvǤb��n�j�r��J��߯Sd4lWWW�B��������!���
��z��d2����tZe��4�������.?�����}������c}��ճ���a}kz A47��F���tw�A���~Q�`��ˊ��d=j���r���L�����!he���"�6??��M(�͢�n��%�͢T*���t����h8�鴦Ϥ�pXS���áX
-�2��������1:-� �������z��;R&�t:133��N�$�\A���QyD���,��ji�"��UJh������U�UN,2�o|�F���O���e3��涴��i]2��͖�j�p}}=�(�X]]�1"""��uvv�����2oJ�A6���q\�����gtZ=Zy;0�������չ���dNK�w��L&���
��ş��,)��(�Ꙙ��{��D"p8�7�M�4�H$�`0htZY'A�$��*LNk�қ��!GBF8;;S������]""��V����K�u�]Z�Ñ�=�����G��͆����~8쇠��bp�\����2�ժ������\Y����ބMj��:�G���,���_�5�����z��;z���'��!�l6���Db�ѐ��4�������NDD��N�5��G"������i���f~;z���	��g�
���0� ��������,�ͦ��Ժ�/--��v���4�MM�����a#��r)��$�"������]X/AE�jgƎ(�XXXP]'�2w�GT��������6�kkk:FDDD��,�899�Ե}uuU��Y���y�R�)��e���atw���=A,wd,-..�fS:�R)ŝV��B��|>?�����쬎i�H$4��b1Ml�z�v;"����,�9�D�Qş�ɔ �|�o�K����c���c��v#����$	�TJ������h�Z����������j��iڌ�������"C�b1�ͦj����˿��F�p�x�'�.	� lgZߴ�˃FT�������� `}}�(�� �$���T��W��KK� Y��fC4U\��sk�P�v �������J�����~�����v�LF����JE�׀��������h�����h4T�-,,����!�*6<���h��:FD�����.��0��n	���fff�z8����sD��J$�T*�OMM�ީ&""�L&�\.��.
���Aud���{d�o��F�pu ;�o�k����/�hj�R��������(6\^^��5""2D����Ņ�:���)$#.��t��l69&�"�����]|
`(O,]t��[��٠Zf��u��m����.�"���!��QѸ�$	o޼Q��;w������U��E�"��������5:��Jy;�s�������9=��ajj
�`Pu]�V�.��+��]�}>ϣ��...P��U����!
�%+V�Z-M=
�x��+�btw�����������I�����iw�G��Օ�y���i�G'""]�r9M�j�� 7�� w�G� �ַ�etw��ٰ���	����-������iM�N��*_�F�,�x���b����ex<�""�qS���^�8�Nlll�ֈ���P���j�4UZ��677�r���.~`h��gʑH���z?,֦݃*�E}�NGq>�(�����|t""
I����[M��766�p8t�����{�����[��[F�pWC;���k�?�������Tו�e���r�������n��1}DDDwqzz��,�����(�=�Aņb�v�ZMǈ�\.�����F/A��9�a-@�E�/���Ql�FU�h݅�{OO4E<�!"2Ϟ���>��j�QZxW�>4�$�.���Mw��5�J%���3�]���EMS ���ԔJ%���׫yS��-*�I��uȲl���� �	fX�6�u�[� h>�~qq1�h�z�g;�N���k�ADD&�j�prrY����vlmm�	�P����uX��r��퀁	��'O0==m������h:�U.���8&��&NNN^�������%""�I�p||<�fp� V� M�411�X���sk����gt����~ �>=�����]t�\.���j�u��}���j�����cUcDm��P(�	=� ��_�U�ø��O�� �no}��߶ZS��5==�P(���R� ����A2�T�yONNbvvVǈ��������p�X̊�tO�H�s�G��ʊ�����?�MЧ�����mdt����]^^����qvv�r�<����&''u�����*��kj
9�s̨݌���?0:����z<��D����i�F�U��j5Y�qrr�f�9p���b�U""�Z����S�u��}N����$�n����fSq������/��/�}�+=��W�O>��������i����c���(vv��l��NDD�Z-C�$�u���v�]���h� p�|�|�߰�1�����@�'�N��v��0H�p8���)�u�F�tZ���,�NOOޘq:���؀(�:GFDDf��vq||��y�f�assSq'�FO4U��_�����|,8�x׽�����`�n1�����z]^^��	��R*�;��|>lllX�)�,�x�����^+++��>fl6w�G���""���a܇.���$�$qf����~��ͩ�k�ZH$:DDf��d�P��׈���F��RIu��⢦
>-�x�c��J�>��hs8@���It�w��fmmMS����Z����$	d�فףѨ��<DD4�����+zb�Gv�!�өxSF�$�E#��r�\x����a���C��4	z�\F��KY?=�ۍ��%�u�$���J���l����8���1==�cDDDd�L777����0VVVt���fvvV�S?s���׿n�c��R�3M�.˲�'2���U8�N�u�TJ��2=�����W���011�cDDDd�B����s�u�@�}KƔ��U<���vQ.�u����C�C�/�Ο&J���[�(�X[[S]'˲b�0]�μ�f�
�����##""#T*�����b�z������1�v�X,���,,,X�9���|@S��5�M�Z����~��\.�
�1��tp||<���f���|>�Α������Y�n���ۜu>������v��j��cD�~�7���� Rz>��t���V������\��9��V����#t:���EQ���g���F����C�3�N�O�<�t��F� ���B��'-��r��?6:�����~@�%�Ri��x2�X,�h4���R� ����Q�������g����p�\:GFDD��n�o�������1�F��x^��묶��o~�V�%�]�e�L����-M�x�9���:޼y3����rakkKq�)YG�������UQ���x�^�"#�E�x|�uY����u��������}�|����.A�|>������X\\T]�j�8vm�U*�}�v`���xx���ht:l���E�������Y���r��*[��ٱ�������AM��w:T*�à;Z[[�tf���F�͚F[�TR�I�z���ކ(�:GFDD�������H��f�a{{�`P��Ȍ�n��qII��l؂dY����C�^��4A�u�&kq8��I����3""3+��x����j�χ'O�p'���bz�y�VS\g�ٰ���䜰���xT2��s���b1����C�K#Դ	z�^G.ώ�V377��6�ϳc?�T*)����|����N:�EH��7oި���%��pX��Ȭ&&&Ǫ�Z-�U�����F��� ����M�����!�	����-Mk����k�P(�t���$���z;��rYq�s��l�c��Κ�N'��o�C����	���5ͦ�a�E"�.�=�z�DB����Ԓ�@ �3�DD&�K��z�l6lnn29' �J����U�U4�X�w���l�N5��s�����$I��٥�a�=lmmi:;|yy�^�.IWj���y&��Ȅzɹ�����-LLL�����������$q�ܢA�o��o�C� �;���	: �99gSr�\lGw�����v�^��|�FDd"�v�����m�B!�"#����W�a-
�,jgg>���0���2��M���\%�F�A������8���)��uwWJҟ<y�ásdDD�E�v[�(5Q���vk�[�pX�3b����e��e��lt���O�`�Ȑz�@� `ggGqlF���	�ҭr����#t:��׽^/vwwϭ��Z-�&������]�i������㖭kvv���F��]� �H�^(���d���!baaAu]����%��P��pxx�v����������^�Α��z�����2N��������Y8�΁�K�Z-ê��������S #�D� G'F�@�����ۭ�.�H�V��YE��P�������u���h<U�U�&P�{{{�x<:EFV��z1555�z��E�T�1"zL�`_��W��-o,��ߤ�(�kEv�]�ltY�qr�1�eje��(b{{�g����\.���p���χ���]ROjU��|�G-���{��c� ߜ���̌�Ӟr��T*�CDd%�N���ƈ����-D"�##"�|��Ǫ�S(���y�{b��bg�z��JJs:���w�kt��+���T�~q�@M�	���Ύ��Xggg<{D�������f�acc�x\�Ȉ�F[*����ujj
���EQ���*�N����$Ilgq��뿮86�"�=,��K����F�A��v���������ԝ�������fqqKKK:FED4����pqqY�����`uuU��?����7n
����d~�(�?���a<�ϟK�����m�Od^���ʐ��<�Yv����������`ccc��B�$�}�V�(�n����
�����S_����}b��&g�[�׿��Q�9Q�o��`���t�����0�z�ѵ������6���Vr�D�����X��NG�HQ��f���&���u����n�c~~~�uY��!cq� ��h5t���gl-���ћSvx�0�χ��5�u�v�����,+�����h��`0���]Mc�����n����ꎦ�����.��N��i)m�f�����"ƃu�ݿ4:�K&��Fg�F�A����i,V&�Q��O�Z�b`�W�ۍ��=�a#"RQ.����k4�u^�{{{���B�&&&^o�Z(��:FD��'�'F��`�V?������q�X2A���7�KȼA��ޞ�3�'''lB���6���P*��^��J�� -    IDAT2ꏈhe2���F"����yS"Q���8�,���>FezΏ~�#�ٟ�Y���l�^��pq�0:z�@ ���U�u�Vggg:DDV��vq||�T*��� X]]��Α��,˸����ٙ�����,p�&���p8��J%�Ե8Y����F��(���������ݓ^���\�]C-luu�t�bQq]*�B(���N��U]^^�V�aqq�����Yx�^�y��ވh�u:����>��lXYYai211�؛��j�~�#�����+��xL�Q�\�U"����C�{O�>ŧ�~�ZVwzz�`0�xG� r��VWW��aNLL`ww������DHDd�z��7oޠ�l*�s:�����ys��n�����k��ɲ��������O��ј�؎�k�^��,���|>lll��k��899�!"�Z���;��n���"����
�T��`0��O�29'͖��Ǜ�����W�:j��j3I�?S젯���m���5%ߍF�(Y���"R��jÐ\.�L&�h4�Sdde�Y�}�3�(bcc������2 B""�Ȳ���k��ܨ����X\\�1B�,�*NLi4����	�&S$���?99�����s'��A��g��7�7��ONNMU�B�%�2���Q�T�K���G0���1���H��y�5�|�;q�\���x]�$����z���Cf�w XYY�|`t�@.�[[[���.޼y�CD4Jr�����d�A��������pU�U�~�Z59�x<���crNw6�xO>����Ы¡�� ~�w������#���+�H&�:DD���h��� �|��u�Ӊ��LOO��p$�I����F�x��)�^�N�Ѩ����{T��V��Z��K��D�V3:��72	������������n��ggg|��;�v�899���e�c1� `yy���Eр���Wm6赮�7Bm}}����μ^/fgg^�v�����:x�\#�J�����F�@���p��ӧ��i$I���1$I�)2%�TJ�����$�>}ʒw"��^I{�PP\�+ig��G����l6��i#�^��ɟNF*A����W��U�àG�D������V����|��H��jx������.�;;;����92"��I�R8<<T�655Œvz����\��׋�"Gq��=��H%� ��	2"666011������Sto�$������}�����yloosr �V�����...w,{�%���X�N���	�Z-�E#�a��j<V���{e^YY���ύ�� x��)�v�i�o߾Um�C�$�����`�P(���.B��Α)+����<{��]��A�N'^�$	�LFǈhظ{���K���~��xWxDx�^���t:8>>Vl�C��������s��tb{{+++|�!"�I������n\׫���Q,I&R�k���y�����tt����Z�r��Է&������w��M����fff�N�U�ޕJ%$	�n�DjdYF2�D�R���R�בX,�`0���c��!"CT*�����5�z�X__�Ysz�x\�yj�Ze)􈹺�2:��3�]�$d��a>�@�R	���<�>"vvvP*�T�G^\\���#���j����}�����n7vww�H$T�=Y��J�V�|Q,���2+~�Q�����n��hĔ�e՛���F���n�9�E|���\jY�UK����$	WWW8>>���@���bww��SD4t�z����7�n7vvv��������������s�Y=Z�{n��~���h����Σ�Z-�gO��T*�իWH&�}��|>���aaa�U;D��zGo���Uˇc��={�J2z4� `eeE��y>���Ȉ)�J��d��N��|>ot���8���UוJ%���G��M?<<�;׵�������g@�D4���:^�~���K��i�5�aQ;w^�T؏e�Ȳ����W�l6���Fֳ���@ ��������U*���#�J��ޛ<��t"zI�pyy�ׯ_+vP���9C(R<w�j��6�
�;�h��n�kX�:Q�|Eu>z�<:��c�}pTn��D��J�_�F2�T<��;^����]sztN�KKK����h�$	�D��0��X���r9��1^�{{{����6ϣ���j5,=u��x��	666�p8������n���}��􈢈��e����r���GS&�A��5:��6	�,��EA���X^^V]W.�q~~>��h,�F�|�r`�_$��g���t����"���իW��W��0>���������͟R��y�#���<�G��t3)
��p�\F�B�hss�RIu�f"����C4�)27�v'''��󘛛{��n�cee���8;;�"�����JEq������2&&&t���U4U���h4P(t���rssêS���t:mt��A�W��x<յo߾e�Q�B��ׯ_���o�X0�ӧO�����G��FW���������s�͆��y<{���9���������N�LFǈH/l�gc��s�hr8��W��� G�$��$IH&�x�����h4��|�+��q�h��ݽx��TJq��W�>??�&p4t�����NȲ�L&��H#�����蟌ݫ}:�f��
���U]�l6q||�� ������o�'Q������=��D4��2^�~���S��Z^�;;;�����<�E�)�RC�\.��8#�Z�r�D�.Ao4(��F�AC0;;�8��X,���B����)��x�����>��������q��l6���[*�4w:�X]]�ӧO9��t5??�x��T*1�Q�,�����0��� d*�B `������r���4���>����:EF�n��P(`zz�����aLLL �L����k�,���"�H �N+��l6���`nn�(�!ѻI#SSS�7�E#"=��eű����L�;���<"��ѡ�#|�~��)�R ��7o��x��zu������D"�l6�����^�A�����(.//UϨ��H��t:����m� `jj
���p:�:FH��������뽦p|M�$�����0��O�>��8�͆��UvQQ�J?��Uw �N'�������v�����^o�Z����\R"�e�BWWWh6��kC����x���t:���9�3P��)�뎮ލD�N��o��oM�d�x���Ǎ��$�������U������C.���avv�@���z����K��Dd�r������@ ���Ł��DzE����cj���󙬫��`����	��,//��v������U�E"lnn���`0���ف�j�J(�J:GFD��J%\__�6����X\\d�72���5�B�����<�*����s��3%�c_�}ss���%6�QKKK�V��]�s�.//1??�SdD��J%�J%��ͽ����~<y��r���(
EJ4�*�
���U��ߏ�����X��6??���W*&�#�^�397��O�{c�xG{tmoo�Z���_^^��v#���`�r����@ p;���:�~�&�@ ���L��T&''��^o4���:FDz�e��Mn�K��n�cee��MFX��Ə�c�D�͆���Y�DF������|}���e\^^���hH��"nnnP�T��J"#��~lll�m��H&��#����<.//��t�T����LNN*΀$��j���V�����p`oo.�K�Ȉ�������X�S�Vq}}�frD�@�e��y��ܨ6�
�Ê����r����5pz�$I�c����.���y�&�&$VVV8nk��E��'?A��U\�v�����áSdDw��x0==�p8�w7��l����T�o�Dw$I�mb�h4��h�x���ȴ�v;���n<Ȳ�T*�:������l��0L�	�I��~6	�d����:V"�ɓ'�F��r����D��i�Z���ڍ)�q��t�N��N�g?���X,�x<��dj�(bccC�ǩ��V����C�U�	��-,,<�I����/_�T]�����.�dz�(�6��0Ȳ�l6�D"�Z�f@�D��h4�N���d+N\.������
�	ǩQ�۷oU{1�33%�|w�9�d����5q����j899Q\���qzz����"#��n��T*�T*�P(�X,�����R�h4���D��\.#�L����|���A4�[������X,29�R�ɹ�0A�9�V�\�������&����d2	�˅��Y�"#z�b��b��׋h4�H$򥛎�m�z�T
�L���hlt:d�Y��i�3��("�bzz����r��b��j��9�cB�$vm�&�}d�Y�A�+{{{h�Z�3����p8��,�V����WWW�Ø����㹽��x������E��y�R)~`��U�ՐN������=���X�N����^o6���1F��${�XϠ��z���ht��N���>�L���f�a{{{�x+"+����F�����{��Z�"�J!����,���"�˩6���l������4�~��=�`0�����G1Z��{��F����#�ð3�Ag��`vv��ؘh�Z���T���l6<y�sn��DQD(���d��$I(
H��<�N�"�2��*�٬�n������4&''�NA ��χ����}�:�wSǈ,�x��;�k��"�v;VWW�0nL��u|��g�3o�wϋ���I���v�199���ɾ%��FCә]"#5�Md�Yd2�iN��h�Xn�[������`ccc�&��'�������0,�	����aLOO�Z���>C��R\�t:����˥SdD�����D"��}w��*2�ˑ)t:�Ed�Y�cJ�("� �`bb���i�8�NlooL�%IB2�T�qE��������G�	������%�e#�b?��OT�2��n��찙 �$�͆@ �p8<�z�XD&�A>���F��ۤ�T*A�����l�B�D"���d5�$�Á��́�,#�L�n<�h9??g��;b�n1n����F�A:��r����;�;�^����<�H#MELLL`bb�@�D�w^=�͢P(��==�n��b��|>�R�4�9f��011�XB4*�v;677n"ɲ�t:�zt�FK�VÛ7o��r��[���4���a��R�~���ܝ�	x��	wgh,���v7s�w��A��.
���"�ŢbR��)�D"L�i,�l6���+N�d2��j:FEF�e<�pL�-�f�aee���PHG���x��j�>11���M&�4Vl6�� �� B��{���,�X,�P(�P(���j6��ϙJ�2���tbbb�p�P���4Vl6���'�d�Y��44z��$R���aX�����$�=�$!�Hp6������,�x��b�^(pxx�$��J���7���v#
!
���C���x�]���Q(����e�z�v�|�n� �z��B��uIcK���*��r9&�c��l29�A��x<�P(dt�����z�Ju]$���;�س����`��½�ۥR	�B���H��D�\F�XD�\x��t����W�A4nA�������5�\�JEǨ�dY���1�< w�-,�L���eA�iaa�$a_q].����1��י��X�t:��r��r ����������ׁw��{g�K�Ϯ��N��r��r��R�4�(���%�� �^�Α�� XYYQL���<��1��d���f�wԛ%977gt(����% PMҳ�, 0I'��z��z��d2	�����χ`0���ۍ������]�R�ę��n�Q�VQ�TP.�Q���gE~��P�@ >��G��XZZ�=.�O�P@�\�1"2�v�}��J��	�=�vxn�,--������Hq]6��(�XYYa�N�G�V��y�/&�>����X�v}�\F�RA�R�N��4�ۄ\�g�r�n+(�� <_�4X^^F$x��׃����9{��&���L&��z9�e���B�$���F���z�Edi?������d�����������w:�ۄ�R��Z�r�]�N�j�K�GE>��6!���<CNtKKK��y�ʈ�S.��(����:���4fff�����Qqxx�����s'��nzM����s8�z��|>ߗJ>[��m��+����F�?Z�j���&��:j�Z���v�����J���yD���tۧ��R����H/�N���F�AC��
���9?+++ �)I�e�����J� �v�����z<��s��x�������&��Z�F�Z���_�n��h4P���h4n����x�3���������8�#Au�e��M�e\\\��}D1A��������͘��(�K�ӐekkkL҉�;�Q/qw�\�� \.DQD���RB�l6�l6�h4F��|��E��@��z���7+DQ���B(����v����D,//#\����n��z��hb��@�v�T���clyy6��_�V\��d I��`P��+�w:���n7����?˲|����m4�M�Z��6��vY�o���������/�w��~LNN��r��t��r1	'2Po��R�v&���tpqqat4DL�A�P�m�C�iqq6��^�R,7��r8::���:�.��n�oG��#l6�v;\.�v;�^/� �v�m��,ːe�$����n�����������,��v�_�>_��v�}�}%I���^\v���z ��p��p�n���p�� �I�l6��� 
\���k:�z���ML�I�ԝ]�����<A�˗/5%�L҉L�Ir�ټ��J�Y�!����� �e�_\#I����ݍ����Qo����h��lX[[Sߛ�f�T����y�f0A$�N777���3:2���l6^�x�xw3����� [[[��M4B�����m"R#�"���Vaʲ�l6�QZ�V��D"at�~zxD�r�5	�x~��j5E�XīW��M���h�����u��<�N39'Ȳ���s���	&����	!�࣏>Rm�T�T���K�5�"""��q:����8�W�$�R)4�##3�d2���F�A:a���$Ib�	 B��?�ۭ��^���˗|&""n����p�\}�w�]�R�;�����j�pssct�#&�CP�VQ,��L��������z����&^�|�26""���z���	����z��A2�dexW�~zzjt�3&�C�W��x<x���bwV��觗/_r�)�
��؀�޿Gs��F2��QI��J���}HX�N_�r���G)�7ޕ��~��BA�Ȉ��h�&&&���6��l��D2���HT�בJ����}���:2���a�I8|��G���V\'I�L&u������%�beee���Z��T*��tK�$���1&�C�ٕ�E�(�>���:Y�qrr���s�"#""���Ǳ��A�^�T*�f��eY��ȬdY���%�:�1&�C&�2�K�� ��������7���k�y�o�DDD"������)���r|��/)�l6=映��ns<�gii	{{{K�z��4���y�����l6����D�^�e�L�I���j�����0�`L�uR.��BL�Ň~8��kO�X�˗/9�����677�^�$	�T���=�,��쌽�	��8z���D"x��9�n��Z���/_�^��i��x�������z��E2���,�����F��0����H�$\__��'��?V��l6�����y�"#"""5�`���p8}�7�M��ܠ�n�YA�Z��'��]g�F�t��0Ȅz�ҕ� ������	�b1����q���^2�O����ٙ�a��0A7@>�G�Z5:2!Q���3���)��e���x��-+2��� 0???pM�TB&��{5�%�2���y󆾄	�dY���5��@������ލ�I�R��NDD�3Q���������eYF6�E�P�92��L&�J�btd2L���vq}}mtdb333��_�E�\.�u�b��9����rakk�@���^38VK��!�    IDAT�F����t�j5�G'E���~�i4x��J��N���@ ���큓WZ�����n���o��t�e�Y���"�ۍ�}�k���U\��t���kVfA4UlW�V�L&y�����x"����n�"Q���S����f�k�k6r||I�t����h4�l6,//cqq� �]S(��f��Te2 EL�M������/�j~~~�!�N��L&�/^��l���q:����D$�{]�$�R)1#M��*ϝ�*&�&�h4�J���, ���O>A0T\W������C�=��~loo������j�pss�&��	睓VL�M$�ϣ\.Y�������177����҉���.�bccv����Z���椙,�8==�sҤ��&�H��r��0�����=��~<s�;�^�ױ���x����h������E����eYF�P��
�I*�B�V3:�~R7I�puu�_����2�?�ǣ�.�N���?�Qn�[[[��N��T*���\.�+�	tj6�H$F�A
���'� �*����x���(���� �(�7��븹�a�U��V��s�tgL�M�\.#��Y�����~����c`�wUo߾ś7oX�ADDc�f�aqq������E��i�gҝ�>oqJ�Ϡ�X:������3:����%��?����t:�j����́;DDD���vceee�1I���dإ��L�e\\\��n
Yw�ML�e\__��j
YLo۠st=�Ql�� "�q����=09o4H$L��^2���ҽ1A7�n�˦qt/.�}����;�w�]�䝈�F��f������&�,�X,"�Jq$�K�\��͍�a��1A��f��_t�A�����ϟ���*�e�w""e�[[[��b}�����E�#�Q��p���[D�Tb2�[��{<W\����BDD4Jb��bI{�Vc�vz6�����BR��ժ�a�E��v<{�O�>�(��I����S�~��������v;���0??�w,���r�d2<�E�&�2�����t�����/?=���,~�~	���">��s
�"#""z<�@ O�<A(�{��j!�H�R����t:�r�lt4"��[L�����%��҃x<|��GXYYQ���n�qpp���s>爈�l6�������uY�Q*�pss�N�c@�4JJ��ɤ�a�a�nA�fWWWF�Ag�ٰ����}�k��|�����x�G,���Լ^/���155��z����14����&�U�����y|\U�?�ϝ=�d�dO
݀���Zm����XE�VA@6iYd/(� ����RE�M�#�}�B��k�ɞ�2[f�{~��̝4)ɬ���Ws�=3�R�7�{�9�3����x�A) T@�`��.����0��,�BDD	E�$�����#���`P��t:����Bp4#� ��Ѭ��; :t�����t]KLt0j�.Daa!��x��F��v;�͛�.Q�v�aQ�����qd��Bۃ�`�C���$����i�4c
�r�JTVVN���t���===|rLDDqSTT�#�<2jr�r������fL�b;gb�la��zzz���F���>K�,�^���O�e��f�ٳ�����(��z=.\���j�T����`����>�f\?+�Ӭb���� :;;9͆fTII	�=�؃����v���q4���f�$I(..�QG�Ѩ�'4j�r�b����X,�x�A)�	z�������b�D3*4���/~1j��?���!""�Y����#�8������
�5���v�����0(0AO!n���0Ҭ(**�q�7�J��7���fL�B�dk͝N'����9%�<�~?�����	VqO1V��EEE��RLh����b�ڵN�S�_�һ�j�ܹs�NA$"":���,̙3'�,�@ ���a&�4k�� ZZZ���b�#�)hppV�5�aP����Ê+0w�\�)�!.��v�BGGGӉ�hZ�j5�����k.���fCoo/�s�5�,���~�?ޡP�z����V�EVVV�C��V��`�TTT`���R�'�@oo/���PUU���H��(���梪�
:�N�������&�U���X[�bM���aU��R�P]]=iq/�����?������q�a�M�}�'�N���j���(���Z��qd��z{{188�0(Ft:�nǎ	�ԏ#�)L�etuuaΜ9�j���RXII	
�����u7����l6������|�)�DD�B[����E��0::���.��Y'�����s�����^���j���x�Bi�n�c��ݰ�l��38��Ñ���Ȉ�(�dgg���*�l?�χ��a�|�GF��n����#�aP�%�:�4a00gΜI��"�)Btvv�����kM&Ӥk��(��t:TTT ??_�,˰�lp81��ҙ��BKKK�à8H��S�ӄ��Aww7*++�
�I�P]]���2���L:��b�`hh��މ�ҀJ���d:�tv���m�(�|>�:����4�������x�Ai��tb߾}]�e0P]]����EFDD�������ʨ�B�^/FFF8��b.`���|(��8�Nq322�Z����x�Bi�h4�_�"�w�^��n�~����GNN;�0dff�8R""�i������N	)�����9%&�ihpp*����s���(**Bkk+��ڢV���hhh@ii)*++Y���(	i4����d2)�B�יG[E4�dYFkk�A����4500 �Z�
�s*�
���Gee%ZZZ��ݭxc&�@oo/,���QZZ���DDI@�$�L&���B�Q���:s�7!�����x�
�8\���$IBEE�Fc�C�4�t:��܌���I��t:TUUE�!"�����Gyyy�u��###���B�l6�n��;J���	z��$	UUU\�Kq7<<��{�tK�ш���k��(����PYY���,��~�V�5j�X������H�à���Z�FUUC�C!B?���wЛ���\̙3������`0���,�~��`6�N�3Ƒ)����b�w�`��S�Q�՘3gt:]�C!B0��lF{{�����9VVV�KDC:�eee(,,T<�p8X ���bA___�à���F���9s��j�
��$꭭�Q��T*1Q'"�e�%%%0�L��;�p8���Qw� �5!�������P(A1A�����P]]��*Q<��~ttt���㠉zii)����&"�AL�)�Y�Vtvv�;J`L�)�1I�D��������<��<j�%%%�����DD��Z�FQQJKK��B����f�q�4JH6�f�9�aP�c�N	O�ף����%$�ǃ�����L:R��jQVV�=ԉ��I�V�d2���$jb�t:a�ۙ�S²��0�ͬ�@�����`@UU�tJX^�7<�}�D]�Ѡ��eee�<MB�R�d2qĜ����@{{{�à$���FFF*++��PB��|0��]����5�DD�i4�L&�L&��#G�)�8�N����;J"L�)�ddd����S�)�M5QW�T(..Fyy9��QZ%���Ŝ�N)attmmm��N�����tJ&~�f�f�y�}�U*JJJPVV�D��ҊN�Cqq1����˲����ɪ�4�n7ZZZ��Ӵ1A��������
&�4dYF__Z[[1::��$I���Gyy9�Fc#$"������� ??�$E�p8p:�Lr(���n����&蔴���PYY��K�(Q	!`�X�����:i���l���#???F��>�ш�����*���|p8�>�$JT����|�D��	:%5&��FFF��с���I�gff���EEE��QR�$	yyy())Aff�b��������f���L`�NI/33�����NI��t�������>���())��0Q�	�a^TT�X_C�e�\.8��	q?JtH8��f
tJ	,G� ���p��Q��T*���,�HQ<���pb���9��t���Vk����R��`@UUG)�	!0<<���X,�I�fgg���,j�%"�X���Fqqq���^��n�����Ӊ��v~�i�$R���w ��<:;;��Sғ$	���(,,����l�:���p��p@�ף��4���DD�E�V���&�Iq������N)��t���-�a���ӌ�H:��@ ���>��f8���T*U�S�,"��������"(Nc����4vJI������RP"��3A����QUU��3(���vtvv��\FFL&����o��f�Z�F~~>L&222"�!�v��t:Y��R��n��l�v�L�)e�t:TWW31���Qu"���x e������P(�1A����jQUU��&�(��l6tww���o�5����0�L(,,�"��V�Eaa!


`0"·�Hs:���|q��(vB\{zz�
�8&��4�������
Ѭ�e�������b�:�%IrrrPTT���BnQHD \���PPP�����!<FGG�r�8ŗ���� �����&��j5*++���*�ߏ��~tvv�n�G�V�QPP���"N�'JS���(((@AA��Ұ�����Ik_�!z{{144�P(M0A���R�PQQ����x�Bs�===��뛴pSFFFxT]iJ+������<*�2�o���Ugg'�Vk�à4��Ҋ$I(//Gvvv�C!�!�V+���������ohD�d2q�Q��j����G^^�Fc�yY��v�1::�*�ք��蘴+�l`�Ni����Sy)�M�{{{�y�$	F�1\,��划�F�ANN
P��r�������,�hoo���h�C�4���Vqq1


�QB�e�@ P�*.WXX���|h��GJDS��h������<���D���{<{#�L0Dkk+g�P�$R��ͪ)�a2��
QܩT*������d��z������6��$!33���(**�u�8��t���Cnn.�FcD�`0��ä�(�@ ���nH���S\��塴�4�a%$!���7�t�К���|c$�������pR>Q�Л�嚴�Q���|hii�:��(Vi�	:�MVV***�4�A8�b��j�F�3�BT�����E4CT*�F#rss���Q�Q���������DS�r����Y��
t������J��_�(R0���,���S�T���F~~>���V����pR�V�ǝ��z�ᤜI�Ԅf���f.�����h�V���*&D�$���n'�v�=��Nfff�xUvvv�:Y�t�9!''����B���n���e��������w(D�0A'�@�V�����(i�AX�Vahhv�]�_ht=��633�	;�%�^���ldgg+��x<��Gɉ�}}}�w(D)A�bJ�`f�eee�[�����j��� ��za�Z1888n:�,������*QO\_K�*�Z-�Fc���-C��C���`0N��!�fs��D�L�)a!��Ӄ`0����x�C���z}x7 p:��Z����p8a������0��!B����ٜ�BI�`0�h4��&.�
�z�ᤜ���f^0D{{;\.W�C!J
L�)������󡸸��n�fP(I������������p@��k�X �u���FVV+�SB
%������)롤�	9�����hii��D������� ��˙�͒�#�~�V�5<��f���������x��T����F�1b�0�l�j����DVV������9n�,��bn>�^��kȉb��v������E�(�TTT��(N<�v;�V+�V+�v��\�NN�B��e���R����9�kb�u����|�#�#�͆��Nn�FI�E∦��񠣣���7cD4�����t:����p8��(eh�]�$ddd�G6CN�rL4�F�AFF233��������l*Y�����p8���ß="�?!����P���(��p�����x�C��T*rrr"v[p��I���(
i����z.eIC�$A�Ӆ�ПcgL��~���p2�u�D�I�etuu�w!�C����,����FQQ����M��g��u�\��������Fځ�Dml��i��/��74#4"n0�R� �@0���?�	�>��X��������P��tJ*�����|(--�;Q�S�T�"rcML�C#�.�V�5��I��^?.����0��t�$��I�N��^������ ���F�}>FGG��D���^/Z[[9��h�0A��]���W����C��8��{<�p���x<���,��0���P�V�e?�$I�V������}�A�A��6�-|��p���t:�����D3�	:%%��.����͐�պ�!��z�{Y��l��|p�\�z��Z�F�V�^N(�Z�/�F�։�J��F�	�]���}��%IB0�,�����Ѩ���(u���a�NI��󡽽���҈$I��[�;��V���r���#�G�eY�Z��J��Z����h�����W��
��=|���^��qf-�ց�]�}ÉHI�.��j�w(D)�	:%��/���B�L�x�CD	$��fee��� ��$>4rJZC�}M$��,�㶔�$	�$�K�C�s(y�f��+����ض����Pl�?�.��fJ @[[<O�C!JYL�)%��񠼼��҉hF����~���G�^�#�D�h\.���x}"�e�G4CFGG������P����R�CCChmmerNL�)��|>ttt��p�;"""��&�2:;;����J�D1��RNh]��b�w(DDDDI)���6�-ޡ��A���u�DDDD�Z6�-�b�#��FGG������P���������LΉ�	:�<���ٌ���x�BDDD���� :::����P����SZB``` n�eee�}�����ҝ��A[[�@�C!J{L�)�8x�^TTT@���;"""��Boo/��%#R�	m�f�Z�
Q\�A���s5��tJK�,���.�eee�$)�!ń��A{{;�~�C!�	��SZ����z�(//�w"""Jy###����9Q��wJ{^�f�6�-ޡ͊P����.&�D	�#�D8�K���N��Uމ��(���n����J;Q`�N4�����AYY233���288���>��%	&�D��~��f���(��M[ @{{;�nw�C!�i`�N��� �n7��ʠ��
%>!�N'�f3dY�w8D4M\hK4���Q����n��;"""�Iɲ������39'JRLRYYY��ͅJ���`�N�p���t: N�V�5�a���/;�Ӊ��R�#""����z������PR�J�Bnn.���  ��ِ$	���{�׋`0���e��0AOPeeeX�`���QQQ���
���#??yyy�j�SzY�a�Za�Z��ۋ��n������������i�^VV���p���� ���C��h0w�\̟?���(//GEEJJJ�������)�����j���zzz���mmmhjj����,��P��jjjX�1�


p�1�`�ҥ�����������z��܌]�va�Ν���EwwwL~v2+,,DQQQ��)�ti4^C��s���������4I���s�ￏ:�(̝;7f5�����o�>��Յ�B3`)>t:�nǎ�x�0A��^�/~�8��c�r�J~���i���lݺ[�n�����p8�RB���M'�C����V�����>m�����r�J{�X�brss�R�,�ػw/�n݊>� uuu��cL�Ӑ^�����3�8�|�$u�`;v���o����\�>�J�Baa!
�
%&�Dt(� :;;9�:���8���q�g`ѢEIs͵�lx����[o��?D0�wH)�	z������;��r
233����}�vl޼��׿�R����@YYY�X�G���    IDAT�0A'����������$222p�g��s���%K��:k�Z���������pR�g4q�9����ϟ���###������ �V+����t:�t:!�2��ej�:CVVV����dBEEL&ӌ\�����W^aQ�ϨT*O���/&�D4U�`��ݰ�l�%a͛7���wp�Yg�h4~������Gww7�E�].FGG��Z��V�a4���.*WZZ�����-��ЀW_}���Y��1AOQ�����q�����p������CSS���g���N�Cyy9,X����Aqq�!�_ ��o��^x{�왑���hDiii�
�Qrb�NDS�p8���$�/_�իWc�ʕ�|M5��ؽ{7�������뛱����٘3g.\���#���G����Cz���A����ظq#���&�)���?����o|#<�=U6�۷oǇ~��;w���-.���r,Y�˖-ñ�����i��֭[�~�z466�B�Ʌ��Dt0LЉh2�`===L��X�r%���Z,Z�hگmkk�֭[�c�����e�3�Z�#�<K�,��+�|��iרr��x饗�����s�91AO&�	?��p�9�Ly_r ����[o����_����NB. ��$iH1�	 b��"@�$IE ��a��ϟ??\����� �������'�@SSӔ_��233QZZʵ�D�	:Ec�������`
�-[�뮻K�.��kdY�'�|�w�y���t���`0`�Ǒ$)CaP��W������.O'�tN;�4L9���Q���x������iz��'9�^�K/�W^y��Y�V�����?�1�f/�I�� 4Ȳ�[�Ѵ;�NsSS��Pb���ջw�P�T�!��@�$IKdM����j�y��ַ�����)�<Y��i�&<��i�DO�$��;����&b���*++q�M7��SO��k��݋���/x�w`�X�}�� � �j������^q�{�}��_Ͱ��K�t�$IG��o ��I�T*���/����g�1�����x�'���sI�41AOb'�p֬Y����)���O�q�F��������!Ŀ l�x<�j">]'�t�fdd�F��
!N�$� ��U*�/_�J?���v��ׯ�+����������B���;"J LЉ($��yOOO��/M���q�UWaժUS���z������M�6lP�O��wdY����v�ڵ�P��Z�h�Q�V/B|�� VP��k4q�Yg�.�G1��߽{7x�.;�&�I(777�p�?�����e��>6l؀���h�z�&�x��t�����3���/�P�gϞ�$}�� �)�3�L8���q�%�L�2e]]������p��E�$����7�Di�	:����l���w(	g�ҥ���1w�܃��+����^zi�ٛu 6ɲ�?�v�UB~0,�1�~v��MD,[�t).��r����!�26oތ_���lM�$s�g���o?h��`0��������~����.!�+ �����o!D�?"=�c� ���% L����`ժU��w����Ig����㷿�-�}�ٴ:���QVV6�b D�:���7!�����ۋ���`��7ߌ/���ɡ�!<��3شi���	��$uȲ�{�F�ߵ��	_ i�������?�����BFGy$���Z�p�	}���n�y���Of!���=I�F�]�_���'�'���o������l6G��$i��)����޽{��lZ�h�N�V]qL�'//�_~9.���D����ڵk�=�H+���0�LP�T���b�	:Q��x<0�͊	e�;ꨣ������������3�<��^z	O�DԠ$I�˲�����w�aPL������_-I��P�պh�"�p�X�|���#�2�{�9<��S�nRc��-Z�Gy�k���uuuO	 �$�Ѻ���f+�xX�h��J�c c�z���*�t�M8�S&}�Ӊ{�o���,F�4L&rss�
�t����ׇ���x��p$I¥�^�n�a�ݑB��ׯ_������� ��D}}}�,�S^x�z߾}�B��+ϟ|�ɸ馛P]]=���ڵ��r�t�ا&�	��s��ڵk'-Da���裏����Ҵ�w����O�$��_�5G���$���qY+V��]w݅�����B��{�1n#n�F�n����Á��N��(����}�݇�O?}�~������{�o߾��F%Iz6>����7k�&�%K�+�� ��o��t�������{I�͆5k�`�֭�jRa����Z-n��v�w�y��{��w��C)m��J��e�Ν�Z�	���f�$I�@Q��ݦ�`�5�\�K/�tҊ��1n���ߎ8���������q'JqLЉ҃��CWW�������?�8��S�K�����������:F!��*��޺���Y6���Ԝ-I��q`˶��s����t�xY���O��g�e���0AO@YYY��/~��+WF��t:�裏bӦMO�!nkhh�8�A&�Ϟ��
����-��?<鴛��.\{�hkk��0��N�CII�A�Q�b�N��dY�����Rz@�sY�x1�x�	���G�k�.�]����O�)��͍���g3�Dv�I'i(I�= 
B�$��/ƍ7�8�h�o��{�~B�q�=����c����>����Oq��O,l&x泋�s��L�$�jjj�� ��צRp�j��n@mmm"M���())�F��w(D4Ø��.�˅��N�|�x����<�L���Q��NRج_�������!&�&�ŋ�x�UcۧRp>7��#)�X�&�	��ÆPRR�ϦM��nݺ��F!�e;f=�$�hѢj�J����D_����ӟ�4�������[oŖ-[bfRP��(**���2%&�D�'���v�=ޡ$�.� w�qG�]ll6n��6l۶m\���$����>�:�/>�� �U�333q���3Έ����\u�UJ�w���p�B<���(((P<�r�p��w㭷��.I��������&!I�TSS�} ���^�h~��_���L�u~���v�}��E�8�(�0A'JB����kzbժU��曣^���݋o�qb�q+�����)1&�e˖�|� �j�$	�W��7��.T[[����c` ���1AO Gy$6l�uk�����G?�޽{�6;\͋��,Y��hY�782�VTT�_���X�h��k�� ֮]�7�|3Va&�ш���I� !����(�	!�t:���������+����_���-[�f�������h4����O{�����l��6 ���<��c��#�D������_��u)AW�W��;�0��7����777��K/����$�+LΧo�Ν�dY��$I���q�e�EM��j5~��n����N'Z[[���?��)ň��Ekk+��ۙ�O��_<ir��?�	7�x����i�Nw*���B�����U*�J ��>� �V�Boo���*++��3��d2�(RR�v#���������W[[�k��N�j�I��Ǭ��l۶ͭ�"��1O�����T*~�ӟ��s�U|������_���h40�LQ6Q��:Qr
�������p�CI�>�뮨׼��>���&/������;�e˖����B��BmeeeذaC�����p�W��ȉ4��V	z^^^|�Ũ�;v���O��$����{͘c�9�<!�d ���r�-���K�{<\~��hll�e�I%##�����Ȉw(D4ELЉ��V�===��6�<~��_+�B��G��/�8�y�9�����U��N��ǘ*����~��*�����_~9<O�+&�q������b��Ŋ�mۆn�^�7�pe}}��1
1����|U������t�M�������b���K.�:%�<���Ɂ�d�lDI�	:QrB��M�~�ӳh�"<��s0�x���ꫯ�mnW�է���6�,�4��L�� �j����3�<5I��7q�m��E��DJ��b�$IX�n]��|ǎ��<69�K�t�����аM�R �q��W��+�����d2a����`>	!l6ZZZ`�X�t����s�z�hkkCkk+��i*++ï�k�� y䑉�y�$I'39���K�K���  `�Z�� ��튯9��3q�u��0J�$A��+p�i�)�khh�u�]7v��_������6�,�4�s��]B�S�Y�.��C=�7�xC�����q���s�� �BKK�����'�L
��������.}�)���x��GQTT�x��'��8�}�,�_���k�I�i����!��㡡!|���GO�r���(�)��/_�?�я�uww��믟����uuu�"͸���=�$�` dY��w��(ܩ��u<�a�X���
���p����,����Ǟ={Ҫ@�L[�v-�>�h�s�7o��O?=��Y�ќ��ؘ~{{�ICC� �����k���n��+I��~̛7/�!���N�KJJ��#�(���l������p�$I7��ս�	���kp p��-�܂�&�N7�p�-[�����Gww7���'n]BDDD8��c�޽�w8I��sύ�;�֭[q����m2n�����	!�
���⦛nR\ʑ���_��,F#)���T*<�����ˋ8q��7�[o!�XWWW�xC�1���?B|�8���u�]���Z�Raݺu��ɉu�I��񠣣���\GGDD����v;��ۇ��n��x����̙��n�M�\kk+n�喱�v _۽{wG�����1t��Gaݺu�}�Ν�[n�%V����M�W�^�/�ˊ��q|��G�cI�����x�bg������:t��Ӄ[o�U��Yii)����BZZZ����D�������(��ߏ���x����j5֭[�8��r�p��7�]V�p^}}}C,c���,˗x;���k�a��͊�/���G���L�,Xu��;＃^��,vI��\�}�C}}���<t����'�T�{ꩧ⬳ΊUh)�n����}}}�1!"���v���Ԅ��V�|�x��2���*���(����;���>�$����wcE����s��!�kKz�!�޽[���wމ����ŗ�R.AW�T�뮻��j#�������[�z@�V_�e�f'	���a-�<�{����*�]�f


bZ�B�j����K�,Annn�C"""�����hnn�{̀�?W\q�⹍7��w�����꞉I`4%MMMvI���l/x뭷*�`�������'�1��\����~K�,�h�ew�ql6[�Iq	�R$!�,Iҥ �����SZ������o�9�!�!,X�'�x���w��<��׋��v455q˴Y�R�p��B��E�3��x��G�6�p8��,8�����I��7՝��x�G��}��8�b[�I����$���?���֝X����NL�i����$�b A �<����_�:�/_��R��`�7��M<�����X������~�?��9��=^x���X0�O~��\�PӨJ��n[[�/$����� �����͛��{�)�]�v-�z}�BK+)���x㍊	��l�����6�����ޘF�����}!D����o��"�f����Ŗ�F#.��<���8��y&"����z��ى�{�r/�Y����k��F��/�0n�$I?޹s��X�F����]`_���T��������bY�H�}�������E�!p��������l�$}��Γ���@���>��|޼y8���cZZ�����ի��SO�.��w""JHB�|>��f�߿�F�E�\s���f����o�6���Γ�޽{�$��g�X-\y'�+��eee�/-�L�~뭷B����7�xc\�1!Ě����X�F����ɫR��Ę��SO=����k���h�exi#;;\p�z�)�Q'"����za6��o�>&�14g�\xᅊ�|����c�j�Zy*%������m�6mڄ����~z��^{mLcK)����8�c"�].��'>�766>��hF�ܹ�# �ǰ/��2���#�����K.�ehi'##���7��SO�{����Ss""�X�x<hkk���������k��h"ڷlق�۷���kkkk�c� !ĝ�$u|�=z�!Ȳ��k_��Ν��RY�'�$�ꫯV<��3��b���B�	!"?Y���n� �EG~��+�[�j�
;D�v�}J_~��{,֭[��.���:ńhmmESS�Ng�CJK����g�����'Vm�mll\ё^cc�@����ݻ��-��J����ѡ�jjj���%��O>�=�XD��b�Yg��^#��MCC�rJ
�/�
��B�6lP�����O��'��h��#I���PPP �V�p���F�Q\�ED��̙��/����8�S�NZ��/��N;-����^�C=4�����w#:R�X�x�; N���2���[�ɲ���;---�qF�t:ݎ;��H���.�L�}Æc׾صZ��1�főG�,���P�?좋.Bfff��"�Akk+�����p""�������s�[���Ϗw8i���B����ų�>;��u&��O��[� ��ۋ�^{-��J���իcZ�J�}��Ŋk�{{{�y���$I����O-)�lܸ1(Iҝ��;w�>�藓��o}�[1��B��t����zHDD�D�Vc�ʕ��o�{��e{��w�G��j�*�T�)�ƍ100:��˸hv466��)t��3ό;��a2�bZ�J�}ժU�������B�V!��� �t����
�����]r�%��<(v�n7�������ժXX���h,�N��}�kذa���j`ӦM��[p�	'����v�t4�����~<����c!����������T*�] ��e���_"�h�Z|�;߉uh))i3���"�|���v����6=Z__?��h�I�t����Z�m*++�r�ʘ�Eʼ^/�����ڊ��A&�DD�h4�K.�����V�;�'�x"�9��w�}x���Z��7�����������c3�B��#:Q�ڹs�~ �����y�����??b}:M_�&��s������*\.W�Х��~щ�Z}}�� �:~���{
�� `pp��ͰX,����QYY��կ";;=������r����h���;O���_{�?����;R�B<@ @ww7�{ｈ>yyy8��cY�I�]�$��5�,��W�w �x~ǎ����f�B /[x��������O�Z�$�2�����ڊ��N�S'"JCZ�===x������	yX�t)�͛���'�`߾}�c!įb�FCCC=�-��_~Y��>��LЗ-[�������۷���'t($Iz"��Q���?
!�	�_��׈>j�g�}v�c��B`tt]]]hmm���0���(!� z{{��؈O?�CCC�������b�������E<{�$��>��c���>+V�@IIIL�J5I���q���6m{�~}}�ޘD1�m�6�$I��T�7oVL�N?����E����a`` ---�����w"�!����FGG��ك��A�G�D��(n��p8���vR{:fAQ��@7p�����_ l�����'�t�J�SO=5��f������B��ޔ2$I
o���ۋ;vD�9��QYYӸ���A���������c�IQ�e###طo����p8�}˗/G^^^D��o�	��:� ��X�E��e˖�����o��8@m0��&��e˖��� �����'�@�Б���ZD'J)uuu�����o��G�$>�KR�f�---B0�wHDD4	!|>z{{�{�ntuuqFT��v/��[o�=�3wNJ}c��ܹ3�OMM���bVJI���NPl�p�x}۶m�Dq%������VL�;�B�    IDAT�D3����b��������wHDD4�,˰��hjj¾}�8�=�H��c�=6�}ppp��EI����QJilll�I���7ߌ�#I�?��}�����v�}�Q�X��W#:Q�z��HV��|�	���/��d��FVO �������\�*.��j��j!I�EGDDS%������� �������#�<RqW�-[�������S)Um�E��,�k�F܏�\�7nTz-DR%����;wnD����ǎ����>:/^�	�e �u�ֈ]�VcŊ��P�^�W^y匽_ ���w�}����A$"�e�,��t���^�7��P(�����?�����<�)�Ȳ�Y�R� ,��ߏ#�8b\�+V@������%�d�T	��+۷n��^�/i��,A���p�7Ft`�>}?��O0�|�s�v���?�x.�4���+_�
ZZZp�M7A�VC�I�KQ�s���������˗G����q�W��eL_���͋/n08p�=1A�����G����x��Ԓ�.��c�Ql���T��*J�,��R�����fX,���XK�,�Kl�j����K��l6�{�1����͛����k֬��`@nn.rrr�R%]�"���[n��a�XX�-M��j���D���֎�iE�T*�^M?� p l۶W\qED��K�2A?Iu�t�҈���NX,��J��0i�1�L�n(>��ӈ>��χ�h�uhII�$�z�Q��~�����aDSw�g⨣����F__���XX��hdY���@[[��݋��&�i��#�DFFFD��{��uuu1��$I���W�N(�ntpI�����aΜ9�J����6�,(J[�l	 �:V��A�Ra��ű+i�x�X�p���_}⚳�"I~�����p8���DKK,�BM ����Fgg'v�ލ��v>�$ �z�TWW�^��Ľ1�Y�����bϞ=}�9��=I��/\�P�����(]�t�t 8ꨣbL2���ۭV+y�G3}�w���<�ߏ��!����l6�j�rou"Jk^�سg���a�Z���ƙ��80�b�����N����+Me���Ciii,�J	I�]� �w�{�aL��D�-�Mss3�~?�Z�,�yP�f���Q��?��Ӱ���s].���_g0���Ƶ�T*\t�E���~6��s�\���CFF׫Q��������":(��ﮮ�q[תT���eL�P�8
 ��ݫ�a�����eLI/it��J�e�����U*U��fJ:�ng�F������#�9�;�s������+���Ͻ�����{�M�u'�|2{챈���:���/�4B�v��v���ߏ��,dgg#;;��:������e>4-*�
��͋h߿��������X�D�EQ��<�s�p�B�����eXI/i�@��?������|��X�D�cǎ� �B�J��;�I�A�|�Ɋ�/��rB	ڲe���#��������N����hjjBWWl6�{QR
Ass3��݋��n&�4-0�MM��=5�, JD�ܫ��]�^Q)���%�zEEED[[[��áݻws�Dzk P
D|6  Z�%%%�f�G������a���q����x��q�=�D�;���m۶�M�}�N'�N'�����������b'D��Bۢ9�N���7�^�%K�`ŊX�d	


�������𵶳�{���G}��۷'�C�t�tO D�c1AOcz��q�֮�.~����D�QtI����zD�wuu��B�Dt��"�h�$�4 ���Q�S^^�=�h#�[�n��j�q4S��{��?�i��/}�K3���,�f��f�A�$dee�h4";;j�zF~ѡ%������z��i���L\t�EX�z5�����������_�2V�Z�Պ�7�^���q�-��p��ݓ�؎;/^l� ���L�g@R�����T����T��!SJ+�$u����c,^$����������8��Z���80�J����Y���с���C*pGDt(��z��������-9_�l������?�q��<���<\u�Ux�7p�'�N�tP�����������Fi��d2A���2���#�&�I�}�H��
?��6J^\\�`�MMM�b���_�g��㏱t��qm�$�#�����K����b��`O��XY����e^�V�###��E�V��s�=��	 ��믟�P ^x!֬Y����f����c�=�����3MUQQQD������H�X�e�S�c�#�I����¨�[)RR$�ў��=�S�DiC��i1<<��'///�!%�Ѩ� ����%MO{{�b��f5AB�����h�Zdee��X����CY��r�022��Y�?�{.[��s�⹙�)u���;z�$��o���ß���yO�������q�Su:]dFFiE���>���X���LЧ!�t���^��Y�*�J5������r����9��t�٥���B��i�h�%���ձ�3~�V�V��$!333������>�N�����x<3���w�b����k��6#?���>��Ӽ��[�{�n�����{�2�{�	5i����+��Pڐ$)<b�fȦ')���\�����JOZ�vh�2V�5"A��YJw%%%�흝�1���D�9�K����hxt=T>33�U��X0����j��n�ܣ�9�����|�ͨ�^ӡ�h�����ZS�J�x �s����{�		�m�ƍ�_oA)E��� ���	z�����h�{Y���Svv�u����Gi?O�^�!Y�#����+��~?FFF022�J�����;?�D�m�(���H̶B+//�:�h���<���q�a�����Gmm-��ك��a�t:����-���UUU�����?��33MN�w҄߷���v���A��1����HУM	�G�$I�U��bn˖-�ŋ�(>a����w|u�?��L:�B��nIh�� rT=�pr���w*'*��ʩ4��
(F��I)"�C��B�!=�������o���dwvv��|<|����y��f^�i�^�,**Jq��,oc6�QZZj7!QDD��*�I�l��׮]C@@�-�����z%�r�,�l6��� 999���/7~W-�&�~���*�
�O<Q�1�$�/���%K��%$$`����ׯ��ϙ0aV�XQ����9J��*�Z��q�l�l6+���:�k�$I����7��0@�K�_����z�'L;{����=h�'��yyy���Ê+�cǎ������t�DT	Y��u[w��n��(�o߾�%���ׯ�9^L&�L���;wV�9�ϟǿ��/�5
3g�T���۶m�q�T9���
�V�i���,��ֿ�������9^Е��PXw�_�&��B���p\�ҳw�^�ݻץ�Yo S�~}ԯ_����,˸p�N�8���t���o^1�>�/�e���(,,Dnn.���4ٲ�(��*�>�������m�yY�|������3�(��߿?�
�p�mw3N�GE��~�Q:￝�]�]@@@�ׂ x���-�)�bq������xӘ谰0�m&��|			HHH�u����Fzz:�;���tdffz��,����!����|M���Nbb��6I�\2#z�F�ЩS'��w�ލ5k�8���|�	���������ٳ'A����U��;�� �;�$Y[�q��U��W�Z�� Qm�eY�����.����zʀ��QWv���
		Q���K]I�ڵѭ[7t����v�?�Ν�dk�7��E^RRbC^TT�u�0&&F�<##�%Ø�w�8t�jѢE��\I���[oa�ҥv����ШQ#dfr	nw�BOD��F.!�b��{�Q@����^�x�8:���'e��*}I�B����-��5��t4�����-Ξ=���t����������NT���($$$�]�vhР�qO�Tc�7Vܞ�����ر��}ǎ��y~���;wNq�֭[3��Y&��7��`�����9^���ժU˶OE�i��o���[d���﷨Vו+W�7j�H�J�'>>^q�իWU��u�^��p}wg�S�N2d����;w'N�����q��)N>G~G�e����A�HLLD�ΝѺu�rC����V�:�zFF�K>�C��mܸ�Ɵ�u�V<��v�[�n��۷����1�{�
�V\ܚ B����ҽ7��I�}�WtG�qԮ]���  Y��Yi��l.w(�(��Z�w�/_V�ޮ];�+�Guz�:�JM�T:�+V� p�g�6mЦM4m�+W�Dpp0BBBj�������,�E�ƍѲeK$%%�U�V^5�FM8ZF��6l��:���?�������;j��T�7n��^�poӧO��;vp��+����`�kT5^q��Htt��gQ�Ui�,˱֟������B����!˲ݒ6͛7Gdd���Cw4C�+Z��AII	JJJ��E�\hFXX��GDZ ˲mV����o���_вeK��A�Q�VNNN�?��w/p�g�+��O�<���уr�{���r��BNNNm \Rďɲ\�zoP���q���?��k�c�e�;˒��o�b��	� ���� 33Ӯ+�(��ի6l���n/88w�y��_�U�j|�$I(***7?� 		�����`1��j�A�b��d2���������ða�p��"..�F�8}���׉�SZ��K�V���СC5�|�fO���R�^=�2��7S���xe6��ݯ��X�z��(���s�"�;GZ�[�,��T*�����Gc��n�ciii�c��ޫW/����m�X,HOO�@E�K�eۍ%AAA�B�5�3�Su�m/))��dBAA
mEDD�O�>6l���]o���شi֯_��Ǵ"$Dy/Wc��t����,�((((�kp�3�\G�)44��SQ�8�ri�!�,Wz�-�2�_��jM��+��q�e/A��Si�,�M�?;�4�3�:���?cРAv���n���k��nܸq��SSS9)�J�kCW���ܭ��e[���N@�^ZZ
���Ʉ��B+.(�"�v�aÆ���5K.IRSS�~�z|��wW��f����l:C�m���~W> U
�lAw?G�����.IR3K"m�t����ׯs�f'yE@/**Bvv�]��
AU�"-J���]�!Sv�؁3fحg+�"&N��Y�fy�2�:t�Ν;+�۱c���PE����5����m��!�b��$�b��l6�za���T1�+i֬��Ç�x��+W���CJJ���U�h�����Y͚5Cdd��>Y���o�����*-��������5�3���ۖ�!Q� �:�.VE[�v��f�{;�+:p�nŀ^a�8�N� --My:j���v͚5��YZZ�p91���O8p ]�t��7r�H��������LY@@ ^x��}�$a�֭*WD�2��0��(,,��'h�� ș�5@�$�x���R��f[w���b[˸u|��\م���?��֯_�]�vA��j�7���U�޼ys��Ue0�p�K'UG_PP��'e��U�k��L���DQ���DBB��1��󚻛����N			�u�� ���� l��Z�nmw̙3g��R㯾��Kŀ.�"�͛�x@3kf?��S�W�ڵ���\�nώ�*X��[��ҿ��L�+�%I��z[[�KJJl���?+�l֔(�0�6l��p���:~����?NT�(��jժF�����p���ѪC�۵�ȗ]�p&��n���r�掟Ԑϓe�`}pڼys�����vY^�k��S�춉��-Zغ����5�"m�$)���-00P�]���oߎ�/*vQjҤ	�ϟ���~�a�e�>&Lp�����Cc�B_���� ��X�g�kG��5�ڥ���֠mm�.��f�-|[�y�e�aÆ<x0ƌ�p�����Ŗ-[�j�*��,��2e;v,���AгgO��8��g:�8���I�������+<܉���	ǎ;�jq�	� �Z�+<������&�;�ӦM����j���������5o�q{�$����k�����G�X�`��y�u/5jf̘ᰫ�����o�>��"�+�"_�(�K�.8p z��e{8`6�QTTI�PPP`��e�*�������ѣG���&ϱ��-��m��\�;y����ۛ���஻���ѣk܅]�$�߿)))رc�m�ww��%dee�N�:嶇���W�^ز��v���ۣ^�z��2�+=p�*�ZN�:e�Q�!I7 ������6m�(��o�yM@?q�dY��坔���� � �璯�f�!))I�'N�V�7���o��@�WV֫W/,_�S�NU�e*<<S�L��Q�#I�ϟ�ZM���7o�A��db2k���_��	��M�.�C���rYgΜ�ƍ�v�Z\�t�EU����4�u�]v�'L������9F��pߕ+Wp��9�kt��X�?���e� ����1|��r�DQ�^��O?� ��U(�<���R�XC�����\~/W�����l�?M�4)����P_�׷8v�;���c��L@�С��1�,��Q.�Y�,㥗^�ʕ+��{�w`�ʕ���/�d�dee����� <�<�L�-6 �l�2>��s��d�V����c˖-~��L�0d��5Jq"!g�L&�ܹ)))��矫=	��8x�b@��t���{�~��*V\\��puZ�+c4��9sƥ�!e��HJJ�t l �C�,wA���`�� p��~?W��t 8|��]@OHH@�:ulA�� ��ȉ':�M��/##999j���N�>��s�b�̙�	����1z�h|��wX�~=>�.�ΎGMMM�{��s���va6l���W��Ξ=�6`ݺu�����ܜ�-%%6lP����m޼�'OV��1cΟ?�#G���sDQČ3*]{��o��Q�9
�lAWGzz:������W�$���h����zU�����[��t��U�{��y]@���Ft�޽���� >T�6�I�Zo:Z�h��s��!���z)))hٲ%ƍW�q!!!9r$F���ׯ�_~��C�p�ԩ*?	

BӦMѲeKt��	�Z���:�����׿��Y��iM�6Ő!C\҅�����]�v=z4����}ֵkװ~�z�^�ڥ]��ɥK���?*�����b���x뭷����𺍌�Č3p��w;<OFF�K�o4o�qqqv�q��Y���+--űc�йs�rۓ��j]eC��J�H"� ��=z�P<���ê��K�*����ϊ�{��Y6����t�iii��f�T#�`�ώf�ݿ�j���y��!22Æ���u������1x��	���q��u����d2�d2AEDDD $$u��ALLL�k��������p� ����8Çw8gEUɲ�#G�`͚5زe�_��6l�Ç�}�݇ƍ�賬k��Y�?����M~�EK�.E�޽[����1c�<��Cظq#�?���,�����8t��C�Ett�m��J��{���#G��e�?R��~���.]��� Ȳ<�~�h46`[�X)��رcj��3�*�gff�̙3v3zv���(Z�G
���w(�Tf4�-ܭ�a�X8�w5I���ӧ�x�'�����5�Yw�ܹs�4i[��)��t�FU\�v[�l��ի9C�-�'OƠA�n`%222�~�z�Y����.�����vӦM��VԬY�j�gdd`Æ�-ώ(�:t�⾃��<t{�w�ƓO>i��W�^��`XbbbȩS��w�?"I�H�þ:u�(���~�/�뭼*���={�zLL:w�\��},���,�c ���S�Nv�=z���j��3dY��ŋq��L�:�ұ�jڱc�O����<O�B~�l6c�޽X�~=�m��!.����͛7�� ��={6:t���(�    IDAT���seY����]�ӡcǎ���r7���~�Mq���}�b������ѡ�����o� ��֟���8$q��ݪ��K�6�SC�<�+g�����A����<�4�������?sڵk����իWc�����#//3f���O?�pN�����ѿ���Ė-[�kH�$�۷/��"���Y�f1���ƍ�<y�ˇb,]�{��u�g��/Qܞ�����4���*'I���c��nݺ�&�E�~�������nk0`��1�,3�׀������ƍv���뇀� �����P�ov�F��5�;��u�t��/��ܹsx�G0e��'�1��HII��aðn�:U�M�'??)))x�G0b�,[�������z�/_Ʋe�0t�P<���X�~�u�)RIZZ�|�I��,ۺu+�}�]�|�U�ƍ.���?�l6��|t{����{ɲ<:99���ʐ�x�z�֭[W��꯿����L���^���b�`�֭=zt��111�ի~�� � ��J�
I-�$Mn��_�>�t�bw����9>��dYƖ-[�m�6�}��3f�v�Z�ם�������]�֭���+W�`�vۯ^�8eI����T�_��~�-���pv{�9x� Ə�ٳgC��U�3dY�ҥK���|�����e]�ٺu�K�EU�w�^����M8p�@̟?�:�8�b��WS�Y� ��a�����ޫx��i�&5��9^Ё��yV� 0j�([@p�N�k���vZ��H���!aaa[_�1B�b��ͪ��O,�mۆm۶!..�z�BϞ=���l7N�&�	���ػw/v�څ�Ǐs��v��-[��24�ʕ+����.x��q��q�Î�,�H�:{�,z�!�w�}�8q"�4iR���ٳ���[��7j���w�⾢�"v�����Rl߾#F�(�=&&��sO�@�8�}�^�(�rS���p������j]��+�/����/�MҫW/4h� �/_ !  �� ��D��^�����n���4VM�$lܸQ���ҵkװz�j�^� P�^=�i��7F�z�P�^=#**�����b�L&dee��ի�|�2222p��i��%�c��{\�~�7oƚ5kp��IO�C�a�X�f��]�F�ݺu��`@BBbbb���<dgg#33����޽{q����ԵkW�������g������٨Q���F��Wjj*' �M�X�С�7onw����q��%U��5^�%I�ڵk1iҤr�EQ��ѣmc�dY�ضm�Y������A���ܻwoř^w��e}XC*�z�*�O�f�޽�6mB~~��K�)�/ƹs����ɲ�#G�x|P ����:tHq��.]��E����  Ȳ< ��1z ���x�������n�8�5k�(v{����f}�������� ��������)�|�2ù����D>L�e�{+A��C��t_RRR+�
#UȲ<�&�kԨ���owLNN�o߮vi>�k��+Wʎ7����.7vI�g۴i�bi�~/Y�������t��%������yk׮��d��>t�в��Ȳ<]��ȭ���Ag}��C)N���� �xm@��>�Lq��	ʮ�]'$$�)����!(���c�=�x����ْCDDD�B7n�P\�4$$?l���,�3mԬ���b���[C��ԩ��#G�SZZ��˗�\�o��~��!=z�n{|||�I,dY����bլ�\O���۵k�������|vo'"""r��>�Lq��<P��,5�"��5��~��'�Nl�q�F���"^���O?U���c�!$$��2Fŗժ��C��M �������'n-�^�W_}��DDDDnp��9�ر�n{XX&N�Xv����K���儛7�o�����a̘1v�ɲ�g39���֭[q��	��4��q��nzB�ӵS�0r)�N!«��]�tA�=�+,,��-Z���d�M�4���e��[= ��� �m}����l���<F���adY��ŋ�=��㈋���E�A�ɕ4O�W 4��3^x���>��sdgg�Y�_9u��m�f�=((�'O.���^�W�0�4-999F��y��mڴ����펓$	|�����:�� �c����v������O��t�N�S^��4K���&�3f����e�9�
�����]�t)�i^RRR�j��K�����>ps)�iӦA��ƍq��I���i>�eY�ܹs!˲ݾ���/����N�@����:u�$��2ܚ9�nݺ��?��x��ŋ����fyDDDD~)##)))��f̘Q�+t�,�o�V՘�`�(��X_W�SV&�	�󎪵��� p��l޼�n�(�x�W�~I�X1v�X���HsJJJf���pӦMCTT��q���;���+5K#"""�k��nܸa��iӦ�ey��h|D�ڨz�Fc8��qkb������l�-[��/�X�� .Dqq���f͚U���s�ĉ�j�F�����L���ӧ���x����QZZ�ViDDDD~/''~���G}�[����e�]�N�R�ڨz$IZ�����/������._��O>�D����O�/:�0n�ĉ0��ײ,�b0z�U9G���
��������bƌ��nڴ	{��Q�<""""�b�
?~�n{`` �̙S�k�(���t�`U�*����
������ދ�*;g��V�?� �}���D@@ �̙����& _q<��� ����f�^c֬Y�[��ݱ999�;w��ps�3g*�dlѢ�y晲������j�Q�%%%��6�<>>�����ݲe�o߮Zm�����b�+����%_���(�s}Fm���/l}����wo��o������*�����*8y�$>��S�}�ƍ�]w�Uv�?�z�C�FUb4�%IZ�ps���s�mش�����9s�.ѯ�d0�����7x�`�?��A��=U
�����c؞�$%%�駟V<v���X�n�Z���/Fzz��vA0g�4o޼�%:������2ADY�� �κ��矇�`P<���^�����*�/�d@��>��V���ϖ[*@���5��I5III=A��  ���Âhw�k����/�\!))))��i�`2�������7�@XX�uS�(�_'%%�R�H�c0 �����a�p���+�n�:lڴI�����tI�0m�4�u��`�4nܸ��Y��q�
�r�^��u B �V�Zx�wP�N�c%I/����yFFF�ϟ��/11s�́(��GI�6t�С�jR9��yY����NNN�̙3�=w�����g:psV���ߐ$�n_ll,>��Ԯ]���EF�q�j �֒��7׮�={6ڶm�x��E��o�>+$"""��X�j��!�}����)S�njQZZ�C���W�8������%�ƍc��egݷ1�L�2e



�,�o�t@��;w:\�1!!,@hh�uS�,˟�~�����(n��9N��_D�>�Òv�܉%K��Y"9��^É'�=���x���nj%�m��w�$�0�#�VZ�n]�������U<���^R�_����: ����عs��:`��-�
�;�^?B�����`h`'�&�m�'OƘ1c�?s��DDDD�����׿��p8��>�ѣ�uZ������O���/�%��������I�&�����ذa������eO��Z�j��?v�mz���2eJ���̂ <�����jE�����F q�mO<��x�	�㳳�1~�x\�pA�
��aÆ9r��� ""y���a�X<]�Mrr2>��C�nӒ$a������om�dY>e�X�?~���u����oY�_�������~�N�x��;0y�d�h>p����u ~� .._|�6l����ĳ�>[v�IY�Y���/�U�?HJJxk��(�G}�<���&�	�=��9�V��סC|��'�.���4�s�Ί3hyҀ0o޼����H��Y�fa���e7_�$龴��_T+�Ǎ;6��~{[�I�mQQQX�x1�z��{�?����o(**R�NO�R@��.�V׮]äI�������w��x�w�.!Ȳ���`�@��+�����럒$�;�
� `�ԩ�yii)�{�9�s""""/�e��3�����^z	�Ǐ/���(�?p��k$''Ǥ��[6������O?u�Ϝ9�I�&�M8��
�����q���(��ڵ+�.]Zqy��EQܫ��[�R�j޼y��h\"� @pp0^�u�7N�=���~��+%""""WZ�|9�}�]�}� ��^�/�P���� ��9cǎP�Pc0:Z,� Y�5i��1Z�P�5�/_�������?�T�L���: �8q���?.���|��nGA��Q��Ct:]����}�,O�n����G}��C�*����i�ƍ��IDDDD���V�����1gΜ��� /���o�СC��7�A���4�� l��K�.X�b��	�\���'��ŋ*UJJ�2�@jj*{�1�-�5�g�}����Y�S�F�gݻwS|#�c4E�0 �u[�V���_ 99Y�=�3f̨8��������o��E�9�?h� ,]����+�y@iii��h��}@bbb�^��J�� lCt��~,^�QQQ�����Ą	p��y�J%�6�@ZZ&L��k׮)���o��g�y����,?�����`0(� �����a�,˟��n<x0>��s�O��f3��y�_�^�R����H%��>^�uȲ�<��)))���;�n�'��:�^�^�6m"U)���{���R��,		��/��_|AAA����?0a�dff�U*U¯fqw�I�&X�h��� ?���O�^1̗x3//��?�����uzA���,�o��Ŕ)S0v�X�������ɓ���?�Q�W��,��|�𗪷z��ѫW/O���l6�7���3g<]�K5l�S�NEhh��KQt��,Y����Gyݻw�t�L&�ϟ�s�7�7���?��̔�Ug���ಓ�����B�͚���>|8^z�%*�X,X�h�.]Zq���� <�����*�z������2�c�94  ТE̝;�Z�r��#G�੧�r�f����,��DGGc��ر��c�������6m*�]��S�(>�����;z���� �,��E��7o���ի��?����tw��<�SSS1m�4���SEL�6����t)��f����ػw��Kq�^�9s�V�Z�.�����cƌ())�t).��3gj�d����q��O���s��q{v6�#""� ��`/#�2���}��/�ҥ,X��HǍ�G�ŴiӔޭ�e��cǎe��HA����
�ܸ�aÆa���~�lݺӦM��`@�,kG�Y�_����Wz���,�S�;v�mEj��hl,I�k� <�2�&���1q�D���wإ���;y�d�C�^U��c�*>u����t,]�ԧ[#A��q�йsgO�����1~��WO��V͚5�O<�J�bU?~���_�=�:t���R �|��G��ɓ�.ŭZ�h��{�Z�F"""θ\�3=88��P�ҽC�-�����Ҟ����X�p!����=�JAx[��>�WM�F��Y�� PnR���x̘1���R�,c�ҥx��w]r���5n���x��gv����l̝;6l��K�;��2=---խ�z��h�'�� <�����d̜9�7�V��ܹs}�f�������x!22�'[X����{�I� �������/)--E^^��o|�5Q	�u���f���9=t�S�NX�l�m��j@��p^��u�\dd$^����3�9t�f͚�����< � �=z�h��������, ����ēO>Y����|L�>۷ows�ޅ�$''c޼y�_�~��<xs��U�-ɲ�F�7RSS���PHJJj%��dY�' (�P�~}<��32dH�7�EEEx��W9\5���-� 7�*x�f�����C��+O���f3����]�CBBQ�1��!]�A�c�=�'�x��>/--�ʕ+����#//���� ,x�СC>�V� �^�,�Y��T�߽{w<��s�m;y�$�}�Y�={�m�z+t/��^z��R%I�ڵk���ҥKv�A�#��⼼�o�u2��c��8q��$I�A�
+ DDD��Ƅ	n�}��_�ԩS��Pjt�e��Xݿ��X�,rssU��έ<\A@TTT�=�|���\�y�3�{�ш9s� >>��㲳������o�Q�P"�W�$���1��ȥS�N�f�y�,�Oh_qbb"�z���<�e+V���w�t/3r�HL�2�O�KJJ��7�`ɒ%��S�)� V=zt����6 �x@B���j�¸q���#� ::��ϲX,��O��{��=�	wt���R3��{8�*--Enn�j���kkbYj���pn�LHwE@�~C�w����ԩSq�}����K�.��?ĺu��_�&�ǒ$}y��1�/1v�؀���> �����fRm޼9�x�	0��R�J�]���3gbϞ=�)�G0�{����*��l6��i�&,[�'�<`� ������c�M$VA����EQ��h �k���������_��W�����sO�<��_~iii.��?�3��&����B��\��R�Z-�|U��x��W�k��=44�j���Q1�{�=z`ƌhԨ�m��~�:���k,_����J�� �HE��#G�hff��ݻ��%I�}� �B�٭ڶm�|C��t p����~�y��!''�e�t/6p�@<��s�WO��M9�,c���X�jv��U�/�Y��
���$I�۵kwlժU�^	���Z��n� �#��  ��5
C��Ҭ��������bQ�?��+�3�(sgpa`Q������׺���k�&=$$����+`H��j�O>�����U������ڵk��7�T�P �����eOZZ�9W�|;:�.X�N ����]�0�UHH���1c� 99Y�;�O�ƫ���C���hǀ�����0q�D<��#U^��իX�n6l�p�/��L�pL��DQ����×j�-�C�q%%%��I��^�,˝A�[���ի��b�ȑUZ��9.���x��|��#�3�W�-�,�sWHg`��u���Z�n@Exx����5��k���y��x���ѣG�*�����X�n�m�V�V�L dY��QY�O����m}��	�r�J�(�w������?I�0�rY� @��c�С:t(����t�7n`ѢE����0�$tѨQ#<��:t�m��u��il޼;w�ĉ'�kip�5A�dY�`�e9G�ouY�#EQ�e9@�[�4P��ҍ7F�޽1`� $%%9����O?�w�awv7ru@gkbո2�0�T��C:�yո2��������v��w�]��	��T5�ާgϞxꩧЦM�*��l6c߾}����k�.dee9s��y��%�r� Y�yO^X�  � �ɲ\@AȲ��־�EF�}�����ԭ��d2��/�Ē%K؝���}L�f�0iҤ*M�Pѵkװg��߿�Fff����\ll,�F#�t�=z�Y�fN�����������/��qe@g`qNQQ
o`%X�#Irrrj�ٚ�W<���G!�ـ�Z���"ҽ� �۷/&M���-[:�^Y�����={�����HMME~~��*uL�q�HJJB�n�еk�*��[��� %%K�.e��b@�Q͚5��?�aÆU��{E׮]Cjj*N�<�ӧO�ĉ�x�˺���z��E�hݺ5���ȁ�7�?��>��S>|�%5��*���zj�X���-���S��.�""##�K�IJ׺3]^�ՠƄ��z�(�w��x�Gбc�j}�$I8u�~��W�:u
�N���ӧ��{q�  PIDAT�����`$$$ 11�Z�B�V�`4o��#���X�jV�\�`�"�>.66cǎň#аa���b��+Wp��\�r999�q�nܸ���R��~aaa

BTTbbbP�vmԭ[���hԨ���k\S^^���[�X���{�+:K�T'�3�׌�bA^^��,ٚX3���W��HUz�=\�;�_1�{7�N�q�ơ���n(+���������DVV���q��۲�'�[���Att4j׮��">>qqq.i�����_��k�ָ7�ǀ�'DQD���1r�H�����iJ��C�a͚5زeg?���t�(..FAAA��ek�k8�y���3!=   ����5T�%�*}�ʕ���U��w1�{���H�{�1b�S�Ե*??��=V�^���TO�㳴�y��F�$a���ؽ{7"""ЧO4]�vEPP���8Y�q��Ql޼[�l�իW=]��넆�B����&�N@@ ����4&�׺넅�\��v�:ù�X�����������>S�*�g���I���+Wb�ʕhڴ)��:=Vݓ����s�Nl޼�w�f���a������;�DϞ=ѽ{w�fiTÍ7�o�>�޽{��qv�KRAu[�X��d29�`���=$IB^^JKK��Zw��Z�EQDtt�ӓ�R�$IB�&M���+�_�l��}T}����%>>=z�@�^�йsg��������={�g�:t��\elA�sؾ};�o���rm���HJJ��`�w�ᒱ3U!IΞ=���49r�������o�%X�'$$�,�uwg8w됁��\���jղ���k9jIg8wQq��%�={M�6-�oɒ%X�|��*�mU�5B�#33�V�ªU��6m� ))	���h׮���U�4����N�Bjj*>�#G��A�l؂�Ahڴ)ѴiS4j��7F�P�N�'�2�L���ƥK�p��\�x�ϟ��ӧ����'t^��t�su�mIg`Q�$I�B:ù:�ο`��kݽj׮���z͚5�,�x����7�x�,�ǖt���-[�e˖hܸ1���� ::�鹤���p��5\�t	����x�"Μ9��'O"33��a��tt/����r_�u

`�X I�m�w���{�	� 0��������,*�e���		Ahh�������W�vm������z�jO��7�	���߂  ((aaa�$��p�d2��]�D2�CK�]ܽPII	�]��u�DQd`QYhh(���XT$"""8�@e��՗���Y�fqyS�����l6�l�Ľ;yHAA


p��EO�B>��U�|�Zc��<�׺g��]}�DD���������HЉ������4��������HЉ������4��������HЉ������4��������HЉ������4��������HЉ������4��������HЉ������4��������HЉ������4��������HЉ������4��������H=] ����h����v>�Ʉ��,�ΧE�(�aÆ����ի0�ͪ�Skj׮���0��WTT���l�ΧEAAA���S��W�\��bQ��Z���P���k���	:�Ո#мys��w��e,^�X��iQll,�qUϹl�2�={V�sj͈#дiS��w��|��G��O�4h����爵�>T=�֌=�����ٳX�l�j�#"�$vq'""""""� t"""""""`@'""""""� t"""""""`@'""""""� t"""""""`@'""""""� t"""""""`@'""""""� t"""""""`@'""""""Ҁ@O@D����&�I��y.��$I�?I�T=��L&^�*�X,��=���H�?���b��ED�i�D�VǎC~~�j�~��j�Ҫ��<=zT�s޸qC��i�ѣG������.^��ڹ�*''G�k=//O��i�ѣG������Ο?�ڹ��<�]܉������4��������HЉ������4��������HЉ������4��������HЉ������4��������HЉ������4��������HЉ������4��������HЉ������4��������HЉ������4��������HЉ������4��������HЉ|�$I�$��e�Y�QZZ��2���l浮2Y�a6�=]��1�����t~E�$X,O�AD~��ȇɲ����Ȳ���\��磨������Ʉ��|����ZW�$I���ᵮ����=������N�:�.�/H���"R:����H��½����z^XX�ࢂ��b��� ,o�U`,����B{�*�7f�<��3M�6�[o�Ő�f�$!//���D�*t"?P�\���b����Bz�*�W\\����r�,H����>�r���hL�4	� ض5i�,@ݺu=X��^��DDjc@'���E�t׺�Ï��"�t7(**��V| ��Q��\�k�=�����/!!,@\\��U�6��$"Ob@'�#lp��vdHw������yZ,vMu��`�ת�wG�ƍ���o�aÆ*U����AD�ƀN�g8��5�}�������W�V0�p6��Zwg�4h��rhG��i:��MH�T7��&4#�U'���H�T��)d�:=�ի���"~�W� "�`@'�S�&6��մ���dbp����ʲ�H��t��E {5�_q5	�� ADZN��x3�W�<�.&˲�*�m���^#�qUk"[ҝ����@�9�D�5�D~�!�j\���d2����!�6\938{�T���u9<^�+((p�z�| U5����D�9�DĐ~�jaQZǛ��;���^9w_���\έ8�B�ΉH�Љ ��#���h2�������f�,V�֕����u�,�Q����k�!]Yii)���x-�&1���5���fO��	j�M,))���e�3�[1��g���݁�:�ݔ������s�Z/���rNDZ����}Z�hQ�����7t���AݺuU;gII�߷0֪U�k�V����=s��������*_����5:�5�GEE!0�o��f3���ΉH���[���X����5�Lx��q��AV���o **J�s�۷3g���^�(������U?wqq1������ê���Z�n����#22R�s���x�����(��:u*����y�=��[;yvq'"E!!!�={6�u���RTժU+���	� еkW��?�App�G��	�(�^�H8���P̞=:t���=E��᭷��H8����f�BPP�G��	���x饗T�V�:��:!�9yt"r(((�f�B���=]�*ڷo�x,�X�y�~�EQĴi�0`� ����_�:u�hj����;w.jժ��:�u�Y�f�ŵ��3g�w���C�e����MH7���D�UЉ�R���x�WгgOO��V:�����x`��ҥ�Ν���PO��6���x��ѯ_?O���B��?�2��V]�v���n��{����R �OH/))a8'"�ÀND�e햩��KW�Z`�JJJ�ܹs��R\N��TPP^y�����ӥ���hĜ9s4wM�y�x��W��R\N�ה5����x���NGD�m�^�ǊD^�C���OT?oii)�=�Tk��ӧq��7VU^ll,�S���t��ϟ�իW�|��lƞ={�X��.]�8���N�:h֬��
����R���:���'O��ŋn��^���Ѷm[�ޣ��5�R}��Y\�~���b���n��^�N�Q���֭��M�����ӹsg��m��I�v�;�é������}��9����R��Q�8p@݊�oO"����@�'����U5�GEE�cǎ��O			HHH���EEE�����#66V�s�S``���Qvv��=66����M�:f���O�z�v���9�I�e�����L�$I>���Ȋ]܉������4��������H8��yMw�m۪6� �����/��v>-


B߾}U=��ݻ�~B����;5��.]���8y_��D�{��A^^��笪+W��r�=z�e˖���9����v�ȿp:Ո�lV�F���� `2�����]<1�]VVnܸ��y��y�檞��������(�ϙ�����l��KDD��]܉������4��������HЉ������4��������HЉ������4��������HЉ������4��������H��tD�4h0	���W�v� ��u>-��������lذ��7n�S�ZӠA��ܫ�����������^�z	 ��y�F��Ovv��j�Sk4h0�@Ϸ�j�������K=]�U�ѣG�z�"�]o���j� jժ����k�gϮ��9�u���W_}����Ւ7�|s��狌�������y�Z�}Ύ;�[�r�Q�ϫ%o���85�q�߯u"���NDDDDDD��DDDDDDD��NDDDDDD��DDDDDDD��NDDDDDD��DDDDDDD��NDDDDDD��DDDDDDD��NDDDDDD��DDDDDDD��NDDDDDD��DDDDDDD��NDDDDDD��DDDDDDD��NDDDDDD��DDDDDDD��NDDDDDD��DDDDDDD��NDDDDDD��DDDDDDD��NDDDDDD��DDDDDDD��NDDDDDD��DDDDDDD��NDDDDDD��DDDDDDD��NDDDDDD��DDDDDDD��NDDDDDD��DDDDDDD��NDDDDDD��DDDDDDD��NDDDDDD��DDDDDDD��NDDDDDD��DDDDDDD��NDDDDDD��DDDDDDD��NDDDDDD��DDDDDDD��NDDDDDD��DDDDDDD��NDDDDDD��DDDDDDD��NDDDDDD��DDDDDDD��NDDDDDD��DDDDDDD��NDDDDDD��DDDDDDD��NDDDDDD��DDDDDDD��NDDDDDD��DDDDDDD��NDDDDDD��DDDDDDD��NDDDDDD��DDDDDDD��NDDDDDD��DDDDDDD��NDDDDDD��DDDDDDD��NDDDDDD��DDDDDDD��NDDDDDD��DDDDDDD��NDDDDDD��DDDDDDD��NDDDDDD��DDDDDDD��NDDDDDD��DDDDDDD��NDDDDDD��DDDDDDD��NDDDDDD��DDDDDDD��N��]�Im
�(*�I���*�h��o�[��#ۃ��>_�s6��7�t�   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  ��ե/ �����~}}=l�|>o��E���ݎ<�i����<O��g�h���ӯ�j�cuY��acQ������ǡ�߇=??������,��ac &Ё�j�^oG�@��Ƣ>??o___�n����>Z������a���tz6uss�m�硛��n����f�rww7l�x<���\�_�   @�  @�@  � �      � �@���9�    IEND�B`�PK
     ^�[/�i�$  �$  /   images/60da03ea-f7cc-456a-983c-41a209708cd9.png�PNG

   IHDR   d   �   ep�M   	pHYs  ��  ��"篻   tEXtSoftware www.inkscape.org��<  $IDATx��	����k�E@\@���%7P�\A@M\p	Ab��4&�hF�#���W@��\PO܎(�: ��!QqAEAt&����XS�]��gzp�9=Kwu�{�����{/s�A���9����aÆAIII�	ꩠ����ν��ʂ���`���r�z���<*--u�çL&�~��X@6n�4h� �s�=�=��#hҤI��W_��~����5`뭷~��|�M����-[�v�ygǳ�>�,x���U�V9��dÆA���N8!hڴ������1�V�͛7j��/�����/�̝;7�f�m�#1 ���{�~��o0�e|Zh }g<��$��ҥK��g�5k�xެ��x�~���;l���ӯ5j�S���o��VСCİ�e�]����O���ĉ]�~L;�c0h� 4Ʉ�����^z�]����g�����{饗���q��$�Rnֽ{�����w��g�|�UW�ߺuk�p��U�V�7n��/~�&L�l���g�}�G#)�) `?�0lذ�'Ov�
�n�|����}���t���s0�/�K��իc�W%@0H��[p�1Ǭ9r�YF���ш/�b ���_9bĈ��>s޼y;�\��Ga�� �h~??��OS��������8 ���σ���;�1c���^{��i��v͘1cb�I%@0�F���c��?��c�S��󟕾��;�8��@�{�����x��?���t��0|�1�z����7߬t��1M��"�e��W6�����r�  ��^{ӦM���ٳ�U�������1���v�:�Ǡ��H�i��S�LYмys�Urꉀo���_x�۶m; 5�G�S�̚5k9�v�m�b�
��
��>��7_�n]j߻.j[���_/\�`��*��׿r^h3��ڵk��i���sQ6/��FA���8BJ�:�(Uf �m�@�����H���^߁��*M�Q \h���a�0y�W�v7P�4n頠��̓�u�=�g�}�=�E�jH�o��uG�$��c���ْY��W_}���(�k�.<x�k�9��{�t;B:dٲe��h6�e�N���M�"�,/��>��#�/\���#����:uj0p���C���s��+`<�g%B2<�����G`��n<�����w_�򥰾��٤0��uMMK,�#-b��v]t��6BjL�����+ ��G}4X�hѯM��M
+q�������o~�s��m.�Z��� �Z�X�!��A#�D�Օ15�Ĥ��o������0�J�bhïhү� �A��_s�5o��:��S��g1�i�SO=���={����;sZU�4L}����o~ݤ�O?��@@�������?��}~�%K�4iRl�CŐ0�( �(�oܸ�{qOe���+���<Ës�:�,���|���`��
^x�����Ο?�=���٫W/ڿ��q�=�[�֐,GR�)���	�<�v_�lϴ̰�|b⺳��N�w\'\9T\\��l��vYPI3zٴiS�rн�Ң�Q���r��܇{�R����/@�M J+9��lgp�m�}����ѣG�3v��)v�wI.��he�x�ʕ��q��Z�|_V@��
�����w��#�������:��:|�g�o]�"I`����k�IX����i)
,��� ��&�B�50��i��Z��g��S����+�o�5�
sF�*lԥ�}#�+�(5�馛�>xf�����O�*5������́�q�|���� �aǃ��͂'rC7·q4�#���u���%�%p�Qt�f�0�|���/051�Ɇ'F������S�),5L5 դ�?��#��|f�0�q� ��k��e�]�8��*T0������@Z�Ӭ�A� ��G��A��p`��S��F�� �T0��^]%ڎ*#=D��Pc����	���g`d�DH`��'��V�4OТE��MD�8dS�T��~���b�nݺS�L	�8�'A�E���6l��EaiQz0j�(���ڀ�1̖���`D��2�+^	��Ț =�L�Gӵ���=$��:���-@h�/^�U�-"�H�b$� P�sJ{�?3<�x��`�<C�����H��&B�� v�9t�f~��e%5N><�,_0�����#d��P�b3I�rY"݋��	��V~+�����l�
k=S��`�w�� :���{�ed��f��hV����:�$#��L�� 8� ��￿��/\a�嫮�Ԁ*O�PZ�	D�t�B�)���	f6����� �Ѯ|�@PuްQG�}�T�HM��:
��D��vm�(jL�0D贉 0�*�ݒ8�'�n8�L�/o@�1 ��҂��`T�\D���]]#[]�a v��#� R��E��0�XL�U��K^��8a�M�6C��w'iG��(�5?��H�D�!1���C��+-\�w����
>)$@����[Bp�K�k��4=D#�z*�}T`b[P� D?|A�����W$Bq��M����f����S��x~�x�`,j�;� �J��X@T<���%�!]P��E�l�{ME适Ѵ������q^P{���n��
O��``+ �d��E>��S��yru��ʖZ	E�C 
�*;Me&R�Gɫ�*���p�qf͘���8��]�PQ�R)�%U����̓�N?�٥!������ϑ0�w�%���">��
�|k��$�����ϯ�L�qyr�9� ��\F�Q��!E�|��DY2�i�aP4��=}@�H������� 1���a�夆�ݣJ����4���,y"�����u_�����l�6_U�C}� :��o^}�U�m��5���i�1E��
�|I�&�c��nV�\ρ����Q�i�I� ����K�|���`e�1�� �C5��D�>�\��4`�@�I4&mf4-�yZj� @j��?�#��8/����f���ZIU��d�_d��ؤ��WG�۴i�!�M4�~E/��� ��a�
�B��¸� 5�dO�X0�%%���~�҂��!�ǣ�-2�|��4�9�0���b��X������o*�; @�~��7;�0cƌ`ĈU@� D}>�A�a&�(���u ԦTĵ	["P`����D<A\}�
�y����x�M�<����"6������q���UEȰI��u�I<�P�	
ӳ��CR]�Mv�|�����w�S^[RRR�+͂Y�&�b1F}��|������tp�?�.$0D���MA�O� �����\��$�G<�`f��'yn�5����u�H>��5P�8Ym���C� H�`���I�Ha��c��I�q fΜY�]X�f<��>���Ft!�HZu�ån�{�Ə�w��+D��昼ޣ�I�Խ�-��s��	X�S΋�Lۜl�'�OF�<>��"e0����W�C�m���W�J|�c���� `���F�%��n�CIk r�s#4U�u!u��R��`�%�+���/���R[�p��^-�,�9�����g� �sF�������aC�5(!�Q�H	 Fk{��I7���Coa+N�ט��Y& �q�|'�x(B4�t��M�J1��$)��KR[��͒9s��{�;��{  >�Cb�X�s'�n��Ga b� �%���qS���&<���upj�S �0��yFK�����Y8@�x+d7ׇP��q̈4 �� $��ɼ�%A�C�:�fTC��e��xWx�Aռ�UBM�\Mr!-I|�~0�}��'�j��r@�qh�g���f��A*5�3i��
�T�Mf�'ϧX+Ɏ��n�&hfr��g|6fd�� �/�����J����Sو��+M'�E�n"��1�&��֙�յ2VځӇ��`���M+'�v�@%%o[�ע���2I���p=�����Bei�$H��I�p������65����kCe��N�Uf�:	�^��MA�s����Q,���t]���B��*(�*v�)�,�0��*�N�^"\�%��D�v}I�2[�����A�]��5MSP-��RH�ˇ��U�w� �|gը-�T��N��*�Y_g|���>��c��ϩ$c�:]8��A ���51/�*���6)�3\^���EW�>^&�"�GN3U%Ve|\9=�>�:��kW��F�z`����IH�)h��~����I
�;i#���:�h1줁��Q�>�Wee�.�_�D�g����n����-��O[ j�ɺJJ�'MP�4���|o
��^�4�S����Q ��(��ɨ����"igp%ͅ@�t������j�o��$D�:�A �=C|*T�ad��gMD�� I�<�����3��:�ƿ�3g��:F�]��e��8Bȣ�P[/$��(�,�*4R��~�
�G3h#�պZY5s����+���(��ko�$��K�K2b|�,p_�������P����Y��H��|*���s��w���{}�"Mb2b�3��&q�̈́Y?��U]��U0H����M���}�a��r����Gwq���9�����٠�dU����>+t�'�b�B�O�E����:$�gb����7h߾���~_�V�t�O�`��Pp�Q�	�� ��s\�h+k�}�w�O��q� 1Z���pl���1�b}�jY�ȏ#���&`�}\A�r #�w���"���4|��1�P�8 I}����	4߳�-双.b�:�扫RW5�!%�Z��^���\� �P�~��w��j��i� ��ԩS����r�'����HRP�dK��f��J�|�BS]���	w�g���G���`Θ���e����Bei/D�h�
��m۶�K�U��E����>��;�^7�"�~ppg$'���*�����͘�5����Wݱ�)A����3�RR(������ɳ��>�hai�.]��c�^ �Z��\��-'�����'�4����h��)��p��x>f0 ����.E>��!�8N��{�k��Y
 P ��o.��eA�>}�''��-��oɘ�(VH�.j�h<ҡ�aJm�?��*#K��V��U��;T����=�P���1l$ 9@x���w1�Td��v�^L�NgX���i6r���9��|�M)-�/�A�� �4����6��*=��f���o�s��U��E�h�D����f��8����]�Q��#!�=�f�9rȇtT�ֹ��;�)r~�j�*U�D"\��u��U�,�+�s�O#���̐���_�#Fi{@����Ӑ�����m)�@�gw9��j _�@{ ��J�yJ�T�ϊ[�#k� %���q<SS�<[���Z|<}OE�
*��w�A�w�a��bg|�cl]���0W9:(��|����Cs
��нT���$������񽰴�C܏�	@�����p�Ӕ��D�P>�pedw	��S�������uh��O��;�[���$��`Ӏ��鐐4�c�6����y�W9I��hZ�x���w��\ep��(�j�W$Z�髦 m�O��U�Ǎ1����
��u�U�o�U��N�IS���x����^Kj�1T��]�S��)fdx	��>W�$�  �ر4�������7�����W�7��k��4���2�m
EZdgP��򎠴#�>bk��:x�� wP0ri�(#"f�a踇v$ݜ��k���|�@Rⴺ��:aGF��xS��*B�HYc���#3͚�꒞:�ON�v>`�m���u�3�4O���j��`�ʸ���5	Px݊�(Җ��'U�� ��TO^��	�S�fkUH��k�Rl�T���q�(�
�QI�b�>��H�[��y�c(���cS�9>O��a��t�dxp��/���F���u�@E��!y������WI�P�S���!�]�P�و?zo������=D퐊�$(�V�5�f+C��)6fKDI=$�����ZQ���i�:�?�]峲v 4��߯iA �@M����G�+hw%yk>'"T�O�txJ�\�1�������q�[o�̛7�]+�ܾ���et���3���z\�#�<�%T�c�h���5d��{5�ϮKPV@�ҿ~ϵH���S��0�Ƣ��[�nݩw��ʱ�4R#��\[�'� �%I3}05|`$�}����'�����ȢE��X�d�b�����^mڴ�}�!��7}���{�9�s}� �d�r�!�����7��z��I$�m�������7�xՐ!CF0�K���" ��0؃�5(�D�A:�@�(ݻw��g��s~��i��g<Xh`�8x��ۯ���q;��l'��F3��!�{.��?�s�9#�����_t��w�yǝ^^�^z�)��0iҤ�v��ѣGW�$W/���IYb��`؋l����6�!V6��	'������
C=��;��E6x{L�0a������_�� �~��6m��A�F0F�D����C�?�x$�O=���;v,~�7*=L�
 � ���h���B���(�
{�&퀄t̞={��ar�'v5L�۷w ]t�E��~��!=z��RRRRWrZ�@F�������kݔ�+������ߵkנ\L�����U�+*�&� �j׮]йsg'9�[+yO�)9A)T���q��-fZv�M7=A-}`�F���v}����m�nSLAH��X�@�����~�JZȈ�Q��f^p�_Y�$:w@PY���/�믿>0�v9���̢Nj��B#RM� ��I����:�(W���3�Ğ�&@��϶{����\Px`&!آ��u�̹����o�!�&fC=�0�`�����u��&�`n0Q-�x饗�hw��ͥ]h�,�?餓�Pq�00� ��Yj���Z���y�Fx���Ql�ǝ��{�]w]��%�' �{�`�x���8R��@���GUl�=��=d[�ar)�ax`�ݶ���ٖ���"fR#ý�q�#Q;�4��D�;n�8�R�����s++��S ��?qO�d�����ĉ+F��(� ��C*��n'�<3�Zy_֖f��gy���0��\��D@��!M?����Ix)�cz{�M�ш�Z�P�5��j�^%��.(��D��4�ei�"a<��/t���>���&9�F9@0�G�� ᚰ������/w ����(f�ۻ���O�ҨQ��~����&��8��Ӄ�����q�{�΍��<���Nv��� <�2����R�+2����xa�%l�B��4���R\`���gt�����|�1V	�(1jqA�^$�gR��U�����K.�i�<�#^�ڄ�ô7��gϞ[xЍb¸]�*}B�a����:����<�Lg�Ѓ��CPS�A�~�W���fG;N#�j��`���D�NbDX���h(��Հ@z»��7�	'1i/�8FصH$�M
`y&�g߾}�d��ƣOz���B2�=�X��ɓ36@n5�ؐy\� 4Q8��Y�f���� �H�G�� ��[�<��W����(�{0�JOy)���u��ô��|�&U#f��}�k��r����� �c��#�<2y���gϙ3g	jRg�����n�m����>��.��Ӫ";0�w�=�d,¼�D��uv�ٓ�&!�L��t;v� $0���S%�D���r�k$4ʠ�t�*�:ˈc�]:>\I.U�7�?�^E��}"�;����l!.���O<�R��n�i<���3�~���� -̀w�ǆ�����JeUftc	#�?�i��iR�.�5�����Lz�M��و��`<+�$��d��*���|�V���ɋi�/z�V��(�/�ÓO���I���iչ�D�b�Is��>��Y4N:�̾����90<�'��i]t�8���<���ۉ1�qJ��ngaï�D�`E}/<b5]�f��R6I?01�cƌ��.�6�ŵ���Q�Ǡ��EƧ��2�T8�K�T�X�*��{P�ǀ#Eg��Z�`��Tr�	�\���ۅ�'�.0T�	q��ۀ����j�4@��9[imv�{l �4j�Q8D�0݋w��a �@J���G���g�q�Ku �C�U���x��;�&Mr���Q�.��.rȇ�0)DY+��D��s.-�g+rV%%� d+���q�\�H�?�3σ ls��@�zZ�A�\K1[)�\���0GF{�9WH���͖��ҨNiPM�&D�@@����@��0Ɠ�ɖ0Du�N��N�YaybR�xY�آ��D���ǹ������M�:E~�h���
���~�(F-I�p����� �q���)�:'w�~`�,&�`"��-��{H����k��*!d��Ue�Zp	Y?�gkR#��«c�Z�� �ֵI���"�FBRޙ�њ�C��(�J6u���$ �������o�Q��)�LF�E�������&-�٨��$b�/���]�}��E9�7��իK�֭��=����M�6�>��L�Z�t�I��}�֬Y�м�'�>�Poq�Yg���~������ꁕ+W~����Z�h�;���|�$�y{o�}�6�ѽ������~����XB��������w6P֔���΢��I$�m۶�`��]��m�y�����&}��mk`��{me�Sbjh(�:�d��,9��ka���;�z�UW�%A)B}��\j�� �ر�X��ǒ&�j��ך��qէ�vZF�`Tt�-�4�ٳ�R�j�c`T�NS'�`?Pe`���Nc�� 1��Z?��W_ml������W܋�A�ٍm�<�m@�}�Lm=8N�7�xc�5�n�쇮C%e��v�����j`XO�TH�Q= F���R`TH�Q= F���R`TH�Q= F���R`TH�Q= F��m)�����Tk��Zo�Ϧ1�k���_�mbPk���k�ƍE�5ڪ��Aiii���.kE���>+
���R�ImU�����mT�hK���V�ZUԲeKݫ��E�������:�+،�??JD��    IEND�B`�PK
     ^�[��
�G2  G2  /   images/ee130f24-d674-430f-bd58-6b2b8a983a65.png�PNG

   IHDR   �  �   ��l�  iCCPICC Profile  x����JA��h���Ha�E�4JL!�b���F�h�;�l�l��_�t�v��70�`� XX�"h�]dҤ���q8�ܹPzBTn�(δ�v��޹��AIN._�	�%���"������S%�S���q��*\�
n
n�ʒL�ذ>���h��9V�6���hx���l��iW���6).��"2���oX��^p�	�ޭW�B���gw���ϭ���` _�ك�X��[Ăٜ|6����!�8G�(v�Z4�c���??�42D   	pHYs       O%��  0�IDATx��}k�\U��>�/s�Ln	I����@
P�>QQK}��ReQZoQXbY����?,(H�@��2�(#
(ނ���Lb.H&�dfz��9��s��==�I�$�{?5�9}�t����Zk��N>I��*���ax�����ix�����ix�����ix�����ix�����ix�����ix�����ix�����ix�����ix�����ix�����ix�GA�Ap;1��0�!���A���d���́un�LȆ|T�T('3�O�� �Q�l�*������|>?��'-<��@��j��x�@JD���SdT��ao�Z(x@d�a��װ�X��'�5�l�g��K�M!���=��8��:)���Eq�"��@�����r�X$���/��JB�����_}�޽8r�Hoo/6��رc�����iӦM�>}޼y,8��S;::l��d��?�8Jbj04��/��K�bKG�}}۶m���+xm){zzT��i��¶�i�J\*;t�H[[ז�� ����E��Y�f֬Y�-P}}����	�3�r�G��VD��@�V���?�x___������������Rl9���^޼Y�~�x�Š��l�*�koo%�R	D����O��d�iӡ������?�s��Zz{K��R���p G:���"~e����à����G��	`4����u�F(1x�3�� 1G��[���8)�����
�/[@'��)Q�&2����ݻ_{�g�}�`������1~�¹��`0 X�#��4���WV��g�yꩧ��`�����^! ���O?mΩ��v��٧p�Ǒ�����{���������v�x�	� :�14��ß���~��g���R�⸂�A�}�P�=��1=xܥ���Y��СC�֭������-[�쬳Κ3g�"��C�A0�fΚ�Rh}�[��_��#H�رcӦM�&H D���ꪫ.���D�zK};\ ����H@�.�5 ��_���O@�A@�!d̜9�c�z�� �ň�#7���Ge��|0dx��޶h�"��^zi�֭�-�
�;,�c�=�}��+��?��9��p��3�|�,2��$��ݥ�N�+����_=�k������/�h��t���B����|�E�W�נܐ"z,oo�>}�����r�ƍ�lْ1��������#=�]wF�޾޶�6D2��Ml���oF���B���w�<CX	� ��n]�ԓy=��y����K�~��ٳ/^��g����+8�����O}�S�r�Q.�)vNN��Q����������>��v����)��+��B<�kl���@�0�%�o��S �9�>S��@�y�s��p/ C�4����'�_}gG'�M�-WCP_8G?���H�����<�0P��Ї>�t�Re9�C6��)���`a'�)�]'	�馛��~�>.Bp���|��n��Q�h�!T+7s���98 ���{���i�a~�{�����^�|9�*����_I�/�/V3��v��Rj� �%.��DN��v��:��~���ׯ��7���<����_~���\�L0����я���K����Z{^����k>x��g�],K�%8�2����0�~�m��aq ���~@k���(�?��C�/���+Wb��)"�����|{;�����=��������p�f͜�G� _��3�F*�<Ll�!H���M�Fi=�=�=��;:��L�~�#y�� ��*$� ,�����/	ՠQ�9�A u���sρ ��e˖]xᅱJ�+v�+���38����]6�
T��9�KR����/~�p��1}�c3�_s�e(�����gT&`uA*>�8n����~=S�R��?�|���5���~�����V��:C���T�>�Hq���qEU���a�?�S�=�\X~GWW>ڶm��e˳SAü?����`ӦMo��� ۸�p�paZ��yc`�,�����$�AV#D��JN�Q o;;;/���͛7S  y�=���>��t3��~)�QY��J�>�{�'�4L��:��T��0�ZD�8���X�e�C(��� ���o��D��R�fȖj09��;؁?\�����u�ց�R_^����s�=�) �$"�0���~)��dx��@C v2����|k�����u�n���8�.\�o׮]3gN��lܸqŊ-�<+�xv���̴(c���J}���?h���oy�[��-s�v-Mf�S�b1<J�9Ɩ�%'�׬Y�c�~k���eg�y�0�{�h��O�U���;�����{����g�}�\!��HO:k���`{C~Z���aaO�{����ӥg.��h�8	|�7v�U�I6�ˏ�������^悂\XM�d�N�mշi�`o�k0`T6��Pi;N�b7�|�v���Y����G��5k%��d}�i�	�;�b��A�L�_OȮZ�����oh��$�,m�r��@�W�cW����/��T�S`$���p� ��Yl���qQ`��������g��Lb'��|�0����p`�=�0X6` p��՗Ԫ]�%K�l6�����_޺r�B��tبꊦ���F���l�x�t����$�)w~����FX��QÛ�	 b�'��P��"���:k���tS����4Q69Y�"�����v���1�s��T*�\��Vgg��4����G�Ď���p���ۖ,����1��3Ācl@.Y�BS�˗�&���ߘ�쫀ۊ�8}9�8�2�TgIs:�R��Ǥ��y�c��2b��1e�K�.��7�����Z�Q�~㆘���3ft̙3'�Z4��~��f���#��eDN��B��h�~^�Ν;/�x�\α���WY��M�G�����)�H��0q��`�ގE�ǫ�C��eĝ��(D��*.�E���vuA��/v����������:w�\q�8�DZ�z5��n0�b8� I����{�B}��U801�,
���{f�.��i�W�*��x���E0�d����_�����?$�DL��H��\��ÕϘ1��=�����p�~�u��gA�~ʢ|�����ht@�Cv�娷�t�i�>������2�:��J5��Ov��ѣG�	�pCO9�I�v���7Z�U:����A��p۶m�X�fR~i�H�޴��F�P�r��oi��u�ReZ[�~�{�����9� _���Gi�X���V��O�w�\��/���տI"���@��[�m��s�RY��q�8���Q�P�/���&�I)��cC���2i�Nϝ��̜9�>�*T��O�,�LҾ,� �	�L��o�{��"
��$���)%�[���ӧ���_f|\hZ���ڲd�j����Z3���k��7���H/�6������ф]{d�ĤPv�~����_�-MKFLd�j:��ҊM��|.���_�W
��~�E۶�?º��.��O��F��d{d��'���՜t�Ѵ�+��H�Z�0��/�'(�9��?
�"V�u����y�p�8u�jl�Fn�8��}9��H����4�7��U����f�>�,u6 �L�J$�@U�1�8p�2�t���b�y�5�I���t���!���dA"%F�h3����gϞiӦ;v����;B]�y��H+�Qg���V:O����6 ��5��C����}=�4W(Rh���V�[93A�����!���_ŕ��v�ʕ8��vغ�e|��k�������>��|!���Z\te@��d�a�=���z�Ov�Zs#�[�Յ�x�+�U ����&Ko{d���$���Y�����U���V�
m���B��D�$����zB�P�ع�~�y��w����s江��� �-ݲ��7o�����+>�+����l̞=�k��9��BJ��]s�`�W(��5�QG4-�#C�t ��72AVRzL�Vn=��i t�G�����>�͌;:�CobG8�
���)%�!�yT�W�O�O�&��Z�s�N!O�;�h������9pv��rxj�dVE�W���-[�Wn)1��<@D�.х�k׮ůM��Ԧ>������}�G$"�˥
F���+����Y�3W*��M�g􅠌�>?`��3P�O13/m]��_�z5�=��?���ĬY� +��OTLpC)�����?��#�g�]���� )��XQ4�����?v�I�B�E�r)[��������z��с@�+�WSt$�IЈdo�&��/k2q��_�5Gz�+I�`H�A�W����`zmK�.���_�K��oذ�ںu���E��u��dMAbM�3�Ef�:��鯁��$��+!�o}�93I�	�E��@Ѫ�Kcz�)~���.~�W�t�}"MS� �֜(�0�fƆ_�߻~�}������ 7+������qka��{`�/��2��%�0�7n���f>|����m���Vg�j�*�wa�`4;�ٴ�n��Tch�t�U��"�%�� W��σ�(�ӕu�oQMz2 ��>}&$ N>��0�O����+v�V��7����@rG���F��?$�<���B��F� �B�o���d��=�Ie�}�1���ۣR����џC��G��G|�W�)�i����<Ԛ)[���1�u��ݻw��m۶�%�mO����ˏ��m�8G�p �5�O���&��@w�%�ǃup��ƌ�
===q���q���2ڟ��%Ն���_��7��! ���ƫ-v��tХ�^
��7�۳g$C�(�ސ���Wj?�L&pU�^a�	]�6X/5�Q25^��Qρ����&n�ܹs���BOVd�~�)�aď����X���+	�,Y·�����2���^{"�#��XeހX��g=�UTݽ�'8t�睝�b����ѣ�7+�C�������^7�Ҧ�~��:4�*el�fV)�*�]n��������������� *4$`�R��>�������K���y��q�>k�99Ĝ�ư���|>D2T3H5Yi���%o9~c��Z �z��Qܓ.4��6M��)�PP�z��`�_��<R]��QF�.2,����Z����� L�L��ijryK� ��N*KeG��o}�w ���ݮ���Ħ��rM,'�ͻD�؀�T����0�+=���wsZma şu7 �S�5����p��5��?�#:��	�&��[���^Sa:��:*��z���4�.��k"د�IT����YA��B�;��c�L�}w�����کhX��+uʂ����I����I�:��=b�Ta����A3ӯ�
�p#�|N��\�'[Mn�&��d�w��7|�M^��0�*de#�ʤ�Π��a��㸠C2z�����$轝�S�b#e�H�㬓������N%	�|�B>$a>��w1����[sz�o��?�X�e��q�������5I���pD%Y�(�?����N�H�Ѷu��r��$k�Z3����]I�L�%q$�$��wِ�c��r.��
2�F���;/{B�?-��=�T�&aD;�z�|.�ւ	s�i %+	i���gI�Y����(��c��QC�}O++�U�KiF%������ȚeD����x�8k"m�#���8����cg����q� {��*(��I���k'pq���>��~�@41��Q6%hKgC��	Q,�qYt�����ӧO�[>^Oe�z�d�{F�5.ܷɖ'�J�(�N��uCv��F�z�8�|�	�SN���r�p�����)S���r)[KbOWWW�=ׇK�j��y���ICu�w�6 ���b��/����>f�([�p'���@�Ԥ�i闌�L�g|�y�m�C͢Mfu�^���ts=����p0�5�-�}���P�+-���L���-7��k5��KMK��G���ᖝ�lϫ��ِą�Z8{|O8�{\�e�f0]�i�.N⨬�N"���DhhZ�e��$X����ӛD1��d����.����н�u�5_���u�΁=�e3�d%r\���Jɀ Rf��6{mZ�%�"ʹ�f	f+���W�?��?���6>&KX�������p�\J�'Pd��(<>{�R>�7-�7nܲe��U���������f�V�B^b-.�̅i�>틙�]���?��<\\	��ٳ����g���n��A�id��xѴ�'��-qֶ�Z��!NXf�C,ӱ����ۇ���\&��;����:���a!�@`c�޽,O���&v����j��γ�]��_]^i�i�o��QA�>�1+�J�ac���_��L�-[�rq��vbgoZ��9�1�===�YZ�4��;�6-�S�*�U��'f8Tc=�!G����篲�"���	�G�ǔN��MH?U�ăZ��ڵkW�X��������U6KE��N���>���C+�xCPɀ�;o޼{���{��ǓnB�	� ��&�}����"z�jP�l����	�-z�����_�қ�j@��8Ѵ���["c��=�]�aW�(���3=R׏s��u��+	�v������Ѵ�[Y���7(r��/K s�3�����UU�u�TuD���0�+�����~65 Amम�>&Pb_�<RT��.�ִ�����R<O9��{�`��hW�׶�x����$0Y��%z�H���نjhZ�Y<#����������0o���������"�Ӕ�R1;��tj'����1MK�L�2�kO��Z��/Auc�α�^ՙh�W5i�z�MH�P+�Rr���M�|㡱�R`f����\Qd%�8p�������èf�B~3�J7��;��Q,r�U*�z�KI1ٔ�u3��.8�߄�I�l
�򫯾*K�y8O̡�Lꨰ��0�ʒ�/L�M��|eC� T��Z�~I��O���4汴R��'(=R(Ԝ}h6�k�jr�{�������*�L�2���P�=]Q���q�ѻت2)�@:�Y;M��Vq�i%�;���tmh�#Tp�<U1'r�,AT!�����Ý(�5�2^4�6���b�Y��磹r���w�?k���L����%cåS��N]P�Y����$���v�g�덲Uq� ��<�mG�RuX�/�P�Yy�_j����Q�I�d��f�l�t�� �+q�6�]�V��=�6�#�3���թ�>r
Q���43� C�˒.� �x$2�dX�L((ɞ"3��L�9����7�v�vѢE�$D�����H�#¿�������>5���8���̝��b^��r%>|���/�,�*egg�+��ޟfe˖-G��Ē�,
>��ӧO�cHk�i�&��Yt=R�x��̀ɐ�V4G��C�T�.�{i��v�i�f͒��&��'P�=����]�i����\k�R(�y��sNK�%�] ({���'���r�%���� }6�q����l}[[���_p���σY�C���+۶mS֢>�8�h��|A�k.�Eq�σ��@T_�K?��2cG��/�M�L�ó�T��N�N"���)#LQ,����?�י�͘ %�'V��f�zHI���djҸ�.K���'�?S��|._���XX,Y�y�W&ƽjb���i��e^�!=qk�%������hJ@ud�@\��J���˭a�,�I�t�"ƫ�)����¨a�{�gtg�/F��=�&B���?�k�U"��J��X�;���.5-�������)��.��d�K�918G�Ӹ�V�H�N5��dT% j�:��ړ��*���
@r|K*O68M�(�X�I��5S�j ������x�ka3�S1A�Ӆ�?��KR;;�;y�%���L��4��CRb�h��N��8��
J��ޢ����|�J�	#��r�p���l&�9���yc1�	��ݥ�F���{�'9j�{5�b[��Tܮ��"�vtL׸�Ę���Dy8O����;O����;O����;鷗�$يk�$\��C��w�~���w�~���w�~���w�~���w�~���w�~���w�~��"�,q�F������~�����U�U>�~���w�~���w�~G��~��?O��Џ8R�!�6�_�����z`�0@��rNf���)���w�~��鯢f��i̟4w%���Q�y��~���w|6���ֆ�3�|��$�aN��c~3��q3�����{�݅��]�����է�M����?$���.���>`���4<���k������r�~���w|�����?��o����)�*<�N���4<�N���4<�N���4<�UԄ��=����{x�]�o����w�~���w�~��"��ŏ��K������{<�N���4<�N���4<�N���4<�N���4<�N���4<�N���4<�N���4\��E��\.��|>�F�I�H�����4<�N���4<�N���4<�N���4<�N���4<�N�A�ck���39�����D��j^8H�G�~���w��*jV�g��U���4<�N���4�?�6̟���`;ѯz?��&��� �Ux�����ix�k!�s��c=���w������{x�]������;?�;O�А���|s����;��N#1��� O���c����;�\N�^��;�8���7 5!~s�����y��;O����;O����;O����;��,~E�}��W�$\��C��w�~���w�~���w�~��4����k��M�_��{�#|\�,H� 	��>�i�=<�N���4ܤ�p��7`�~��u_��G%�\�~���w�}�0��;�g9�Q
���|�\�����zd�N��2���_ƹpF�皛J��3���f�A�7�E��J]=R��Z.�q�3��0xX�����f��A�]e+Ǔ�S�9�q�mͣ�����5��@u|��"�ĸ��Lp����i���0D�i���.(��d]�_hfA��z�i��! 0"1���0Zd{����"5Yp�� ��^A�Uc�χ�N�q\�������2�4��u��;�2�*'�C(����aY�I�{�!]<����4����ݯ{�'M,�����p���@�L����P���s��[!C�sc}���C���z�7u�2~�נ�  �Ũ��9��J��|���c����b��c'�x�Tjoo3z]��¤jP��WӦM��O��/�E��5��h�~-����\����Z[[1����ޖ��Ę�0a�G�}R�C�ayǪf�6��}���g���A�'��ʘ��D�>^���N�s�?�w�~���\��-���ة���i3��k��\)��zagg���&�я[�q�r���A�`����`���G�:�sa}��=�t5r����[P�-m�Y�: 74S�1҃l�Z���m�P��Rv�s�ɬĒ�/.	F�h8G?�2FV�=�|H�t{�?1�B�P�/�9CKp�.�g�2���9���xׯ���!�����������>����?W]uU9*�[�1ō��ݯ��k������~( /�>�Ae'�я�Kj���z�؆�3�B4���JT�[��F\�h63?�ׯ��GDO?z�o��a������~Vr|*c��XwǴJ@}Om�.;_��{��KC��(�c���:#�9���3�~�;���o��?��꫙q��6m�2A�I��3Զ��c:���;�o/^�s�Nq&�{� ��_a�����{����mlI-��L'�{P���h��wގ;�2��_�@�9�
��je��	�����DH��]���o~�7�\s��͛q �O�����s��v3���*���t-Ѡ�n�0�4�a���?�0��+�|�W��d���_������6�=*�6�;/՝9>� D�]]]�-��+��.�%�
�&MB̩��Y?�Yp !`������3{Á���6<�N�-��G�u>8�W59)?�\��gl����)�h�`V��8˺u��:���o��رc�9��$忪�p�~:zR���V�v����� �:���+_�Joo����q6���D��w�}�M7�I�s����L��2� -��u��)�t�_U&�I9z���L"SǙ�W��.6�\�����~�Q����G/2r�6(|R	���3ē��/�-=�l��=z"8����U�1����Y��5�Hd�����JEs�����e�������}�p���~�L��#���Jϼ/�>6������R^�`�wsd�~ժ������=s	����v�?����[������c��ٳW��/3i]F���7��?#l��[�w�o)�@�9�?�r[S��+V� �a]��_O('	k)�,��>�L<���!`JUYv���@Y�+�g�-��:�����k�N$s�����|� 2G9�N\��{V����9�%��PM����ѣG;:;1���]d�r���%;��d����`�wÆ�Jnx��$LH�O}��W6�$ �f���N��v��"s���&�d�Z���%�=���k ��g�Y�l���8��+�HE(�`������ā�i͸��/L5��/��,��!_�7�����~��~�M���G����y�O?��;���믿�[����m��aaz����8G���q��2��ۇ~q�O<q�&���	��H�~�c�`ƌ0�^z�}��n݊�����;���C=D�#��Xs�N<�C�xr� uѢE/����ŋ���w�}뭷b? �>ew�E��Z��?4��G�{����QBh�W�X������n���z����O��!�0�3g�|�������|��L,rv2{�O��^*��l���'�|�;��o�;���}�f�|>F'��s����������?]y��-󐆅��7�Y�l��R��񙹀�(���R�s98��5M׼0��J%0���!z���ܹ�?��O=���,����5��h���L�_c-6������.gr�֗_~yoo�s�=���}�^���W_���OS�X�ş:�����R�����s��ƿ�
&q�A��Y�w�%����?_�d	~�g�ٹs'"��1�,]�N<��@�2I֚�6�)z�H)sH\���+J�g���s���[�ʉ%���V�8��NJI����n.��o}�[���W�nkk��B�O���?
��b�ӟs��w��^�ˊ�z�7�޽{Μ9�1�;gΜ��/��9���d�s��\~�i{���O.���_������D
�V����;���?lKC�O�(�<��'/�\0���|�_\�nݮ]������7~�����`������d��A<�?���0��\3��1���������S�}B��dE M���cM&�=p/�`���?
`̟z꩟���>� �*~��W�v�mk֬I�H'�)O�( ����w�|�IeR�x�����W�Z�~�>��n�1��q�������w�sÆ�]v�~��g��;� �l��'O�( �W]u�g>���x�կ~���o��oܸqǎ��ϧ �٧�(��P�ի�3�?�x��_��׾�5��v�ܾp�[� )��('6A'>�;vx�G�;&�����}��� v��\n*Ox�G=c�sܸ����,Xp�Ek�D��x���<�i�I���ѓ��_���y����R�ٶ��۲~t���?
��� ���s�=f�~��?�yy���	�Z�+O�X����	ܛo��y��n����,~.���SS��Q ��C���/��o�g�}����%�� ��]�����?<��?��A0�����gj��\�[��R�􏎽{�~��� ���w�ҥK�U�����i�&ĵ�^�Z�Y�f�u�]����X�u�u��x�p	��A�����t��{y��~��M�6q}֡C�0
(S҃���k���$|�\���?4Č3�٬�"�����ejA�I�SK<�)�������җ���wܐT�T��)O��Q`�=Qn�9}���)����)O
�9ۇ���'C�=kYe嚰|��Ğ<���h�4���5*����h��0�{��5���Q���q?@�|�2�A!�~]S��5����]cH0�.��a��rn���j[�|K�/�ݒ۱WkL�:O��w�~���w�~���w�~���w�~���w�~���w�~���w�~���w�~���w�~���w�~���w�~���w�~���w�~���w�~���w�~���w�ŪX����    IEND�B`�PK
     ^�[��Vt�  �  /   images/193bec7f-e59d-4bcf-b15c-6ea8617b7acc.png�PNG

   IHDR   d   �   f�  iCCPICC Profile  x����JA��h���Ha�E�4JL!�b���F�h�;�l�l��_�t�v��70�`� XX�"h�]dҤ���q8�ܹPzBTn�(δ�v��޹��AIN._�	�%���"������S%�S���q��*\�
n
n�ʒL�ذ>���h��9V�6���hx���l��iW���6).��"2���oX��^p�	�ޭW�B���gw���ϭ���` _�ك�X��[Ăٜ|6����!�8G�(v�Z4�c���??�42D   	pHYs       O%��  wIDATx��mp՚��鞙L&��T���hI��+[�Uֺ���X~�uK�`���eQV��Ze�����eE�J���\��%1yK $f23�g�s��3=��LOs���k===���<�9�������W��a��˅|X.��r!���\ȇ�B>,�a��˅|X.��r!��[��:Wʷ�p���3���`�&�q�2.HFw�3�����v��$W��f\���,���>v���9�� ,��hb�����}}Wz{oq�#�D"�uu3gά�������b$˼�nt�s3��r�Ŏ�|�׳g�z�L�H&����o`3���������s�6��@`�ig�#ß�7�ԅ�}9�:Ւ�Ա��9r���H$#���Ph���e��������������o\;z����.\�bżysa7�ih���B)7Y�Rzn<�˽W������kJKK�,l]��:sfciiy0�I�6�Z*>�-�uu���/����c�=�H�#T�&35����K�B��������f���@QQѼy�V�\���7��S��Q-
�Dj��5k֊G9y��ѿ��歡���^��Ժ�`���|�r��YE�ѝ�|388�W�^�|��p��(|�L\A�-�	�\�|������cnsӁ���	�Y�_�>
����E�nY�P�x��W_}uch(RY�O�[[[�S#e��fܕ�񤝽�\�����aÆ={��8q�$����~�o �������s��m�S��������[rD�`��4D��A��0�F	�/��y10�u�֥R)h���pǊGf�?��[,<��e�5k�,Z���8`VV	��L�r�Rؾ�y�A�2k5� k׮��b===?��CsssC]�ɷ5�/�`�˗/C��Xi鲥hk@E�4N��蛸(���O�R��af�Fjg?�Ayy��?�c��(��3��wryE��e��}b�r����7oVVV>��=�I�Ȓ��!�d�tW�����5c�P�;ŕ&�˖-;p���ӝ�D[�5C/��j$g޲�v�|�K�������V__o%ʚ���)��]f-gjD~�\��.]����S�[�?��S��&$�6.-<,��/&���={vxx�����1�X~\��r\_cW4��2�s㪮��oɒ������uuu�}�PxX�&	HS�d*�����3t^%o�O�hl���EMG�,쏑��ڎ�	r�h��2[�.�/<,"x�e]��;�w��ϟ� 0�p�
P�T1s~e�]��	^�jn���ʊ*�;;;!#Z��aB<��s����`MM]CC=ra��C؞���Leat������pSS4C�����p{���E��@�x��uX������*�	^ <�Xs���ͬ}�M��D^�B��.�XJe�I&�1�ۆ���h��nRN�%`i��n�<�O��555���c1��--����E�w�q��ymm�G.� �ƕ�Z�ʶ/\�� �`0TYY5�/��(�!)(�v���0�!ZVh��,��bU��ga*ᑧ؀�R�+~�遞�
g=����=Bu-,��Ԓg"�r4�׬�������4kK�	&�H�u4�`�yղ�����B�-c0%�B���Ǟ�i�O�(~�$�{!4�����6v(<,́qYDb��b�,�����r��BL*��4�p��+�B6�,,���a�v�a=IgK������9��OD%��۾���hw@��i/X�@��)	�N�=z��S����3JKJg4΀�)�t��)�:V�^��� v�8b�Q^�`n���%���}	C�!�.��\���=�@0i ��������Ԃ8��o��t����L{{{II��p�����p[��.��Q��%68�D��n���c��p\T�40���3�緈1A��湮s���@@|y��ՁɌ�Gz��&	��@�$r'̙�.�V�(�rӄ`bz>&J�*x�d2��o�F�ݶ{b`J@P��pQxΜ9��B�=z��E�T����,.&~n��0����w��麆���+..RK�.�{<u�x:t��{��qY���w`9��"lrU���멦����%��i0����,\�0����={����n#=aV���f84+��0.����`:ﻬ�R�ַD�V]]�d� ��ϝ;������^�T��b4��UG�o�d���c}}Ckk+����.\��FaYn��b�9�4j��%2#фt]wzh 7cƌ��&�)�藄�T0$� ��4�I!f�h�?B���%#������������p�����s��X�*�^��UC�Ar��Xpf+�d���!"oll@V�Gx�4
��$4�e%�%rH6 �@����d*�I�3��/�P�4%87xu����/ dm	�2{���وm�4�0��C�@����s�B��X��8�Ɂ��=��e���d�V�u�ET�:�ǵ@`���L��K�#IIeDR�x����c�ی��2Yj�i����0
�E+]c�k�`�f��MVc��f�bdK)HTL	ȣ)*�Lu1)�xF����}5���q|:/gs�DRF�^�g���v�K�c'�!�V�k�]`'��Y}�И�'ٮ0w)K����:�[��=�'�&F̾�@V�Y�'��r��Bqqq�$RTβ�I�	{(**

ɯȪC�ZxX��bhBpZZZ
qf2�*)+]02��"����V�!���W�IO�H�Z���Q?ӊũ�6�@%�d�V(gsK���GZ..;�ݤ?C��e�!�Q1H����+t|D�Z |��%��i�Yz��+�������C�=�N���AL�U�u�ʕh4
�����|�:;�@�I/�^��੏�z(�U�eJ�]�
c���Ç�m(Z�lY�ް���^��o�>9����uwfy{��4�8�<�����s���vRSS�Hn�������������)��1�E�"��������vX��I��X���;��;xx����g��W��<��0�0j�!3c.u�q��`"|x�ĉ�{��ҫ,2��B0UYY)W::xk�����9wj@')��V֐b�S�
�b��Y���Ҝɢ���'8y�?�ǅSQ\��JǦl��̉�M��t���ߒx�Z���ЁdY�	/e�v�lW:��cZJ�P��;M���ÂfQ���������u��S.��8',~��<CG�S8w��(f�hX��aW�D�_$�o�����pZ���Ǚ(�Q>�C�"���^��`������o����[������2�u/VXN�	�4ayC��Y��kbز�\�x1���Pм��;�L¡����d?T�q��_z����H$���������X����
���Tb֌�UUU���-�p1�Ƒ@'8ڂ��Ú5k�ƍe��m41�?;�����7�g�����*�������C�ayNo�ڵ�gςs�'��������c�=�`�|���ݵk�a�;:V��S�$�13�ƫ���Ж��2�iP��^!�'���f�K��\��|?z@N���7=�C��mw�ibF�����Je�l�%�I��u�� �!Y���s͸��[�M�YEXR���� �������9DJiX�i�
c�4N"r'aQJ�lwE*�r�:ɱ;��2�H}Z�����s��5?[*��G8�1gW�i%�4,W���ߘ`.�4,Y�q�Er7�4,��ŋ=H㸧�._���W��a��˅��eו��R���a��˅|X.��r!���\ȇ�B>,R�]V�
�z=K)�%w�a��+W�>˅��Yx厬�3-�	��h��R����H
�B�X)+-J���BT����U�Q���^�^�i�G��B��!�$� ��nGp�d����i�T��P��B�K)��r�K4����|���-扪C�1���]ɇ�B>,� ,���b~Y9w�ޝ|X.�*,��)K�2C�����|X.��r!���\ȇ�B>,�a��r�ԩ#��r�,)2��)Ua))���\ȇ�B>,R���J��M�O������x/6�P� ,T�ݥ}˚D��.%��Re��&�����*�Ld|6(W�����P7nWD�²��\�]��레�y�
�'���i�>�\E��ʮ�DuX���ݙ?�/w���ɇ���᳘n��q�+��\HYX���R�^E7�-�`Y�&*J9X*ˇ�B>,R�6e��54=���9ʦ�n#*�r�cL�Ai5a9�?cݸG	)K<��5O>�IE�v�G|�w��"�s/�6�%6�	vy<�Z=X��9����'ڞ�C�wQ����Oz���6��B1X|�5�pZ]ג�c�ďjϪv���rޚ|�����%��#�J%a�0�n���r����0poT�?y*Ǧ,��`(���>/��H��8�vqg�ʢ��Qǣ�*++V�Z����rxj���|�mmm�VX�/���'�TC�iq�@��I��U��Vv�m���!<}*�6���I>�>�x�ل���y�?���F�s�ҥ�;w�����=_WW��|��SVL�{�����^�3g�4�<�m�,��ֶm��x㍾��`0�ēOΨoH1��kD�S!��իW_}��h4�z�j�5��S��ӧOwtt;v��͛�4�\L��q6Y@����z'�I9X``V���<����@>;!Ԋi5�j�֭�V�ڿ��O-X�ᵪ���;���h�eD۷oܰa�OEj�B��7��`��[�>���M�6͟?ކ�a�8�<[9X1f�[�j�o:�O����_}�̙#G��ٳ�~$��А���Ղ%�m���/f�C���m�]�#�LA��74����f���ֶ�������"y��(��5�"���É&��bƌ�?�a%dKH����y��6l�gh}��|��-[����N�aQ���B�jll.**2�4��FuB*p�L��8��[�������ZB�T�Q�'�ٵkW2�,
��}�"I����6��1+n ����=��3��t*іZ����	��b2S��tfK���hgg�ŋ�|~�apv�#���`��������u>�Xv�8S���+W֯_��e0�͛7���N:��)W�Ղ���8~�UVV���[`A���|��K/-^����==�%�y:^?&�̬��x����;��$iY�r$�5���>}��>;|����GK�<q�Αҩ��R���r��zң5V-�/C���G�B�|01���q�*o3S�Sp��
ك���_�?�x��_|�O��e�hoo7����2Ny	V*���	�� �c�¨�z↓'O�?`aaz�3��MKK�z�6�[X�d��޽{�޽���۷oojjj��i��<��9��c��vww��'�n�������O�4��,�󴱘�,6mڴq�F�!,++#�����u/����/�n���֭[��+����ʒ8�ٳg���,�m۶C�ݺu���ܲe&4�6�t'y�����ʎ9��������URRb�%��<���^z��H$"��у,��my�U ��ٳ/��W���A�Ǉ��ߓ��X8����~���_&�Yj�D^�z��=���C��Q����/��}��������/���0}yV__��͛a��f �v�-��7�� ,4�D"�f͚��ax�:�=`Y��!�, ����~��\���"���]���fE��B(�+k�=�g`Q��&��
j/�"�Ä���ʇ�B>,�a��˅|X.��r!���\ȇ�B>,�a��˅|X.��r!���\����~ϣck    IEND�B`�PK
     ^�[	��} } /   images/bbfae99c-8036-4c5e-89fd-a87441410720.png�PNG

   IHDR  �  �   ��ߊ   gAMA  ���a    cHRM  z&  ��  �   ��  u0  �`  :�  p��Q<   bKGD      �C�   	pHYs     ��   tIME�#Պ�  � IDATx���{�m[���Ƙs����8��GսU���袍�i�4��A�("�q�6'9�Dq��E�HEVd��HX�d���&�Н��g=��n�}����ךs��?Ɯs����{����f�J������k�5�x��p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8��}�𵂪 ʳwQʄRZ����k��{�Lǁ�%O�h	*T�J�`011@��#�QD
*B)�@ FI�"4"L�Db4��L[�>T	
4AU0����11��*��J���N�L� ��m��l@�(`\m.@aW��7W�G�|������%���<�Ç?���p8��h��@K�J���s�H��K���EFi��_j��R�kh�,A	P@	`   �jQb���!f(PA�U{�B8��W? � �FE}E��z�T�0b��P�t�>��1�yPr�P)[��7���I�����>P�+��T�hT ��ۻL���J��ui� ��5%Nd?#��z�vH
U�w�[��}��rV)R�""�%' ��f�v�U!�bs�!lJ���x�/.��Σ�~�S�����G����7 xD������%b~�]  A�=��~l�,!	"bz���
�*�E �
$S�
t�Nb�Z�L�WaEM����DՀ�Ĭ
�h�AU���!7�(���?��˯���1(��a��%�۽�����]���$���}i8���U�5�ժ��T�[T�GE�C-�J��eC�����	d�VE�RM��F���dQ�liO~M�?'0�w^d^�b�Op�x<��L�$����3x� T"��q���/@%B���w���w��ڄ����k��3o������k�q����:Eӯӳ� e�n|�Z��	U�M"�7h�Yr��((W���� D��@U�����y��䟽��� �6� ���X��D%"H�T�(�R��0+���	|KLO�x��8L����m.��>��m.@aa�]�%����P��/  �Sm/�J��eM�7h.�SD��J�$_+t�RM��
 ن^X�f��@�aJ��QS�t��k��纽o>c8y�l�BqĻx<������{MH��sF����J�v�������U�v�+��K�������]^\��^��������ԟ��|�^�/�-�p����; t�0�>]=����_.���FD�[%���P�)	R
b�K)PUÀq� ̦���2���_�+t�;������2{��W�~N�D�DF���k��q( �fB8�g���90��2�d�����q��o}a�X	�@�>�G�ᗍ�VU����n�./��'�����/%�n���Z�K*%��Pɦ�T d�ά��H��Du�Z�9��yeӕ�����}N�]�v�W-�~��;?��c|���	s)(���QJA�fB�C`036�`6q��F��,��j�@�.�q�}�_o��v�y�~���g��W~Ƌ��Ǉ��q�`ڿ�_�o~��-������<�Β�o�o��V�|����D2��\!���!F\]_#�(Q�W�Y7ƽ˧3]oqǕ�\`S���"ZM"�� J�jTM1+���y����M`��P���ϙ�gƟ��~�Ke�q�1^\!��1��,���;�������/b�]�����U��HI�Z2 ��"	���`^yۨ�j���l&��mH:��@��l�
^P]���u�{	@��9��s��{<��s�7��.���L@��i��%c��؍6���1b�<b�#��E�0�+l����U�_�������b|�_n���7^^���, "���~����g~�G_�2��W����O�����%�v��7�i��|8n��[���R@*��PJC��`�!9���E��^z�U쮯�(��RU����� p� )�z�5���5ki_2����&�5���5�Ye.1WEO�����9
�'����e~������3������1ݾ��}�������o����!����?��9�.��T��9���I�"')�
�慢�B{�g�Z{�^IU��mt�Y�8��ieٮ����$��qԮ�0Q���.~a�9|*���ÌL���9�((#cF�P��BDĆFly����.�<`Ѐ�p��Kx��|}��[����/�~���T�O@)������W�������~�ǿ��y��/a�yʘ��b�]���o�Ͼ��2r�~��p��3,����4�P) ./v�$ bLsƓ�^z��x�ʫ��
� "���ӅA<�t����<���])U��kH��Wy��P��]��� �r��G��C�U�/J?�!�(��#���,o�M���#���#��p}�����u�П���|�G�|���������e��_�|+��*�Z��BHU��(t�ͧg}	yK���*3
�U](y%@hM߯��@���a�y��`��s����N_�8�@IAA���`F �!�b�
��1�6<"P t�J@���p�勏��W�`xTv���8?I<��ƿ�H���4��.��C   �7��+��4�i�p�x�xx<D
�:�ߖ�߭i��A��8o���� � �3��Md�H���#��9g�./����g�N	�^~��������Č@=Q�z�I��;:_���LV6�^�l��H���_׾6	�<vQ q�P��@���Y���q�� �o�D7x�c����@�P���/�*��A_�����폐����_�^�����Ayz�� � �J�h�V���c��S�w�Vν~I5!�)t�j�/%]š� 뤸��P���x=@B"��%Ct��@Q2��j�H1�Z��JI#2fd8!% `@�� 	!d��������F��:��?����R/�t�{C�o���6=~��v��o�~�qw����AU�RP��Bd�p�:s)�ó�?V4��9�ߍi���p��·m)�I��{H:@JB �%�'H�(iF>�Q�H4(�>�@cA�	�M7�i��;()D �%oz����q�9t�:W�dg�o�;��#����u��I�%�X�a���|����(�߮y�#!���@o}���8~vs���[_�N
��~$�}�y��޲,� �Q*��9�%��kXӀ2A҄��4�z�P���oYY����aJ�E�*��j_�*�cYXk�PN��l-(/4;��.�S*7����S�����	��IZ
� H�H�.� K-��"
5�d0�6؅+\�x�W.���xix	�0"`Ѡa��4���g���e��2���x��p����-!����n��K�u����9��3 �����͗���o�*2��O�\~_��o���O�i��N��y"�3Ho�Z 2!�#JN`"��9!��r�0�nn )!��8D��r��E@q���5~�۰���FFV3#R0Yc���Q�.DW��ޛĉ�~��P3	j��6��*s{ͪ���O�u�y�T�����UM�0(�X
�'a:��C�i�ݏ�{|����Ȓp������/	_W��/}�!l>���(�Z��-��D'@Dg�(D$��I�\��%�-h�Ӿ_|�U�v7Zy��1o��B������״}��;��"�ܴMȋ�iT�b B$�j�,�JBT�[J�A�X���B� �غ �H ��`@)B�6(��3o��4��4 �	�kL�c�O��g���8�0��s�Ͱ�~i������w1lw��t-����@��m�$�9���M<|囯5��۫W?6�~�j���K���U��n�O!�-�dYfhI�r��-E��	I,^.9!oq�y
��0n�u����3�4�c��ͣ�-bܘ�#��a�K�J��J�S���$�U�ng9��޳�R_T�9�h�EƂ�@�����OՒ�J�I9D����)㯕0��D�ߺ�<�����~������������O|�ʬ����O�ւ�Z��!�㿡e�(�)G�r�j2[���T�<s��qن�R�T;�Ψ*t���F��9��z�Z&'銢jT�4*���-���9��ւ�Y�]D@PD
�H%�&����Q�VC��H*�b�#Ka�]"�Lϰ��pF��~ʀ(
�y�&��M��7s���Y���t��1�� ~!����g_�t�3�C ¸�Ї��43�3���/�ٳ=��
WWeh���u0����#��̀�rP@b-}�j%A���BH�L@mX����D���Iָ���Z�X�K���jZ����1�}��p�b��`@IJ�A��AT0� Ί�2f�vD���q����Q��0E�t�c���
����v���}����;�y�%��j`���A����o��I_�"��>z=ݾ��*�E�'E��Z�5D8���h�C��	�@��|DIGS� H.ȹ@0�	ДQ�#�t � C���05���uw��"_? �&[T$K||�7�ӄ@������u�{��KoΏ9\����%/D��=����f_tN��;EJ�֛R7J_#�@uF)�e��{�O�����~����~�w~�w�����V���u��o��|���W�|��K�H���"G�L�2�lJ�%ͫn��1F��Ϊ
��w�yL��M����E)��z�ž6^O�:��׾�aU �Z"@�lB��;��,O�@����z!�$(J��ށ ���l���p0R�Ť���3bQ\L��-�����A� ��RB�v������5���������3S��8��"z�oso!�o�?�O?���q(1��%��f�tv"�w��T�Բk�a � J�s�a�q���	L#�iF�G�M3�:Z2r���<�������}��ʟ���G�q���D��2LE��FG�b�c`��B���L��	, )�M��`bb��Y��I ��H�tr��7�>½�
�����_R�U�Fji����P��
U"����V!�K��R]
E� n�b#��:�Ah�t�����p!P �����^������ 8>y��h
n�S� xh+�Q
�60C�~a�.�J�s�JB��g�o��}�f�g��]4b��� )�����/�9^
�Hy@�!��H�q���7��oW�߂r|]U^*%_�f�P�W�Vb�%��@�y�e>"�(ǣy���-e���'@b��%c:� D�4�e����!�@nn��gL9B9X)Z) ��oN��%�T��G�ÛR&��!��Xe�$��nғ�A+��.R�m�e���Ξ-�K��%�i3 c)lT�D@��H��)�''�o.����nz���O��#���a_+|���f-�a�0o����5_)�R�Ũ'�H-+SA˃T]�oQ�a���g�8M�X�jU�X�6ֹ-���s��2�kѩ
Z)�wR��G�؅["D�Ь(�0A� 6A�(g(B��g��#B�dU*`Q����)^C�
�hA��43��A�!��A�^�^"���{�BxF����D�%����ox� �q����ՌF��� r�0��N����N3�W��z���y `_��"����.
D>����d�"ø9��IidC�qP�AJ� �1�C��n�	1��R؍X�S�4A ��(TsE��*7�\5s���C��L꒮oZP�7�7T�/IAbJ]�i*UΩ�Y�(DETUE��Q��q��THJ	�E��,Y@9�EU���PJ�&*��"���T�\��-�˂�-Ƃq,�~�_�9�B�R����٫Z��*���l��r�^�3=��C�<�������`�hH�޽P�E�#��HyՇy��\i�;���9�ΐ־Y�'ת
J� �(%[-�<��#��M	�fS�R ()4%d�ӌ4O��0#猔R�P#�b�R��0����f�� sg8툩9�M�5[���Kύ& ���K�{}��$ԭ����ԍ�ƪ��ηváv�_=]��p�b� �d�I�oU%��w�VDE�n��2��ܼ�i\����zV��*�ӻ�'{�q�M���/i�sH�G(gh��V�V2���>���@��L�QSƴl�N�t^~��۷}JQ{]/1��Q�&�v���^N� ���M^[�f��FR�`l8��#v�E�2CHl�Q��I�d���I�zp�`��DDe	 &&��Tn��u�b@s���\KE2�L��  03�Ja$#��� V�P�C��8&���(4�(QS&��L���U���(I��+���� ����k����v
�<;��T�i�����a���2���(��r�BsR��H�L��HDL̡*_��i`Bd!��͆i�/]1^}i
�U�K��q�u�V�����û��|Խ�6L+MD$���Ｔ}L_՚����R/n�7o+%Y6qVe) e0���([�DDC9BDTPP�([P�P	[`���P���VG��"�%�HI��R��Ǵ���V�!T�T�c֜7�������Z�̌�{5Z�v<UHUI�����V��b��*K� RX�0����b^}�P�*��g��S�Ħ�i�q	e>�oQ��d�Ϥ-�Rl��������
���cJ8���%��ْ�b b4�:M{H� �S�-iM�@cS���YS���3=]<4e�L��&��7��D]Q�2<f-��w�n.�~��G5�,"�mb%S� ����Cx5���k���n��4r�x��O��Z����~��C\~��雟�m�������'PI֛Xg@��=��F"�j��V��w~" O��~M��S4����z�}�,���歯�f͆��ڇ�d��fc5/{TƆ��BϬPeX�2��Q�D��p���� +#h@�!����!?E. �ƂѕD���huRTC��� �"�z��`G�� ��o�����Z�&�Qz�w��y��CUf�<eL���O�xrTd,�X2B����$b�:
�xf�<�3{�D*}K1�ĀAB���0!h��̀a�������D!�����жt����M޻��o�[}����F�,��'����ͻć��ď*A���Rt�-^V��$��%b�p��[HA<a�`� ���tܢ�K��щ�P��-!l*1AF��lbM����l�=Y���
{?�x�=Y��k�
h1o��Ĭυ4�C(�"E���T{OT�ԩf])tj��u{#I���|����) �֬�~��j��|D"R��<�8���8D���M�l"B$��ʼ� ��7S�(�i>�϶լ^�n�ﲹ�l]���{��*���F��* �:�et�볰<+2O�b芚���ĕ(�Q	Py���P��}������ȳ�O��)<x�[�aǇV��~����@���4���n��*�
��5Ͻy�B���4��*���{����z73׍ghq������K������������E1[���
2�P��  ���
��b,�F:� E�Rz�A+0p(��\`��y
(]Yk5����C#��jV��!�׃V�q���#�g*w�ξ(�/pW�j���1�$I @�3n�7�`�@����D�;WDP�@T0�	%[�b)&l+8�b76RT�	��U�h�\�	~'��}����N�25�6��~��	Z�"�	"]��l�
�{��)T��!@��t��i��#Xf��`�
@cy��4@C��-hs�v�n�p�{_�U=4�¼(��8�2�M�[S�XN?�m�(s�5	x.�5>�3��j�I�z�K���O�,=f�{���'��=@5�\�]q�P�#����JNV]R�0��V�V�3BP�t�����^_B&3��R�t ������ߢ��h��t%��2�O����T��^/�k �Tma��0�����?{�J�KM�CϷ��r�若�E�� ������������'���{�	�|�Sx��oy�g���R��޾�gሇ�UM���K:��G�̖"�f�Ve^�~	��!7�l�n[��%�ӂ�-J����ן�)z�+��O7�J�wLZ{Rj���5�X���ʜ �2�H
��N
S�\@�M�Aњ�7Ȥ"(�}ge5�t�@��r�1�A��`�8T��湒V:��}�*�%j�ΐ�E���m�"H���:��`�ύjڽ���D[̀�� �#O�,RD�l1gV�@��5r.�sF))���!R�e�0�-."a`���UjhדX�3���=(*x>V���-LY��u�� ��=�u4� pT&�NвM7
SX��0���vL3(O�<�'j���J�TD  <��:o �%�`�ov ���^rZ�U��Ր�5-mMZ�ЪL�p��Mq��g�n��[Bz��֥��m�h͏��_H}F�Xy�-��׽�O�}��)��a��$	��L77fP��
�����mă�s��2w�v�n��Q&���	6�U�!��o�N�Jj�u5��]�r���5[��ht�ʘj\���AlD���^�Q�2�~�*��~`�L3�j�Q���`���69W`{��$
�����O�G�+����`��e|X�S�
���ޔ|�'$�T�<hIF�kF��PG��r�V�V�̓v.+ֶ�Im���'V���wS�k�ܳ[�u�z�<��/[�]ey�)��ԪI�l���w&�v�@m��d0g(�*��%����6�%P�Q����4`�r�$3����л���ٵ��^&*�W�*ШUi��P�,lM�����Oj��w��(W�kJc�͆ ���Cf�"(U�81B��� �\��{�V0P�Zl��-×a��|Ļ���u��
H��O��T�C��]�rQ�͋�=����v��(��b�.�`���.��9�ƺrD��L��Ϫ	(
� �	�� %�����T "0,��T�2�)��!� V�._�� ���M�	b��GX6�+��:ٻ��5m�*��Z7�6���S�|��β(������h�Z={ċqQ=z�RKK�2��,Dl}�I��,N���9�!0(0r��b��#f�-V"I���`I��7�f���ۍ�<�?`:$�3dN����z��
�:٫��{�����5��x�M�wơ1w"+�[��`�G�����\�3���}4̌��OU�#֌�z�a	J�������9=���G���'�����q��gq�!m@�S�7��T���%����%�XӒ�e��l-=�]����+���f�����j��$��Ic�٬R:�컀&+D�F�¼��,����*�C5Fd@i�DA����2�b�'�f5+�Փ-( R$�FիoP��(2�5��Q��/#c/��2n�G�A���vo����Rf�;2\@� ���l�r�@�Ӣś����O�\ʲ2wj���k=1�B�l@R0b�u��	9<�f(P�le�2Z�p$F(&���d����Lur�Ֆ�R��
�12�����x0(X'�&�-���.���[����J	P�o�Jm�tU�띪�ꋵQz��-g�R�N_Dd���	:�V#���Wg��
��`L�,IrU�TD���*
���n!�-�b��PF 5�����B���O#�-�e	^�@lFT���<'�6N�5׵Z�ֈ��贌����3�L�Z�ZmHͣ�&�+����o�
o��vT((�e!OG�)a�8B�`�7�W�����O�<��֔��|�s�LG��"6q�V�K����YyY�nJ����^��:��*p���T���85�~�4�3�<�ET_������J *5�*˥�v3���k�$9�/!��O����ç�K/�>T
}z�H��'�|�Ki>|���:!�)	��lJڒF�4�Tzh���Bk1�"[�R��tE�uO��V+�����oS�M6,}�[}d}��x��
��!PH=�k%�����(��`�)�X��>6�	!��MHP��D	3� �z�,G� ݮ����,c�f-�|q�5�u*���m�cB��5���+/H� �������Ѽ��x-$R�9�T���9�Br�� 8��ԗ	`A���
)3�
���2z��@�R���RlT-�R0� S��`?r��y�]>�k���ݵߴ=q�e6�Z���<�~��{j��mˡV���Ȧ�+���6*����D���̥� %�L�3�c�j�V��?GS�f`�	 {!*��C@k¤�A��^I2&��0)jߘ�%le�w2�K�C<�<볳ؿ���[;�K<[����V���.��*!��m+��Y0�*aD
D[WHE)���h��!"�3?~�9M�\I�a`!������./���/DH�1����iF�%3�焠-n^�U(��Da��O7_Ջ���׶6'������ڴ��pL��idJ��.o��oK�]�����M��`�Ř��>��9zB� ��o�7_��v����[��/�>����Q誊��/!�Ã��͟+����<�J2�\l�o+�`�D¢Z�E� 5~��$�d�F�-�k�}+v]�D7VX2�W^�J�T����i{�	�槣�!U2�bk��Z'��`�[v��kw�~�%2� n�>�{�8ҌIf$(PM�#�f0pD�4� &�����܎$t��Q^)iՓ�5������Z�t�i�a=�R�P.��	�2$)����<!���JѶ��1FcD@�hID)�T��"P��{�Rޥ*-�K�=�z������(�^�VN��BJ�F�<�u��'5�AD�O���[�q[y{FEP������PB������ws�fԁ��B$���0K56YH� P��8��1�8�ᵕAB�~i��s^���^'���w��DO�ZU��_�.��B^����!��?tf�����0*~=DJ%�>���Ŝ��[�yBN	77Oq�&�֫���k��/�q��BDPR��`���'����'8�(s��4M� ��j�����@M�yW������BS��o���3�(���Bn����\������nșaѪs �_Z��%�ތ\�1�������O��;�����]|v�o5�&|(����������9������<�ђ[R�1b��%�Y\1KY-~�g�7ũ?���@��y��Q�%�ף�(zvh���3!��n�;�@�����7b�線�F���J�Lv�"@z�0{�v@Ĕe��$�P�g5�V"w(3&9b�	%�`W�}��j�����#@JFN�QJ�`��P��r �լ����h�"�(�F�׷�>k��F��Z%�2 �)f��~5\��@�i&���y�R�#�1 F�u����"�!�keA�sQ�T�Ů?FFL� �ϧ�q'˵�H盡��]��8`�ce���4�e��1&K�9��
϶΀e��ʘ��a�:im�|ʼP�T��R7��{U�x ��h� T�ʆ�5T�/D@f�<IP	�o�������c)��%~�i�n�/K��C��nG�V`(j������k�gM�=�S���I�Z:o�v�TK�<"BQ��������equ��d�>}�y*H�#R�8�v�ǓgO��l0������)%��<�\
�	����Gf��%l���7u�,,�%�ô$�َ'9K�@�r����:�җ�3Q��6�h5Z�:;-����)z�LY�u�2]�r=� ��2�������Q��|y���ǃ�+>,����"����]|�o��S����<}ea6��՚��I
�-~���Xr1�doz~d�z���������j-a�3�W��X��L�L��1*#��e���5_]p��aM�5�A{G&�L`����Q2a�#2f�Z
 B�� ;$��5�02�x��F��x����0F�U����W��r�%	���,KZ�v���߮�sk�c	�F�.��j��S�-	�Z7S��pn}�T�JAI�s.AB�H� �(IPf+�4`�ڎA�%F����m��J�5o�HWR��{�'�����e�`�t��S^�g���JʟP��fL'��d��`��ք�Z��e��["�P5LXZ�F��s�X�n{E������9ke+��u�v�1��Q^+�sZ:A��.9�gJ�mW��E�����]��wj���/	5����p���J�Q����R�tx�iNl//��G^�~������ FJO�1��r��a�ʌ�xDJ	Zex�)�sO}���a]���㥯�k�;"��Ȩ��\^c��V��$����z�S�W����I�z�^#3$��6B���?���/������}��O��cߌ>p��������7�v�돤��?U���J:�%�D!ɐ�{2��R��s��r�~��K&o#�j�2 �z-6Ӕ���9x�ڼ�x�h���z�,����|�r-be(b����q,��2n�P��0}��S��j�6���%aFƬ3�L�2c���l�!�pG�C�ц�l ��xF�R���,�z!��OX])t�$����x�,�{_�V��1w�J�
��� �1a@ҌP
B�Z��X )c.Y3rJ��>�gD�F���E)+R*`hQ�ڞ�4�*������S_���5��[h�y��������0+����e"��Q�EiA��iz�7&2Mlg�$��0��T#+t���Ĭ-�ь 5�Ό.!K�5�l�n.�����ڪ�_)�x�ٛAsj ��v��
���F��I�7���W�S_��("]�o���9\Փ�����QE�d�C q@*�<g�R.8'l6#�FpQ�qy}��|�u���x�����}�� �i�8L38D[����	i^�,����3��s���Qp�F��$c���oxnI���J�\�{j5�:+��8n=1L�����\�e ��L	N��
I>�����0=}��}o���x�o��T���%���ax���(��G�|T&�Z��6�	4Z��K?�Lړ��k��S�Qd�� K���Xka���Xv�2?��Kq��/8��V�t��=ʿ%C�6��"F���������ѫޓ�:oAT�X�M��Fւ$3�L]�[�j��z�bε�e�vW���8>@���:C9#�Yp�����S6���εRWt��}�L��n��lb1�w `�)،f�
��֖��c{(KY�KR��X�%�eA��`�C�hQxUkKlԟ�n�?m��
��;Վr���G-�g�hԽ�h�*���! %,^��>FcQ�GҌ[��5-�7�޲��%���q�8�&�ڡ�@�Pڹm
�Ң���[(Gc+Dj��T���E�:/����K�����װ��Y{R�H���3��(��#pzx{�W���2o�C7ԛ���3*�[�@ss@�qq�4g\]]���#���8N3�d#T_{�%�~�d)x��cd���T0�qs{���{�a
��rFN�ĠYd��lRks��t���8Y�;����K���:�������H#���ۺ�I�Z���~���B[�f	�"��A(vn�:m?rI b��t�^��/��>���;�>��ۿ|`
]U������_���{~����h>��2A$�g#����	�j<]!@� �Z��&&�-�D;�5i:��d�V�D�P������e��k���y�H�b:������;�[Љ
;�Ӈ:�KA1��0b[�Q��)����ژT�@�2*�n�aP����lY�(�R$HP䈩�"˄P�B	�C�Ad��$A�%=����!�xe�j�!<d�Bt���&a�1)���u��{+���E��qq���ŦTJ�BEj��"�pE�����焒	4bX:X��Ա�@$BΊTj�
� I	b`��`?�΄cV0�d=�j��P�h�0�e:��I��v% +ͣ�̖��R
��.���?ۗllPh	�U�	`LK)(Z :!ȡ6	1!�4����$"����JMk_]�F&k-j]�
��l����������4�����	����E�֑ �)YIT��ֹ'���ւ����v�m[v�,�Ѣc"]�-L�:�gevF~�>5�n�Y��+;��i�����w�l/����ݣ+l6�4�����f��^������	�b��<���,'�x8����r�m�{5M���#'
�}y���vΔ�q����L���g'���t9 �o�u]����C뫯'��Z~�U�؜�j�$��I~�������������߂����|�o�-�������=���I���t� 5���,Ѥ��-q2B�Y�u�A��ن�W]j��.�`��O(������W5��w�Z���|�$윾�Y��\� ���7}A���[�U-.W։)�M�b���,����f9X'�b���-CY��?:���@��:C���L��E��������� $�Z�o����,ٺ
�nNUa��ߝ%�����D�c�E���m$"d�q��fQ2�T�p HY�&�D"D��`���5z*�\�X7-����o=S<>�K대dzZ�*ζ:XNH�ԖF��=��c��Z9���a��\�Jw�)Ag��^"E! J1_�,fK����rWB����Lw��(�Evk76Hm?��[	(��a����e�`�|v�������a�Ӄ�&�E�5�Q��f��J. �}�j� h�H�S�f8�Q��q����z�-sga�Z�jkKZR��i\ (6�t6`ETPJF�'����#����a�-B���RJ��v��	2�9c�#a�ݠd`;��n�SB��)8��)M�P%�J�!�,,sKe��{�x>I�<Y�;G�����z���c��3���Fw�c/_���>
����:�	l���a.�24-�D"�%A�d��_���y�}+�>�<.}>0�>=~��똏��W��GJ:��Ɇ���#���T�]J��Z��5�^��K�.ٱ���ߟv�[���`
y�1�f�)�=v}rg_��(],����p
�u� m�.�bD`
��jrגd�(�H�ſ�P���EfZj�U�u���Z�EY��U�	a�#�	*���H�,�ea������DKM�Z���0Е!Ж��0�H(�\=j�GV@R��j�s�&��J�zܘ�$"g˼�LP@����Aр���@V�����L���18��ߺ�qCN�����CS>��;���@Kz����q��ǵ�U ���mF�V�3C�2їw_�Gv^�a}�hM;��Ty���"���d"Y�Bɦ���-=y���=�P��� ��"+O�5�i}�W�\=c�)�O�w�V���*I֝�t�m?\��f1�g��i��[_��&@5A���^�j� ˄i>b�#�`�MeZ.���߁����A�f3"��'X�RPJ�dWǨRs�Ob�f��f��}u�V�ק�)�ޟ��q�峽�����Ým��xr�r"_t]]�Ƽ
 *���=.�2�1���O�g���?|�����	�������UzH4g�o�B��$�w�:9M{)Z������dP9��E���U��Xj?������[��7�*rfMU���ݤ����sZ�Z2%���0%�Ɇ���&�B7Nl���i$��5��דs��SR˜O��:#�D��#����<�;ͳ5��d�&�N�������`j�nBAd�z��^/�s�B*�lXw[k�o����[���L�o�m��a� �%�Υ�Bd����T���U��CR׮������x��w��?���Q�]� �����s��vJe�X������֙��������J�+b�!��i��[+�:e��#v-���K^Rm���/�ql�^�:U�
ъ�4/{CZ��v����7BNAulks�AK|v	�-�	�>9�X��*��_���-�R\
3n��|#����)��A�@ ������vLs�������^sr��@���%��n�#�<M�ӌ� ��<�w��u��{KM}ϟ�����-���'��:z�*���V�ja=TÔ5�Xȥ�L�Kӌ m��@Hy�.�����|��o���>�m��'�s5�Z��+���m��_o�������_]�[HI`d�f����j����ZG�5;�ex/����<I����4�y1)�S\��� X�t3=�=i^�T�S+���,�co* fD�  �)b��V��h�,nZM�B��Ų�u� ��h%p�Ե� �p�������.j��[^i��*Beu�u`E�ʢ�O̵%[M�6/}I$�,N�K���B�;��R{����-�c[d��[+������S"�4|���#�\[̮"��;�t��[������?������$��0��.m?�?R2�5F�0��ތ%$cЪ"E����wژ����v��[��Z��z��+��y5"[0j=^�ʹ��\vHK<����-4�ʭA�'�����{=�=w�2p���i���-	�˂f�BK��?`�����
�,(*8LGp B`\^^ ���W^�v�E%<~�m�\����`��y��B����0�RrgS�ڷ�Y�b��������c0���g�wΤ.N���Z�ʥ��yYRs:Bw3��X�s�:��BbslFg")��ռ��o��o���o������k?��k��U��x>���%M�?O7����3�N��*(���-RȐ�@��̵��	�^�J/�ܵ�[��?>�b����+�6}�y��^�:n�ĈȨ��C��3O3í�zS�l� ˀ��	܇*�c��=%Q�
q%q�����-��X&�e�D�D��Źև�d4X��Xe|��D ���1ĥ�nsS�G��.����C-�8�d,��;�a�z)W{L�Q�	c�"r1ee��Z��h�t�0* �Y�S2�z���kAk�[�"YF<�g��E"��J���&,���������/��+�۶��B'�*��w  c7
�MR�#@�+t4���|)�Z�6��3.�	]_Ok'[g�3B���@\�z[�$�W+O\rmM���8Y�t��Pܺ2R�`�$���s󱭳�X��'�:�V�^-�g�>���������c%�|�*/8\�v�~� ���<ς)%�ĸ���؁'�����g��O{1c�6O�@a{�E�)'�4W�_��C�Z5rNo����؋��9�876ϙ���`w����l�K 3�E�V����$����R��UWC� (׮}���Q�ux�J�v�q��l/���n_�D'���B�����7��ø���i>��r�}%�#4Y	���敷6��(T4O�� n
�y|� �y��Y�Ve�R�W`�Cz�����5�� ,�Ks����l�1�����W2���X�dS�T[��hͺm��)�*���R�[Y��,�)��/��QɹR��h��z��&|c뭬�<J[(,Bz�G6���F;wA�9�VZ��m;��aE�v؍�0�=�f^�Q�1Ty��̵N�j[��yW  �lSڄ�����Ҟ�W�z%(��g�M4N=��/ܞ�#�t��m��z3��Q��5��S�}��Gh��"���޻��u���mQ`�z�5'$�RCkW�/� i�EW��]�=��]W���q�qzv��\�h1&{:�?�x��P#��7��|�|��[v�H�3�[~Ƹ����
yP�h�x�q������~}�5��?���/ �#^}p���#��<��^��ZA�5\rz�~�Ej���ߝ������P����R.w���@��3�)úGl7q����rv��kc�'
f�5�3�}T� %!���a�o�0�Dz�~��e�5S臧ORP��g���%~MI�������l�W�7��׺W�H��@��Z��N�u�,�RA����thZl�5����l���n�s����A�6V�Z�VJ{%,�W)� L�1�ujS���K�w�w��ʭ�����ɖo�;��PK��("�4�Ig3@�Y8KD�h-t#��m=�ﴇ�1���N)���)���Ӻb4*�F��V��J��Xp9L8@��c�
e�D��@�mp,�[IlP2PR3�IUPuN5��L3�d�T��($`�`+�w�����0B5Ygi����fw��oE�'��(�n�Q��P��3�����H#Ѯ��	j#F{�{�F;��]��(� /���L��Uᮜ��̴�s7Lq�����3��{�~qB�.�C��������j��ɯs/�u��G�!+����f�� ���BHHl@#A�`�[�������px���$�ݸA�{��b�C�#J�� l��jr�����ս�By����֖na@�y�����V��v�Ӭ��X[1�?YJӈ��p�����}��Xߤ��æ��bU�(/}Z�	P������c�~7��I��;�<��0��(<��>���|��5Q���u°�����u)�H�H������*����Zfh>2[-�m�:�eQ*�x�zB��E�%l�\����B�8�N�z�Խ�J*�+�2j��Qq�Sl[��*��6��D�m0{O��^��%~�5	.��` #x�R���Q�����:g�!����@T�"KX�?��Go�-�K��R�Ӟ-k�z��ۮ�e>].��ϻNAl��Vf�c7������B�,(��deL9)��W<+��	`%���[��U�)[׳8 � �8��J�t�h����Fo�z摟����t�N֮�&
W	E�=����Pq[Z��,K�0X�����ӸI� k����:�KkV��C����b{4��L{H:�,���،anSW^]���Ӕ岎��:�O��w�W�N��W�ѕ�������w� �_�aդ��$3���1[\<��������C�Y�%!�'�4c�8N�l���W��%A4��f�1s�5gِ�ߵQW}~}�Y�����%�@ݘ��,]1w&�Wj7��g��T�ڛX�j�3����Y��^e;�A*����*� +7���v�B�)�؆�گ���|��)��@��^y�o�q��%��5��o��<6��o�<���飒k�m��j׷�k���R'��X�;��V��إkTU�k�z��O�6�Z#�v�Z���i��}��鲉��>��%�K�����]���,�@K2�G�&\5���}f2�N�Ϙ�-s�T�ր���5���T D�jMD�D!��p�~w
�a�?|qo��{�j��Y��H�Q?���Fp10v0�i2Y��P̛��i
���y��6 �8@UpLq����p�/8f9)�i���%�4å��N�d���{��('��>�xH��H�ɇ(D`܁�(���6aX>�=}�gs�tc5	�v��s�d �$�#���k%p7��ޡ������<�O��\��rg/6#K�u-�2Al��-$�%�k��� :b��@�C��ѣGH�Ʃn�4l��KW`:������n/A���� F#�	�!C�#(
R��l�6|�:7AOBF����������٭r�� �JݘlFX1,�\�����������e�q`�`��T��7VT���h����*P��º��dk�L o?��~����Z���/��e�_<��
������݃������2���{h�!�6��%n��NK��gh��в��j	�Mi��ePb��\��i�ƾ^�u�d���4[B�	��%|��՜�����z]����k�n�[fk��V�<@1#�����(�ڶj��f

F��P{OB*1E��K��`���TP`�Ig���JR��
}�ث�Lt�+N�c��8�/����}5�̓�{	�:����� l��e�P�eEfE��."@jMgH��z%���ƪ.���v�EF�r�1)��8j�mfP�j�m�.}��#��X�-�Uo��;���:�?�A�ڞj� l�@�:?��,�5Ԩ�F)������ޒ�t.X��G��ZjY��[��^��<מּ��x��~�2�p��Wn�]3��\x�;�|�pژeG<x� ���%n���"l������C�f����K��n�!�	"2vW��!�"H���'dN���?S�11���0��+-gq���e�/���sMm]U̵��-9	�6/�tG�ܕw�k�P�=��Q�8��hg;�:TZ"rc�V%���ԉ����\�N�8|'��C��m�����l�^�없��B�g�0I�0>�L���H�o���x�2ی�>AMڈ�6��&ĕ�g=)���5����qIu%�Esr��k�[8�5��m�C�(��,�f=��]b�+�e��fP�JԖ����J���&�{9ࠊLmrي�V�uB����{�p���
��5�A�x��*�gɘ5�:�f8����X�_U��_.�"er�'���5w
�<gZ�S_k���F&l�a�@
�-KKQ�e�}�51�~����$dp����VZmÀY��8�Šh~Z��}�g����*��S��5�{���ݤ��"��q�\B�K����[-�b�-����PY���áf���
S�\2�B�%������?�~nD�oX�W*u���~��>C����j>G�{�'L�z��\X��J������D�,(qD^~����n��G�o�b�靈2=����T���C#�w[d��Y�g���m��3k�b�D�]������O����,���o!�u.��"�sQ�зOO�[Bx����)�X���S\�?�(�t���"��4B�� ��5F�Ǘ���7��}�ZP�_5�>��BJ���K8<��o,i����$iߕ���iu�r���k/�}k����uV�=	�	��X��!%SoJ6p�=X۸U(�,�T�=x�K���o_�����}Z��OX+ۯڶ�)��H�FU�����7$��r���y�@���Ba ���Y�� k��V!K�5#iFAO��I�{�}z�=كϫ�~�8����s]�ks�{��%[3cc L�T�Ú�D���ux�kB�5����\p��E�ՆZЀ��'2���:L��Lh���{���#i,Meb�yu��)����yU�H�-�hIo��b��kyd7.�g ��n%�������8�`�a883D��?/��ד�֊�q��z�מ\_Wk���dS��l�nF��>�C��@`_\�2n1l6@P� ��S��)��裯���o�`�nno1nF���ţ�݀I "�AD"�.���ah�0->��$�{�_�7� ��쒯�N�a��5��h7TE\�n�hj]	V��8yԶ��O��%(������%�K�@��&�|/1m~p����p��?��oc�|���ܗ���B ��c�� ��b��$y��(�CoʼNX+���1��&��zPa�g}��[�����"��,曶f&]!0�r&S�= S�ש`X��d������s]����ZJ�h���*��Uk+1����
BU��YۖZ��x֚1\=�6���X�u�9���O��{�a���4�}_hd�F�5,z�d����)��\yX�@dB�̢�@�Z�E,�Z`��52�PJ�V�!�E0e ��1�Y��S�SO�z� ��;��4�b��e�W��,���홝@�?�ٸϓz/���{T ��/B����?�`=�{�����sK�wu�"	$O 1Y�hZ�]E{�}���Yb��Q0gk�x��_��c�gk���nh�`�M�ٰfCjb�x����5�,	�c�2� 
�0"�$�#nC5�6dG2 	��&"F�$[��Z����dDkBk{�������p����z�¼(L'��u�Z���O�A���`H}_����'_�F3��'Y����%((BMn��Xcm➅�*�,5\l�ܯ1��Ç��t����돽�0ח���BWU��\\}�r�n��L��'���a+���^k2�f�t'J�@$V:C���VZ���,�'��j։F � ���0�u%���RK�L�4�ܼ�:I�Jg�0[BA���xemC�pk����}!V�$d9�G0cF�Q3�9"R 	!"`����j��q�mR�5�4'c=����6�cD�@(A�����&ݽ0s�Ծ�OA�o`Z��+V5�R4����Z����i糖}]�{u�g�"JA$j�����Y�P�9 Z]�%"�ጉ9�D;a�`�)����% ��CY��`T�� A��#H��~�U�6�	�V�mF��%��y ���3�z���r��� #�*tp�B��z� �<�(�V�&��P&�Z��ԉc rM�C#* �� ]���s�#{ُm���yl���r֦���L��lu���̩:�C���+�w�-���ۀ"�kC)1bă��\\���"4���1�@1�Z����e����K��x�Ÿ�8Z`�a�NV����8��3�pY2қ��
;��3��c=F��e���;�����`�:dy��B��UUPX��"�Vm/"�*�ɺ8�8�"A+%���t!՜$�Z�.3�$3q��C������O���ӗ~�����*
���~W�����=�]%�L:<�(y��r�^ �6 D{��� Wk�Q�2WS���|AM�iZ���[�7�
��8��h�!��$'��ڗR��A�4�
z�u8���\���r�%�ED�D���w��/h�}{r���D ͘e��r�Q2
8�0�e����5bĀ�G�&h<b�J@Q!��Y����g^��	E%��xe��ŗ	R�ss��	oX��~��PX�˒���c�e\k˺�V�96�U�����z(�,� jT��J�c%��b@!b ⚓`�������u�<Z��XM�"��"��rPeD(�3D�?=�w_H�%*�)�a��Kg�Seֽ��Y���������z�L�X��ژH	��^�P�Ӥ I�f@�w&K�$������Z�bN��źr5���^���0�:H�e��/��JB�7w�m��%����q�PhZj�@5 lPK�^c��lm	ow�QA����T��@�݈a�S����4^��� �(GP�QR@�;�������؎#<��	�no���*y���"jȤU�gW׫�yzX��	�ȩˡ&W��'x[����T��4�~I��Ő��˸Vjlom���.h�5"V��fК|�0Y*
�ĕ2���s5H �BTg�#�y�
�����r�����_�;���W\�����{x��s�����XJGk	ZR��[�[�c�;G��z�z��S�;H14���_8�R ��;�0��и��j�se�`od��^3����B�fL�ק���>�s�qO~L���(�tƭp[�أ`��ܺYu@��D	�D4��:�qd2CI�oy��b��TD�K��^V	'[��B��E+[)��z�p���K_���Z.D����] �!�ZՆ�T&�ƃZwd�gE2@���])g 38k�ôE��|���bh�s6���j]�kr't�}�֛�t�\���3�Z�J�`�� ,OČ�Z�ީ*To�NU�������Z޵<1õ4�.�y����~��>��A{ц��W�%�� ^ga!��Ujg��h���w`����Tp�zߵ�'x܀���K�p	�> o^�#�� (yh���ƈ;��+\\^�ٓ'�}�� ��K����MYS6��K'>c�*=}O2kk-ߜx�]v/����J�tMO�֏^k9�Z澨"��Кoo�**�(R�b���~�"�4!�J"�+��_�������S�W���WT��G�X�����9O�ߓ��<�!+���;ݞk��ORU�u��������2��շ�w�P� o.�����6h�(J��4C�h�1�t�f}��)���iC��{a�k�
^_�П�Da����(Gܔ=����q`%�8D� REfhIȚ��l�ݣM��楪��4%�C;�;UL9Cj�j�*],]�5���-1���Ig����)�JǞ��1^��� _'0�L��4�U�}e-H%#e���U)G˒堰��R�X��@#�1I�X��Z��R�ʓu���eo�m_����^+��{>�*�v���'B�y��������u�_3��R�Pb�W>�>	�<�F����a�6��ySpP� +��0ԻE�9�痽z����w��R���=I���ܫ��*����,�oz�Gݓ��e�}ev5.�1��L�#����+���a�h���T	2�@܀��|IO1�Y0O���x)���4(h,z�S�����yt槷���|�3���n��$Z���uiy5�_���NX��<|[1���;_�c��٠�Y�͗0���7��O���>���q�_1����SF�8���������f�t i2��+�d��9�ǘ$ϐ2e�t�tK��BO�@�h�vYy�-M
��+��)��#��5#�($g��OG��4�=lИ.4N�bP�^�꽓Y�}zS������ϧzn%�I�*�t­�q�G H<`�������b;4��	�6 rDd�Ԋ�l�e�pT�̄X�F$��5 �U��V�є����Z��J��=����B����C������.���w���B.�Bj�C��:u�fl���DB� .@V "
d��ÚpX����ө�J�4s�=�(���N���k�^����-9HWR���s�k[Ә��\�V(��a؀���J�Mj�j���Lm�*z,ݘ35j3XܝZ<^�|tB)�� ���л��y��e]Ob_��M��g�<ɰ31g�l�K��^}�RW�R;.y �2��'T
�9ˠ��_�x�1��'`�,Pw����Y&��$=��^B9c�#�e�=�JB:�.�V�Z�~v�C��qT��z_6gf����	�� z��I��>��UC�-����K�Ӛ'�T�75���H�U;(J���}�*4e>��0����DM����-�_����W�C߿��=x���������%�oAe����$��s��o�&�U�O�&��*o֚�~7��lr٩��#�C�\!lV�����!
P)�$h��!�(M}-�q�����z=,�)��qy�����zs����Տ��3-(:c�#�2#�BÀ�6���l�Y��1R �`3�À!Z����AҌY�L(�P 
F�ȴ�J�QB˕^c��~n} �IF�fdQ�tv�������U�]Z�)���Ϭ����j�DȢcғ[k�{3��%bY|��]�	<%F��5k�����QVh�R�GPb;�3�=�q�J?�<���kUg	�M�4�5�EkExn?�ӪҀB	d�(�:�������KfhJ�N�#k�ޛB��5]f�E!�*�v�5E�l_��l�������-�sf��8��טr�js����]�������,4�;P+�ۂ�0����q}C�a7� UwU����C[ JI��.��2c���&Y&��ץ5��2��ē>�,T�hw?�51�^�W��./a�u�%��yF�������-��@��Z(Hebdɛ��[������ H�Q�ï`
�V�^�?�O�=��)�_�B����8N{\���w���������&+��Q�g˾�t�J�ݞ34�2]��iյ�Y�ź��5����r31B��a�!l.��%4n!a Q��>���9� T9+d>��	����#\����k3�վ��ž]Ss��5�B�����[րH��k0('CDd�h#�`cgE��9?E){�F����2�L���Y�g��%wn�<�~�p����ڳo������[T����]^�b���]�;Yͧn�{�� � �ܛk����GjR����5-��W�ք�TC>R�q��ޠR�M��I�{��ŕ[� ��b���:ɮӎ�ۭQ���]�֞�B������?��Ѫ�[��t�0��V+�D����JR�&{N�l��➽��*O�>�}}/jvr���E�S����k٥%��=.�8�J�a��3�1���6�1 V�j��"(lL�ǫ���3��"Z7B�2mP;�Ae���sv��D�%gD&%����F������,t9����(xj�?�:t��e��慷�������M�6My��n{��1�Y����s��4MD��)���n�W���_�2�_�BWUdI@�1���y:��<��|�A��%X��kY��i�h��"ٲ�A�M�W)>���8n+{Yh��z��F4��<���ф	�fٚ`�Ƹ;h������o�iM����~����Yg`V�������"�!�k؁,V��\l/�9���`���l��aB� � �
�"b�V�"������_�Ji�j�D��/�a���]K�[ؖ�O:/�Y�%؅:*%��߮��b���9UO* !�1�����b�T���꺔�\2rQ�"(mR��b� ��L�G�����Ę���ݧ��#��#�sݱ2 @�HW��"�7Cc���<�P_*j�[hآ�����j]>���d�G{MO�%@�헚cCdm��(4[��h���P����FX]�6ñ�Uܹ��ʭ�n�2wd���㉫�iL��]�ڶ�&��!�(�J���lz7��IA��C �<nA�N�Bk������9��:T2(^��^EH�1�e�˴ǜ�eo3!<`��,��S�ķ��K�9u%V��ͳ���sWKN����������約7��-��>�X����{c�qҦ��\��������;_5�znB��f����V�,����VAdά�iSb��4�G����o�q���)�W I��V��e�ovWy������曧Q�[��7ŝk�j����(e�JsՄD+eVyh�����e�}�Mp�	���r��X�h#)����-��@ PV�6\�BW"ê�4�C^�U��v��-T�]���x�)9ka��D3ـ�Y
�*�H�L) "��1�כ+��Z�Y�(�ՃHFQgt� �8��8\#�g9���r�� �.h,V��8�u���������i��M��s�r�u��)�u��B�s���ֽ9=m��H՛�'f��1D(e#��"�6�Yj�W��fBa+��`i�f$)Hj�4	V�:q�3!�ơw�Y0���,�}X��߹�3%�ZW����YR���^�Zk_�uS}J�]�/��ј��Lа��B�(ı
��.(����~�����`D�Y�+26�(�Y�Hd�"A	��4�D�n�P�0��)�n0��n�>��A"X���X�qbʀk���3w�n�E�6",|��MX�e�i�����j1j)ku��Y�#t��$_�>���J�0@e5݂�����e�x�3G��̆IB�	Dl��f�۾0z`�נG�`Kl�:WC!U�W�pe7�$T�~&]��Y([މ�0�DK����ʊ��� �XS�
@3��ٝ����@ �t�[q��O�`X���B��d����������)�L)a��t��������r� �Ǐ�}��|�
}~�E�+��G������?7n���g��%[bKk�
IPI�bY�Z2T��shy��q�U��r��P�%��	}��Y���� �n�2o�e�j��P��נkņ���Uٮ�
��̛'Z�O(�R��;��VoN#v���K�-��H�1�#]C�D��4�0!)��_���+�m_B
�y�})O�*�*��vTkg�zl������2��̚Ʊ�&���)��J̖g�;_�xO�[���iĉ{���m"]^�ȇ���rm�	�m�������)@(� ��qS!LaNQFD0���ϋ�G﹧��:���Ӽ�j������`�7���E!ZZU�R'd������F]��~�c���X7�hQ��/˯�gY�+z���;m��RkힻS���J�8�ľ�Y�<�U�~lʼ��6j9��Q��֫�]�(Ue(G�q x@� �@���!8�`b���Ⱥ@��ҥ僄Z�Z�PH�t�q���3Ó�ȼU����=+�?���KP���u=4���Ժ$�M̀�Ϲ(��%���Ͱ.�i�槳]R���s�:�ψ
Y��]�"�&�3*6���QUf,g��p������Ӛn~��/�J��
}�]��K���_�y�w���7��3Hڃ�T��%���uQS/K+y�d��*%���%��[u��q����H�$7��uh{��(Ѿ3M�1� �q���Jn���@WnX�]��Z���(,_?�C[2C�J�Tj�oD���n_��h�<*
���K&<����.no'���\?|�_}#.����� '��|��6�*���v���=��(��4;���"��k��=�y_g����w~�_Ӄ�R��֫-{?hM>
dT;,���0ԟ�q����T�dƜ2b�՟�Q�(mV dUL	��!�J��w/�ݽ,E݇�����z�!uo�����ĝf֚�@�lUzS�zl�җ��t�^K3i[\�ACj65$ؠU�J�����ݙ�:�]IS�R��T��\���� �'o��f�/k~���)@��~�ү�gu2{��ٶ\�
��A�`D�&0���İ}�x�b[{T��=�pUv� ����GFjܾ��}]��F-�Z+\��x9�kw�m�5]��J�z;d{�b8Y�~�Mw*�a����re�Ȫ$�WA��q����J���n�递 &0��������2t������N�� ^��U3@�f���F�=@��䧆���Fn�z��O���|����R���q�3v����p��N�gߕ�O��(�M��*	A������ټ�R�I���.�G/�g4V�T�@�p(�d.�����Z�0�!��oISJ�8�������3쯵�
zO��[6����rP�
2	�����#<ܼ��p�Q�\;d�FTk3aƭF 3T"Bq��^��F���8�|���̄��;�ᖷP�w����F0��֔�gZi��͗��ti�Y���^ѕ����E6N����D�Y��"�����ǫ�^��+��	�h�~�t��l��by����y�\����\`C5�ص[��%����	�j|ϻV�^[&/���U:aIN�����2j�T�r9@C=w
H�B[�)�ɮ �	a�h���@��|���ߡ�K�]IQ�aս�~�������wQ�m��{�-���yv��:�FS���/����:QD�׀�Ge�F�x����h�
;h�����zK�[�ZC)�0hI	AG`�BV�sҜ��,�\�z���sسW�궩
ͼ\BAf�h�R`/Iu}�I�f q �h�kA<Խc��@����e�䄒&n߂Nπ�4�b����W{�$ɲ5j3��,���Ԝ��᎚@K���%���Ų�e��
�2�Oo��_÷��4߼���_������� ����r���|�����c.�H2��V�-3��+b�:�w��@b��J�B����_� Ӿ��M�8ڃo��Ą1T���E,YAD�5�ɳ�ʣu���E��J��hu�����hy�f��UA�bY� L�_p5<�[����%!��X���v�c|�Ww����#\�+��I¨#F��[ڢ �uU�4���Վ%���{͞Nծb����ђ8W��~Ч8�{O`���g/	;m� �j���r�C@���`�b��U1P��f�_a�Y�<�T � ��c�8��V�����������|ߟ�ö�jm,.�=��ژ����<����51l9�`�6�7 �y#��U�������ː�u.�c--,�(o �ސ�V�s�2u�x��ܗ5X��֧1�u�.mq�uX��?S����o�K����q�����Vi�26P���%(l���=�$l��^�kv�ld�ʭM�D�\�`�ɘ��Ҫ�5����Z�l��ץ�b��Y����R��A��� Es]s{��֗�r`�#�"�:G����aD/�h��1g����h�Q(���q@>��!T���ٺ���:���ۜ�����v��ԫ�o!HR��9�����h�%���̓7�EP?�(�����蛦�����x�}6�t ��h�2�4�Ħ�I��<uz]d��X -����i�G�g���V�ڽ/��@Sb��K�U��%�X�\����6-�5���Ք�)NsG���P;�u��N��^p,��#(J�]�jз��x�6@���C��t�`�M�Q�q��f�!��������!���f��y�m� Q�Y�8n�[�[�6(�,m]e�����bG��:�tM��d �~��R{�B�?gs�ΠR��ɠ�E��Da�Ը_�m�U@����ݰ��fkS��(C�"� ��%P����F��_|��9��l�Q�N;�R���r�˄���ӳ|Oּ�Gܼ���^Ŧ�	��b��[� 6��8L�o�PZ-��&ݨ�S&���04^@ɼR�r3�J)h��E�V�v��N��Z�Į��t�f����l��R3�z�0��%?�Nd�赗,	�=L�.���aİ����#4�P
�!�#��5��Fѿ��u韮r��[P�@����� g�L�4��^r5hN��b�-�ag,t��Ka�g�*���#Bl7�@W��}1#�!� !4A�#�a�8n7W���:����� �`	�*�<bsU�RP@&�t��@Q��Ȼ����/���;ZbvԚ#im*ղ����9 
K�.f(���_�a���?���Gt�D��!~�x_
}��	Ⰳ����r��J�?������2=��E5j}�>EU���)�˽%�L�[)��˼���baXL�y�Mq.Y�V+�F1J�#Y	g(U��S�U�Cj̿��!e���ZXh=���R�²��O�V��)�ZA�����Z�
-�&�0���1Dly�_`�[l8b3�@6A��#X(%Ϙ��WyM2C��pa`/�ܦg�ϏqC��q�0\a`�:<Q� �ڍ* {BU�m�(P��yH��@�x)O��noc�f՛����/��Oz&�:F�|�r2u�,Gf��:8F
�d޷���B!P�ҡ�	�)��4� b����YB�Bkˤ�D�ʬeX��
�T&�d��=��߶>ն��WyZ�׽G���'Dj����� 3ۭ�0��]j�3�P)6@f�!\>��	�fH�}N��@���Qfh$�m���k�w'�)�0�(K�s����,��:�ê�
y5�r=��i�Z�/#E��K��&�j��=I �U��.  � IDAT`,�� l�4����/!k�����Xe׋CN�qX��j����,G�t��'h`Pe/�2��i�M,`)uݖ��+c��������^�ꥶ��v�\x9@����7����h?0���/@�7V��e��h��[�TD���9Ȅ0[h�ە�Z�v�?�q�on�<�,)��ͩN�@���Z���T��#���4��B���*�..�'e��R���/�S��|�"���'�V�?�e���� y�"	H��֞C���tD�G���$V�2�)9Z	�����ĨEi��]-�q�J��"�ʹ%d�B�tDψS��ob%��>���j�Y�f^oՅ�0gT�ԕ�m�R���=�6`D넮��{�'#CsDF� ���]���-�a��.0� bE��(e`vd�DŁn0KKƠ���%�7�P��K��n�4���F1�0"���W1n_�̚.jG+dj�H�VE_U�H�P��-�V��BJ�}�P���dZ��b����P�X�ݩ6����C�f �Q1cGT0�3�K���)�H��Tg~�	(e��q�3�9C4"�F�b����{X��b��rY!ZVa��K��y�E�/J̨��T@)ٌm4��~�51��lS5�T ���v��
� ��I�#�8_����j��@a��Q��Q��ٔ�0�6��G�}�1`��R�ڌ���՝���?�����@o�K溶��'�;�P��,��W�Yz�=�:>��$&؋f�����y@�=; lA�L���
 c��V��{Й�׺N\@�Vהn���5:���hA��4�\�"�%!���o��CK�DN��� ���PB�E�uJ�v�0�Ȕ7x��6�6���ot0�Zg��/�Za@V�Ҟuի!@�����yzѣ�Ij��Ѝ2"��n��2�L�T���\�Zե���J���FD���nC
�P �L�8�/y��u���cl���� ��e�|�. ���4>��k����_ȇ�����2�@��!%��y�טۺ,=zƘs����|��jwUu���v����F�b�8a"% K��A�� +	�eǎYF� �KE
v�H�\b.����۷v�ۮKWWWW����{�5���9���=_Uu���|�m_֚s�qy�ϰH+
�T�����v�Ik��#��#�8�O��9����|��yR�*脶^���?!��P�IoN$3��G�Y���Pܔ��ω�?���^�D�M���u������3���'*`%4]q�O��Nt��`)x��>��z��b�{]�����U}��5���N(���5N?�	w�.��_.攈Dy��oƙ�=ݢ>M�7��K�X����At1�~'��ȕy�g�>��
X��+�T���dI�*�ԂR
��
X���P債	.�a���Ѻ�cC��l�[�L5����d]�Fn�A����@�r��
=#x���y�Y�5�ܨI!0J9A��`x�@]l��W��c:{!-`-@i����<~��~���}�����*�\��r�K�<2�?䱯���'I����F����)�k?�����hj����R����N�M����S���9l+�F��H}��8�L�R�(�W�z�l�`Hc";�~ݔ7��'2�W��+�\�i�����@�D[�u3�dl{����3��1�z-V���p�YUp�%��@�dj�U^;����p~@_ΐ� }�н�]:&�n�Yٞ����$Qs�qꌲtD�l�ҧ���gk���Z^��S�7���o~�~���(o���zk����_���x�3��B�+>����{~�>{�������m}����cP��ڞ]_����h�
i�'Y�WF�(��U��m:��c�8L�o�`S�>~�YD�P���"�?S
�Ջ�ċ>�<8����sl&�Go�8�Ǣ/�]��W�F��v(���0��$0�**���k{�����-�3

�r� ��� R+XTi(� *�V�Vp���k����QO�Q�/��e$����y�e�3>[߀���v�"ɨ�� ��+Я��l���T��aN�l���X�`��T�v�'}:_9Yf}6�T�sQT%q+F�z��өb�\±#��B�k\y��Uj�o���1YM��d �z$�4�;53��7��ʹSߡ���y������@�,�k�xq�
�g�j���	�ɯ����b���f
��=��� �s�	�}?	@��@_����c+G��m�Q���ki3���=��$\~/	�AB(����]z��_�x�y��7e~b�J�Vh�B�3Y�l� �D�_��'�t7:d���gg��+P�\�(�-��R���y7�i8�#]�'9r����bD(*)tKgٮ����ݧ3R=jq:�����s.���R� �6ݭ��9�����b;����#o0Іw�x�@���^���{2��z.}���(��Q�|<��Vl D��E��(��S[�����_[�?����G������b{����_no?zC�\�oQޠ�G_����}����z���������mO_�L~�>�����iޮ&�="����}p�>�h�xi�B��!L�f��3Y%���!w؄��Yu�a�/�x�<��!FL5����C�������^�Ƶ�u
:�P����C٢h�q�
��q�.�l\�S�C%,�ONjF�����l VT�(�g��	��8-�V<���'c*�>�ؐ�uW�����]��q��mX����3����"���ZO7>o��G"���C��ۺ�p��,X¹*^UE��]�5�鼸1�>�a0�T��X�������D0�*�p�B�5�ucT�j���QDy�����1�a`���N�Rw9����G�M,�JJ���:Z[Bm��nV��c�:W@�@���i���>�y������ ���v���A�R��@�6ɻ����&�:N�i�t�T�s{���<����á��u!C�
iF&%,��|��j���޷�(�>��@���$K�V�/Nhå�������<�@#u���P	=���+4��ܩr�~G%	¸,8���(�.�֝K���
��d8�B���+�Ā�[�:�_|Ljj�<9}L�#�iԳ N'�,
�t �k���j��- 䱫���������|������!�з_���;_��7�x��[����vy�ej�_|x�/���?���/�?��U����7~���Y���j����vA߬��*�;�wHo�	X��f��.aT�O���?-��yzꇈ�5�no��:��C!,���\y��|��=<
��B���S�N�\8��D��1w�����oq�����N�)�.T˩����j���
����	[��, �"��(u�¦^��k*��,1��R\�:[r�PyK�U���T�T�6��9��P<mh��ޣ�RQEK!J�Z�-%�v���kx���qQp�h:�g�F.���лL����غ�IW1?bEaB!E�B���^�)�`���(�Ƙ�����ķ�U-�B��x��h~A�Y�$�{ 1��4蝬����
�#�9W�� �T��Q3��D+��"V�|��d�� �+*���;�A �C4$Ip3*�G���|��v"BQ��݃�ŏ����Ӓd��X�ݠ[o�BG+�Re����A����/<�L�"�"@{�^ߠ���-����O�iUE���	Z6_���0E�z=�s'�ȓ�2�"3%�rwh��Yg�^X}It�qW��f����NP�է̙~�I�	��5�P�N6�7"t���� .[�hD���}R�1נ��S�D���P�h���������S�.��?[ϯ�����,^zԧ��sr��W��-Z��]�ٷ�K�<�}{�E^���ڟ�m�+z_����B�jB�F�!�iJ� !�α0{���� �yM%yH�U �=?���f�J��U �H�����T6Po`�J��ny�~LQ@���ï���L�=�*V��	�����ͪɹ��&�����L(�����<��S�����v@q�o/Ox{���U.P^��g�͊�z�sa��/c�*�Q[K�p(��Z�	`:�+�@�9?�����쫥H��6��A�1���G��ɣ+���X
^?0F��3"h�
R��3�R��pm �Tl1�\ԩ_G4@Xj� �;ZS�n���HV���1�?8e�<R����L��t�FGEj��܀��+Sqv7�uq�n/1�>=؜t�|�B�����%�w3�_�hӣ)}=;������8}��|!�(�o�����rҕ�H)��ie��������̍NKz�N=�
��������uȋ-%{:
�A���3X�TـM@�t��i��>$�hϠ�-�]��[��d�-3�Pj�8�O�zE�f�E�����I��2yd�n_<���J9�Q�
݌��r�K��!o��y��p�v*d[	U̹��Es9�2���r�t�����
�N�0(�h@�����;h GsjFwN�X�H��a�=9�*5Eӭ@�?�^�~n�G����7r����|�>����ǅ�PW\���7��K���|zD)�ԧ? @�'H��Z��v���f�U��l�8����~3�Pv0W�~��K�1�/�̣K��M�y��H�)mt�x���SRoW#�F*�F6	���+��񏾧D#Ű_�P&,���wҨ�Y�DVi
Ewv�M�6<h��g������9�#l�.�1�D7@7+(%2��ޮ|�UW�z�U.h�rmD���R@'0�<�e�`DE���M>�P�L����f�5�
��٫��<x�Zn6h���5�@�&HY#lq��P��2�
����6�B���{�s+��������G���	��
ҫ� �^�'���$.w"�tTu؍d�:<>$��+�O�x��&GA�k6�tre�� ��٠`/�R��|Z ��O��y3��VK�vg�}{��Q��-���|h��R-�B>���G��#�6շx��<p(��&+���ɍ�ʒF4Y\L?���m�t�`�Qg$$�v�d�]BP��q*S��B$�в��o㍻��o��Z������V]�b+��+П����'k�9�B
�.�ֆ��f��r����q��M�hJIL�H��(ȓ��BE_�~Q�lЭ���ë�q�aNw��`��
ft�X�����LK�68!2� �X^}�V;	���(���Ay"�!I&��&� %S��(�Q�t���v��m=E��`��p}���T~b9���?/��~��X�y��ׯB�!�l��v��_�"��_Ƨ>�Y�+DXW`{F��]�_[6���@�8,���10o����(���BD���5u�a�H�d0vB�1hͪ�IɊ�8f�GH�j�$�Z	Ee��5i�4s!\��%��$�yq�,�6�,L�����U�ʨ^ ˂^*6U4o���x8-hz��
\����9ٮcE��\�[,�!6UlҰ����EE����S��&`w\�v��-9!r����Q8-ֶB��
�E �cU��j��@B ��H�;�Ժ�dC�M�8�ՙ�xR,��Ʋ��]	�z�e�@W�R�h��;���@A\�PϠEAm�\Vh/Xj�b�z��6ԥ�C7�W�mw�MC~4!�(�DH�8���0�h�8!y1�.(w��j7���xP�ttS�tk� CB�-�0PJ�/�yO�����#X���ryB�P��j�_���1��yd��G�R��ܣ�(f[2sVd�c�]l�FW��2&��\����ȟcgB�{���Hq�s
�21D����m�mC����z��S�p�J��[�R��j���ؖ��2������?X.֍kueU�����l��:W@����'$�d��,7Q�A)��(
u�\T)�5��2G�: �a|񔎢A���Д���Rn�F&�Q'� 1C��RP��&}�ٺ^A�
��J�K�b�������罭��e#`r�4�v�b����j��D=��T/�44R�Z�:$��u]��"��g�]��<���6-˟���oy֟��F����}�����2-ݮX�~��7~	�w��c}�Lܝ�]�p�{qlD_� %�KDgn�)����/�!�8 �)�����G�Kǟ�s�=a#F�nހ:j�4�����{�O�}mx�/�����~�4�{ ��;�'�|D]6���+���Sõ_qٞPE����	B�k��k���䊭=cӆ�b��.���(Y�Ђ�Ū޵����W��A��2��n4��>��0JF=r����rS�JT��`�TL4�,c@��٪@��P� ټ�ETr8�Q��t��(l~�L̌�i��E
����BN�NaWb,Ո~X?@W�ed�(���T�z9��D8ג
[I�����FT:�!�v(W,4C��9�62�:F-�XM�@���P~Ƅ2Ph�f
��9�>���w���ޕ� ��զ���d�(8^
z��`Q�|���o�.��g����@�[]���zG�BA�8��>�Z�k!���]�Y�i�&��w�B�1��9�cLg8���N�XJɌ��v(+:YMJ�s�^a��:�#VT�i�n��E;��aݮ�v�yfݩJ1���3�H�<���5VR�+0X!r�&��g�U:��#3=�f�
��kp��qj�@A 
�O��A���f��,�z��CF�;�����5�1r��Ό���M��7�<�v�_[١=Q�n<}��R~h�$��7o��@9�����{������������Q��c��
���;�	��y�m}�~y�����*�p�$._�9�0����c�`��1��&)�o��;fJ�#���o�;�J�Lč�i4�7Qls���~��{�AO�}��_�!� t]��36y�ϸ�g�L�=�\�X��*&�mõ]\�+D��M$5�q�V1��F��`�����
 �] �B��c��(�{����ChV8I^deժ>瘼5���[4t��i*`W+�"hm��r�N��
:Tx��Y��$��	�d[΋1�5�iw�
���h�lmk�O�����(^=���%ИXd�y Y����=�2��0�AK�����A��D ��o���Fa���EUS��C�+h��=��8�+�Π�ЭB�g��{-ZP��gm[�T�
�~t���)��5t)��������	{
&:J��$�P�Ls�3�>:�{W�Y8��]�r��(�E�C9�����a�^���wb*G�f��*�u5�V�|��i����jzK7k�m+�]���]ѯ�6U���M �{�'r=GzpvZf��ᨧ�:Q��2n)	�ӥI���j��r���C�B��zq�9�V?eN���+TZo�����~|�&��χb��lz0.z�?�պE͖{��4�ϵ�	�i����LIa����W���t��S���?-��O�����˫�!���J����:��a���O�_�~|0:�S��F�2�˳:�M���ѻ��m�nu����bFr��LO�/Y��x��$#7!<�8\�Ccj��o9�o���q�Ј�.h�T�;y�&,M*"<`�} �L]]����z��p�J�x�x�+<���k������s��+.�	�>� v�%��Q����̆"+dSl]P��6���	Qṩ�f=: �L�:ds�85� ��ә�@6w#_��y�v�P\Q�l�l�n%JP�jGS��Bj6�����X7l�Fѝ��7lm6`[����	}[�[�R��x�N,`uR*�x�1s���(�J%��K��a*<e��.���9蚽�(@�y
n��[9|��5���<X�Y�n ��H zs�+tmЧ��7_G9 �؀B�ӌ���pxzKT�"�Ha�g�{^�o�L'�����_��g��)E5���Nۥ����hZuؙ=%Aݘ���/��>F�rF^,��`��͸B�o�����zIG!+�%7L����BXN�4(�]8a�w�<Ń&���"�>	���5�T���0j�/�U��08�UBV2tթ�3C�*��qdH���/�kV����ޝ%��9����H$�`����slZ�q�X?��~𖾜�� J>k��������g��������K9����0�z�[o(�	��4.X��'�	''��= ��:q?K�aO���4�&�Q�	H�`(���w�����v�~Sseo�	� ��Ͳg}xD#J�8����c��=]0AX#Hl�`�c��Z���D��bECG�R���i�z�0:z���]m6��1�i�ł��7���+?㹿�S{�k�"׬���x6�f���\��).�D�Oq��ϱ���A6#5'�����`|�$��B�G��m-#2�Rs�T*�&u�֛o�=���E���s!�����K�"��o���n#�\)غ`�����x,��FDUlr�S ��ȳ����i0�|�ff<�N�5�E3�1�<��|5�{BdU�������.gT4`�B�	R��d��-��7C\�+��
m@��Q��).!�e��}��:�T(N���Q(����h\T!2ڙ�ԁ@Gwzt�|�	�TU7��|r��L�թ���q���<�Q9�Ե+:72�aB�\�׷~@��TG>��P_�=���\?�^>�\?���z[����[G[;.��u����� UΕ��n��w��@V����Jwƴ�#�G��m��)o�\!A"dd. G��@�D� yoŃ�pܠ��!����T�����]�@��K>�������Ǫؚ�{��i�z�g��m$��sFJe]�lo��#��Ղӫ�^y!ccr�׷X����V��C���'��:�sB��Ob�(���&k!��6�`�Ɓ�ӚE?쯔�@��m�C�ǔl�X.�`F��C�Q_��wK1��;d�a�v�т��;�Q�:ǻ.غ�/��s����PX��$�njк�k�nxӁ�����{���y�e|Ծ��훸�7`�Xѣv���UZSM ꄾF�����e��  Q�ut�D="Wl~��Q������]�`���r�a��8�0gP�	��h�hM��P���L�BY*�+���P+�'��J�V'S�1ùsAg���a� 8��&̚�YD�ٌ�$0dDd|<���ߴB�:IED�H�n��vf�b�+��YA�`���J�@؜�� /�,'��ڊ�r�"�b�B�3z�,��~��P�+t}��BsZO7WN��<z4Ek�K�Ѡ!O�8���3��[�w�	��
a�ς��fj#��x����"�D���Z����)E�t��z�^���,��xOm�6���<}������_�-�!��IQln�ۺ���:G�r���N�"�R&F����i2��Uy�
{����@�ϵ�N�S�$*T���^(�f�l((��s�[Nei��{J/�3e]F��82qWLޝ.�Ƕ���j����]�\̝p�%�^�J����P�9�n[��ޒl���rap%+n���_���_C��W���HcC���s+��ibˑ�����tSp��{ĳ70����vp���O�Zk��l�2���ߘ74�'2��]�t�˛K)�%�h�t#!���G�	]�C��JX�к�����&�d���
��N6�h�hҽ�Ԕ��/��|z���o�'\�W�b��sW5�Vچ���u�t%)N��iЅ�OQ�2r���s|�Y��#�ɠ�n����hE�J�qL!	��g����~�i������o���� ����4T&�P��X!�n��X�^�:���NU�rfs��N�P������9��t2m@hL�r�����y-�M�M�)��Z*�m�oP�L����ؼj�O2ť�����[����� 0Y�NZ��>~�I��q%���������\&%�8􈤁�Y�&u��mhP�E94�w�z�� �H3z=G��D�Ll�g��'X�@�؞P�[$7A������,*m}���u�� �o�/^Z��ۊ�:�)����s��������m�>H�kBZ�e=�Oq�?W������R�ѻo^�G��!�NX�OT�g)x�_�-��� �ڞз7��Ջ��ta��7��4���#f�T����3n���1��/%QT��@���[��|Ӂ���1C{��.�UI_y�	� �گ��~EU��kk��2�c/R ��z���%�8����ɥ��*9�u���P(1���!sZ@T�Z�����
�9L�^Sю7��P_�(�	SN1�����7����>
�f5ցgB�|y�5���A�����'W���0o���Tl�*�����}�t�mo�XW,� �pU�"�UmD��Y���*!�F �^�D�Ԋᰏ��� �%�h_/0j[��"Y�N�DE��`9��;z߻������=�5��FWkœmZg��j~�J��ֳ���U�z�支��V�b��k3(z��J~�ݨ5� ,rX0z�:H0%�Fp��N+F�="�ؽfa��C�ʚ�*�6(��cR��R���Ũ �~�� �0Zˏ��@V��M�������
*����庁zGc�d�AB'��ijhHk@5+jjT�Ng�9�t�����N9,��u@b�"�������u��8KF�dϑn�!���sC�J	w���q�C��P�Ů ���Ӗ���U6P{���/�П��X�'�j��-����7X�>�N��>w�U�}�X���s�7�8I��S�}��U=�:8�^�z��)W���J
)�*�6%徏��{K�=�ih��M�x�{��R"ڡ�f�t�v�����}��}�� �W��͂T8\ng�F��u� (ڡZA�H�ϐ��6���^W2�,�hc�à�)-ÎhJ3�e���eQk{]��3��a����+�Ӓ�i�S?���RR;F|9�p��0��*��d�`�:`���FN�y��Ë�@�x���y���B�+��]�e�d���!�}NP ���8��"=[��u���u�<9{qQa�@дa���@���5zF��du�Hq��¯p�U��t��64����gT� �8c���[{��dR�vs�:�)>*��d��! ��׾yk�5&�����+�y�F/���+�(�q:�3"�����7��+x�,�o�n[S���������Z��)s'�7)ˬ��H�$��A��ۉ?�<�M%��pBU��]��
Ō��W�h�
�iA� zD�oW�l�A��A�|�z��N�/b�$ h[Q�'�u����xOV��a���1Q����`T#i���B=��G��@%��d��Tq$-ȵ8�S��*2OӨ��GQ��k�:UD�ӹ6��~��QHgU�$�������|hV�.�<?���[�4h��}���� ]��+�nX#�g;����0��'3�9)Q�"f�b�5��&d�Eq�z����<󁎆�R2�F��t�F[.�"
�F
wju���(*���L�"`�&�;i�8u6G$�Ug���$	�:��P�z*Ղ�dnd��Qε��Y06ul�	�	�{�C�Gk�oF�As�-��ذ<DԜ#j��1�~�PD�/�تs��Ugn������B9j��&��Nަ|Qn�M���ܞ����G�x�y�Y/p�u�I����l`ݬ �/\5�s1c���a��醆��l�����*���1D����_��'����Mqך���}'��!M���(Y�����c�J�a,���	��K���}�q������9.�(\mNr��`9�ZNX;akFw{]-�ۚ�DֻN����hǶ�/��*��a)���Q�zm�y�Ԝg�� ��y�C�����n�(�w�k��f�5uj�h���~
*?���`~��^�^4�D;�X�?������������T|>�N' ''�q�i(��#Z�hr[�h���2��a��#�����O�����L�����8�}΅3?&IM1��3�=�0�S�m���ѥoB���6��,` M6���>���3��'�������z�v����
��u�X�ڝ��c���ѻ];��T�	����ޏ��1e�L�F���ӳ�7������0����rA�ϐ~�����{���D�͎��o��C���g1t��ɓ�E�fsS�&Թ/L(]�xGd�Z�;S��������w}��V�6k��+�snL^�{6���8%3�0G iؼ�8�)�d�I�eZ��x�	�U�b����v��`x�Hd|޻���:���	��:�`*"h[б��B��rE��[6UP!H�·&V���4}���7/�s��Y.�1H.f�u��/h�-:@�-@)SMA��!�1̀!�]s8'�Gv:s���ڬMN�ރt�27:��9R=��N�D'��(f�A [�>E�r�u�!�-�
�W��ݎ:�4��2�X��"(�)0���:������:bJ9�#��r*�O�<�.�.ש@P)�#��^��#(��VeDE ��N�
���lx�:]7�ј:�I�@{�<9gy-��P�����#�@����rD��9���z�	��=Χ�L�:�8� b�̓ZtD�B��y�kn���]P�"�����u,����B�+��g��P\�|�7��5\޼�	���u5c.��ʨ�V��m�d�,�Ϝ�~@���O?�g�>nJ=�F�g~]�hO�HI��N[Ic���s�(`����	爴}y_������'

>�ƽD���`�<��ݬݬæ��$#r��Vp��H�H�1���^�nW�^��}�1ZW�ϯ�u�z}��x_3cky#P2�!A2���7�p����ޞjrI�@��Q=ڧj�[Þ0a���g���h� �N؆�}��o��8��M��}�5`{�5,�� �`�c�>uUl�{�T�T*V�% `��M-m{i���
�킫nX��r�"2���M*��:)r^6� �g��U�=� [���yn*H��vW`l�"Q<4+��%ۍ��ݻNQ(Ie���ܶ��nx^��J%�Z,��<GF���ɸ�;YL��'V�^��`�
wDME�:'�9"�@��~xr����RG����[�E�K��k�Hv����h4�1P���h5�U���7��3J=y{����(%&�m��HV@����@����Aj`��	���c��ڤsxR���_��b�U3 ���������pB��޵�Я.S�^�����B����ր�!W`�z��]�,`|��_�}�7�^���m}ݬ�:�IfN�"W��Ϻ N�q�F1�Q�{�)0��h2�����fyJ�>��αWL����������~��m�4�TZ����#-u��)�V�i��i�#�3��_RH�l&�`���'���F�:ə�\�pFb �TjoA|E[?��7�D����M+.�'+��x��� �?�� L8N�&�g�^,v4��q�q���!�ʱ��ا�}���d�!�&
�s�C��?�!�?kD=\K�	`�Ć��+V��j��

0�d)C� 6�.T�Dq��U�EM��8B׎���'yT�o>K�ɀx����'�ݱ��_1��Y[�qs�\�@_�_zL�S�ۖF{���@9G���{������%��;����
<oƿ0Ё���u4� *�xA�hG�M�w��x���<�@���C��H�lǡqE����c�K��u��J��i������70X7�� Z���؜IU�bI�{��=���b3�9W9&C���Mz4c*�P��T��EU�,��ͨ�H�"=셭����%�猼Y� �*'�,6.v��pwN'dk�q�H$�LA�ۆ���7�V
J�3���z��u�mE׎u-�����5�����3Dt�>%Z���
T3���=���θ�;������]|B����D7�zE4������D�ܝ(����@��9.�y���<��`���H�Y�:��p�	lY�E��*�+�������A�#F��l++�ШCP���7�U�/op}���4J)�}�z�ڻ���؛��hIF �t&�6+r�ۚ���ꕂN�p��gwrǫU�w�gm��� � �8�gH��y�q�$��#��-����ݣ����l�\��3?�ay�C=�B�mOX7E�ŋt4�@��)p�+6l�����.];�V�����#�oO�dÎ����S�n9s�d^˺�"*�*�h"ن��E�|$/�MhR�;�fhZ��6��H��+	�>{��u�xz^q��{�a8k��$w<Q	v`�Z���:Z��fc�;���E�P�Aey��`߶&�A�C�����2����@:���
J$����8���(�kcE���
���m.�g����[t<i���h��Qt�̷H���{���֢(����E/i��J�',>hMF)�N��X��Ƚ��^��>R'� ����ʶA��f�K�6(f#i�9SNy�`�^wk���36�Ƭp;c]:�n%W�z\>�׷oPT�ʸ�}�δ���zE�]P����x����l�뛊ys�b�&�#��؍v�Dt�i�<���>(�]F�7��ؾ�������\v��uk�N6�r�Ń���]2�+i�1��8����裳mS ��R�#�Ք3�;WOqG�^�{�u�&��U֯����h�ety���7���uE�T��]!X-R��#��BHN�*�#��'CRޛ�Xe�Y�>)���-�O��� #��I��)"�ؙy�G����"�_'/|�@i��*B���T�E��}�*V]�;p�
����>j}g��~�ju�l��:�l&4:_��8$�s�+mt�.�O����kG�l@�/�w�Q�TGof^�P��;�v�<gJ��D��M�% ��OnZ*�)eC4�e�_�+bk�ѵ���-�0�#�q����V�aU��wl]�MQH��F>�+��3�מ7��o�%���8�*��N���\���Ly�"�X�#�:.�h(�����U�éKm��ϥ����hs��.`}kH�����X	��RFR/�2��ΣݿW��l�3�_@��ܖOT��O=��ߕ�6��|��F���,b�C�1(V��%�hf�\���(��Jg�#G�ԞQ���Ԋ�H+����ס�(���b�aU�`������ \Q�(/V��l���>�m+��NX��uC��|��i��m��z���2��=�O:9�:4�>���{Ę&��Y���9}f��iD iT���II����<�	V�GD�q?�:�~5٭�ŋ;&A�Rk�C1<�L�&���M�� ����H���P��}�m���ذ�5��-�&Q#q2N@� U����'@�"���=�}
Yӎ��Vo0#M����3�-����VF3}h-SԚ �k4�S�<���.��qB��=p�9t��Y�����Q��ݼ&Q5K���tM�v���.����*'\�׾Z�I ؊����s�J2�G�~h�Cx3"��Z�t�[.��V�:%�,(�9 ����ek��̧����I�����z���S��lQ���o�B6`@Ĥ�����ņ�(l�r���&�歞�h��Ώ'ŧ�~�x��R�)��]͔�a�������ԛ��E��^�s�$��k�p��@:�љhR����Q1������֙�0C�N�h�ܽ�ɹ�<r����[�����7ٶ�M�3�����cT�?�+a~f�i�B�ר�>�ң������3��gyu�C�uK�j�q�VX)I�R������m]Q�G����Ӳ`SB_W����Y}r�)z�O���h���'�v5^�-�F v��q���*�}�7�8��p�"�KcJ�HŎ��k�G����9�p�kc��n�|x"f!�|��a�H���Qw(F�v �R�)����
�gڜ���W3��l�z1�<F�`��R���;c�>cY�Z	��h���W�2��kBS=�|�g�VD$��צ��N(��0Uj���X�r�w^����E���Ǩ��T����j�Y���ȧ0k�hF����������g(VcC"��D��'�4���sdv��S�s�s7v|�~�6�<�c�6��k<�Sz8���-��y�zBG���G^��*��=2:Ӂ�ZA\�1z�dd0��p%�R�z\� ���r���,
?����W�K)�L֢e���;���"�ދڝ����;_e�g�]�{A�C�U�ZpN[*-�Gz�X��
b�͘aC{'�Ԣ�;���[ݜJ3�An���UB��;e����3��Y~v�iʢ�렰3���>A`d-���\��o�yK��p�l����k����{�ضRB��\�u3Z���#h[�Z|1*Z,Z�1�Y�n�j�i}���
)ya��S� �w�9�k�N�~"��Y��I�K��#9�=�B$I��Yu{�y�+�=A�ã������������d��5;!��U;��\u",KM�4����fr�ά�Pg5k�J�?�瓳c]��Q�!R�)��p��
$$!v2>r�79����:�C4���}�i�U3B
\w����������;zX''H��/�߾��v��p����qe�צ�X�_�L�TP���{�p��**�ӹ��0 ε,݇�(;ч��|��!w���G/	�⛟��܃�b�9��/��(k��&�s�8�k=}�D;ۻ:{t��Ϭ6uM"kI�����b�GN���Ƕ�'�w>|�x���0:���_; ��}�2`$�y�宋���<�
�\�8�X��[��~��	�V��*����f�[uv�T�����yad�R]�K�S!�1`�qpn4��=�[9�c=0����i�1��4����hO����[t1΅������K�?�
S�_��]��?��f�Sx1jYe����p]ַ�D!q�Z_S%�T�3 "ض��̸-N���N�N�;�`�O�3�e�kh�42L����b���,��`��{�.�����Df�O�32}��A���N{!�h(��:�r ��XĈn���B��ƀ����<��T1)1�?k����	�Bu9��/+�u�i�ц}k���xof#�E	�����+�ً,���X�#{so׀\^vv�abЍ��%όm���ΌzF�:��X���=�2�+`��eF�kְ�O�C�@��\*�r�Xk[�xLAZ5'#�a����v/�2��{kY7��G7y�I�������	FSĉ�[履#��)꜍ݽ��D���q��b֐���F���}�ӁOc���fk y!f�X�U�{Yp����
�טߧ1�B�X�;�z���5�!�8�G�E ��=�EyF��9��8+(
ubN7�bx������$E[aF�q�������^g�]'���ܸ?�=����@9��@�lW���͉.���@��}dlpB�MJd��J��qǪw���io�ڶB�b�v�@a9p�h�:��y �l�[C��Ō�f���d�-z� h��H�Gn�����0�٠��u���b�N�����G�QgS���=�b}8	�:�;�p$�H#-�4;���kĲ�R���:�|P��Y�\^`�Ҁ�#����cumDT��tA�6<>��ȓ�FX�{#�����ʾ��!a�>�������(v�zG�-�_��j�9?O��!�����[>�/�������ތ��E�6 %zh}�l��*��x�+
*��Q�@u�G\�)����$6��]'�A��E~S~Ky�)����3;6-�{R��Os?#�Q������#);X���'urVH���'u熺�ִS��=|�58ѣ�"�N�X���(Ҩd����DбΑ7��Ý�6S%��6�ܽ��2�mj(Σj���g��(�	��`D��v��ՋWI�n�'NŐU[s�h3�mFZ������cu���e3Z���T���^"��D����
*>���0T�����������2�)qA�շT6�ZAUP���X퇰b�}�ذGY,�V@A��Y�7hW_J��	G-��YާDtzɹ��M(�I��Q��lu,}$Ӛ�2 ��0hZ�]�?���o�srgh��=��!SZ0{j����7���m��Y��EE]1~��ʗ�)GG�Fu�v<=]QJ���ds���� l�7-%6�V1R}G��(���	�|˹�������$�6e��gR��ְ�`����c��_�pA ym�*��*gŎ�!���J�y��3��jᵙ,�
1�\7�J�/<���39��􊮴�jB��HD��J.����D��,���dq�=�0�\ϑ�9@d�P��K�s���ư�]p��>W�(�n
��e�2J�2j{ѓ���� a��h"�?�΍kC��3�y����G���(�ʳ�^1������;3���-T:���q�~�Dge~{`�-���ɻ2B��P/Њ����w:oq�ُ��U��S��+8̤KȽu�������z��5��ȿ6T���@�̤#�.θ#���jS��DֱAu׺X�T�S*
��}}F#�e��tr�Y�h]aL�+̰Oŀ;�gBG�3!�߫��Y�7�ى�����|��%�c��ĵ�:M������H�#��\vNǄ��^�uN�Kbסǥ�3��O�km�b���r��G%�R�4��,"��Ya��] �?� �����+D�?�QСX�8�"Yճ{��:Ȟ�E �9���z���v�غqZ'x&�!��"�}� ��Ө�r�3������Ɏ����ع|c|��F��+ht��)��	%��lchO�~FEEe���!��Y�����k�h�{�U��&���� ��z�#Y�]*pf|��l�=�x�2c���Y��ӛ�T_�ݑ�Q�������0�>�n�.X������]RaĴݮPqs�/.��Po��?Ԭ6z���E��U�y�DôKP�F�-��BvSu�vKE8�5�2u����2W�n�GXgB�Y����V��A�)}<��P� v�(i�BV��yĮ��J�w�qԭj^��f_6� �v���3�T$��!9�0�V=��x~N�aLR�a�_����߈ '��ƹ���O���q��{��3�����ڬW���=�b��\�@�X:��Sk���mPK�:�1����h�!CβX��4E@���n�/v'Ҁ��p*Tu�%l7�io��N0tM��Ri���H��e�_�S<�p����b*7'?^�;eb����n\c�.{7�@���`tP�:6����g��W(*�U ��j]Ћm:�a�>�&�	~��kh-K�ة��ܴ;?�S�ŰG� ���Jӽ$CɌ/V��[�/"=���O�"q{C�peJ�_�v�L@!Q�9�A�����C�c�|m!�D�aRm$l��EpXA���&��`��?ZG(ׁ\i�lnuN�b�2�!�k�@�:�BW�4�W"�}�����`����9E�~��制��{䮆Θ�7x�a�a�VKZ�L) -��&����M]��3�A��[��-�����)�0.
�&�������)[���&��P9�sm4*��4����zEi��0���r' �G�""{��
vN=D0��l}���zH���J�]j+(u]2l�Y�=el�����7�k"���K��h)����o��?�t֦6�� əR�eM�3Yx'�B���A!��TA��T�x~�n7���ޡ�c���{1�5K�$��@E���S���6�x>��G���Sƽ������B���tDZ�%a|�������3*�U�r(��@M��r��4x9Bv��m������Q,2L͵��X}�|N�ޣL�Z���* �i཈a�&R��Z���64�C=�������lR��hq����?`���iᮩ�~��_�]��ʬ�&���Q�p�sgOt��p�\� ��s7ex��������|��&��T� =���hS�1�1h��n�]����!�a�"s��ØZQF\�-��7Fc���K:���h}/��������ޙ���"����H�
Y��"Fܐ��a�S,���tϣ��xTw��<B )��q88&�p�������:9eq=Z��¥���vSR�	�*��C��b�������xE8WO�	��N��$����V�fb�؏{����{�{��`_=�	�� L4�ҚFoO���X�]��+Ԩ�/%X��!rsV�~E�(���\,�'>a]7\�+��+��y�fuA=��HpI�2�=�w�3{#{�u����3�����QX���榰�et0P�|KhE�+TW(�DHc����8[�P�M��Z楓]z�a&�1�׾��kN����G�z��� fF)D
Q��EP�BE����EQ£p�c�t��_A���L6�!��@z�T*v�uN��d�(�+�	�@�pw��+���犃�4��0N�!�`�CT4)�]!��w������ �� �v���
�QyA�j�l*F��FF~�̷�X��Ƹ�y�݉Rd�X��(�����J06Xq���;�k�W�ɎG��?���;����r2g\'{Q\x�ܒb�b�����"KR����h��w��|�|�At$#��;kp[��1����y�4�/�-_K@2��2�|��u�.(W0�u����]1:�U�A���P�ކ!>Th_e@���oPF�f�T��5[D�\ݓK+���1G8`���N@ɴc�Ƿ���Nn�C��e�{&��Z|���IϿwtti>�h�TF�6�vу��oX�뺡7A�n��'���3`-�u'g�\$<��u_���$������ڞ3P�q68�3�~dN��
�>��
hAg^��\���q���F9�����A�~t+�w��?��khl�KJ)#�6uT�ʐ&�m�E�bJ���9]bV=¢�d�i	;�S����kG���qgto����B
M|/�!*�'c��^�/>'���� #r����Q>u��x��
i�\v������XE*/(��|oX�������N�9X>(S@��Hr�A@����ɻ�K���e�s�	��N�P�ݪ��G ��d�B�H�P�
��s�5P%�t/C�ja,�`�֝����ZfJw�f�Q<�ֺ��I������{��#�?�H�?�C1xǮ�ńL�=��p��ו�TPJ�p����@���(�6��t2(u]�PS����}TFߒ��DL���-`w�>٨cB�w����f��q�;��RHS �ņ{*�Y�����H����+3����j�~{� 5����k�P���i98��;��z6G�Q {���O�����}���2�hu�4���B��,td�y-Q��f$_�, ��lG�H9	��,�cچ�ܑ��G{��i��U�V�~ھ,��$0�� �]�ć�
zj~���0�à"�ao��W�3G�s��8�)�;d�n����ў$q8�u�q���u�T=R@��F��J$�(�	�q�&%cn"N�C��Rt��(�o!���m�S�*�����C�Js ug|n���z���u�#�#�L� �~Un�B�WE�������	(�r������O��.}��U�/�ϐ�ŉ���w(�c�=Z�cY<;�q=�Fw=S�����Q�P.P&h'��oA�Q��yޝ���D㔎�gx2Q�<;�v�]jfT ��dw�S>:�G9����2��'>#qCF Q��^�}ެ%R`P�.o�v����ӂ�*����e�[Jźٽ�N�Ey�u��zu��,��6�o�Tx��60���uO����������x~��u��۞t�di�m�l6Q��+d[� 3Z*��ܖ�� <R�ש��&\LoG������G�z��t��!�rZY�f=�vY�=�E�Iޭ�,������	�U���b�����|DV�zz��Et��U	���-E�˃9wpq�ˉY�B��5TI��Ü�F���hB5�3&���K����p��{ւ�DN��G$` [�� A��٪�_É�������E�E]�U�yY2��8x��=x��_�ϛ�d�o�ҳ"�?ؽ	f�
�ޞgU� ���e�1p����o��WhF7�KG*�����j��{�D��޼b��(�ؙ���J��k���#6��)�d w��ą�6�e=�b�0N0��c{�c5�,i��a/}�j�=M��ٺ[� `F�D��m�Y�����=�!���"�����@ղN&
��ȏ�����cT8;s���o1��U�^��gU�R*��Y�0���+r��Sj��5��s?#�i�H��T�Щ\���f��
B�>\��1DH-c<�X0N>�mr��Y����i	��S�O)��gبy�>y���)���HTP���X!��l���B��:W/:у�<9�f^����(��)�>G� ,�t��ѓ�us�2Ⱦ�S��+TGaBx��U`�(�@in'�{׻�Ez�b��A�#�M�%��/ZMjDV���ǁ*T�Z� BJ�9%�ݞ'�G�ad ���}N~�j�,?_I��T!�h�u��'��5�e�>�2֏�{����#��$J���B�=9�uc<�y?23V��Qٔ�Am�y J���,ŤS'����B�.`�!�׽IG㫡l�����ȇ��hɋ�#��L���¨ѐ�{/�Q��U�S�j;�����
'��R���������vM�ɗe����^�U��b��"Ppj)4"	�yB�����!�G�yr��3?���n�i�\�$U������;���8�w��v�?�T��r�'�}�ea��6z����b�z������r�(����Ʊƴ�ӂ���j�]�E�ur('����K�ND�z1���q�P]��snU�c���~�D���c�p�%[��
��sC{#��%�.��>Z���A��Tv����fX}��d�-�r�H�t�*JN�BǞ����Z�n�n����-��0"�o��E�PVtCl �A�������!����E9���-��ux6����aΛ��="˱�aPF+�0�(�4�Q3�H)�`��R��=�l��E���sX��m#J4"t,b� �	_ǭ�G3X���
 �V��)�H�1b���g(G��u`bp3U���É��}��C�9����Y'��>ϕU���^�;�؞[w¤M=��M�2�zw���\�@�l��ȹCt�`OV�(6u"���5O)��8ס�2*�<z�;^z�3�)&�]c��@�o��o��b��ENЙ3j'�j_{]��
�5��q�
�A��@ݠ�`Tu��1�;��L��g��C���D�GO$��Q>��vK��/^4G^�a�3-t����{�]K�� ���u�tA���O�6��Y�2>C(}Ak�m 7P'ȲX�{]@T��.'�[4�����̎�]��U=�GE�X3�[c8� �w���	�sK��s�P�^�F���;lV	�i{F.�K�[Ѹ3I���vvhx���l�ehiP�Zlt���G�o�X�d3����6P���A�ѣh�l�������`��//�P��D/Wb��I#7��m��u�Q�8A#��|�c�L���1����;��/j�0o�+���)�����|�AP�$ƿ.`e'�]d��`��E����N�)0�N����G�kc���-f�V���6g�� ��!
�j��co�:2_�Q�'.�|b�!"#:�mI�%�(�Q�}�o[�'ӹ<[L��jI��B���2��?;-\VurJs���;O�B����U����fY��{ħ�t
��3�#S3nh�t�|h�
q?r:_�~F����Zv��LU����Bϼn���C�=���ƝR���#�����+My��5>'΁�)�#R��3��k�^��'kY3���u�)/��
�܉(�X��;{�ɶ��m��(˂�,�Z!��bw��/W��e"��3�c�ݎ��r�����@���;>lZm��A��� �~�T�?$��Fٜs�w�v�ns�{:f�'�GF���(�E��1�9���>����I���f�IFU�$���((*�WP����w4(��0���l��B���8�܉Bo����q̥�Wl����yq�n,]~s;�sˌ��l��f�΃L��;���3��g�1D�CW8gT��I�/�F_R�?�<��~E���m\��UD�/%��&f�:�o�q'�6�� b>#�*_w���vg&���?"��7Г(���)���ǣ
9qdn�P��w_��0��ş�N٫�Έ���s�&�q��`�8:���f���s�i�i� S[������m�D#}ـ���,�P7�T��
��E딒s} L���N�QR���q���4��=������	����I�f�!�w���*��ED�t�S>Q��Wmv���b/�c\�6�3:Qje�n ���jƜKF}��=��0������C��:�[Co��a�#H��]_���h������%6�A��@��E٬�,��k�A�T7��6� F��İ@���X8�%��sDO�l@�73@PU�kSH3X���ZE�K��s�5;�S�� �VvBI��`���ts3-/D>�����=��X6�r����i1E�C%��G��qwo�;D�=��M���Ӑ�@�B
���������ܔ����W�����r�a\�uν�;����Տ\�-���9�KQ���D����`D��}�T�NF�&�r���$'��dF�a�ZԸ�}78X�BG�HU��'&��P\'��䓓EJ��b������5���e�>�|�`�06�p�,R��8c�t���H�&yn5�J(���A�6�Ċ��8��ts��,R�W�i�t�*�3Й�}�p��3�p��#�r�NU�;���p����E �,���	�V�ɀ ��-��Գ�������[[Q��. .���[��s�I}�'��!����㬏����ry)B���y�7��7F=́�Pv���o�Na��N���B⻗c)8k����S��-κ}5���oH9r��$pn�-�6eY��u��2 l#�I�,����Ñ�(9U�*�����T�8ˊ��[,8�dy��c�n�+G�oB��K� {��dnQv�����^���^�;���ѣ�?N��".ಀ�Z^�#D"��U1D�C����_�������չ¥wE����K�Y�g�F�7(�z�9��T���ڑp��A4���ܻE:ꟛ�9*���^�Y�Q�@:�&��(�Č�uW['����bѢ�D٤����-RB�P�ec�"��F���D�;	Ԯ<��n��o�q�xN��i�?/]�H�JG�x�^�JΏ�GG��g�5!�ѻ�#���.�@�4%Y��ᡝ.�qYܙ�;ڎP�q���]Nh��Gbb�7ϛ���X�1)%D�����F�{�A�B��
mV�ޛ)�bP?�x�y��z~�r:;����ఇ�����9��o9��CP��Š�NjU����zءk5ϔN�N������I��91��@�w�=96�ԣF��,d��+H�,pc�ͳ4t���es hx�tA�v~H���}��o� %�o+D#/hp/���?�}E�y2%��8dcJ�p`�;A��j��~3f������;����#�sO0~��t@�G������g��Xȶ�)߷��]����+�bdEkB�F#p`E��H\	�s��P�����fnQh<z�؀��)�,�=p HrwMn+����,�A����Y�!
�s��(<)#�d\�00�R�� "r���	1j@��;�NםĂhǴ��B��Vɬ(k�#�n؉��0�@CXZ �6���)w�X�w!K�.����_4N�8����
��p������P�kz"�	_
6����3Nft�HGۤ��^��c��^� ��ޯ��yt8G��v��$g�N{�*�%��2�)Nxޛ�ZP�*��NtO��^�Q��ԡ��y���D6b�{�Fyx@=�@�SI�=�_jd���F������@t�z��)l9���'Ο��EpH��n:=f��3�-4��M�T� ������"=;������d�o�Da��'FA�CdF!��:`k6�k X����_�I��Q��n,�ЮoѯO 4s��xn���r.��Y+h�x5B����&�s�5ȸ7�v٪cy��͜=�/#����z� W����|�^��	���<A��b0C���h����1=�\ׄ�y5�� ���`t�:5�O b{�D�&G-
)B'G;a!q4!T���
h�iX��k{���tV��{��$��\�xF�7va��+t��Z�ڤQ}�8U�IG*-S�j���y=��-b�id��%�b}s��XW.2�E�3W��s���$�PBF�U��SC��}�0���	�-FD1$qj+T�)9�=
�
A+��*tWh�>������
����VW��N�fA�z�C9O���]p���e���|�fԧ����tgT���9���;M���<(N�G�55	��
��]-�Ĉ^�&1�)EL�Dњڷ�l�Wo��HS*(KO�yt��ڝ��wH���<�Q��&'�z+�&>)�ߟ�#���ǽϛ���(�w#M�@.s4Gؓ������py|��z���l� RP������k!
8�rPq����RS�s �U�
��hJ����j}��?���*Z�W�.�O��o�.O߷>}�(׏�킢�	d]���@OڄP����s�ݠ�r���<G�V������g��2�q B)%����{>�q|�[ͯL8s��Ul�<�4�À���yiFO��D�q�}��Du��f���"A����r�n��H�[���fs��@!Ik� 44t]mp�Ѣ��u�]�MȨ����!�<&e*�z>��i����P�4"р�vxʹ�,���I�aMF[K��;���P��E���W�w�����,��<#R�VPF$������1ʾ�
�T���ۄP�t��07���DԻ�2M��=e��]��5A�������C�"
[ZD<�o�_Nk:��z
�^�ItP�N�a�lvH�>뽓5�Z�t��K��:�x��p�:�Ml�촻(Ӳ����cG:�lq����>)T���Z�M/��8h2��b]4�^g=��2�~[4O�+|Џ�1N:���m��D�����P�޻��/j]tvcT]+���9I"���VR����Q��y��'�����z���F���9�j�5��DG���r~�������J�������
п�v������/���|���#Oo>�O��{��\��1]ߞt{���!?o��ʽ����	e����JC;A}��d3��l���1'�߇[����`H�,o{�Ȁ��������.7��mD�?MCvR9|�Ip#�D�uD
t!�"4)7$��B�S,Άf=�Pꝵx��3��#?���ל��.�:��P.<��g����x�#SᏑM�$@��F�*c����pnsf"6�X�P(����!.{��e�t�7�XC~f��x)Z�����M��Em�n�X�9E=��n[��@��&���J�����1ǟ��,Pm&�����
*}@���-p����9��v�������[���_FE�+�À�]����g�d3�:)�"���y��^#����0�Z�Z3���\R1��d.�j�E߼�4�ra)�����o��^b����9���wA�|����Y�3}<��=s�ߥ�i��DRc�)z�U�I����M
�U(���RO�`׷����_h���'P�`��?�����^���?�]�K�~��#���~Z#|�aŶ��?�_�[��7��������^�>���?��$_���p��(g[t�JW-:dT�igz�j��P-?`�K\s:D:%J�~�� @s�Y�=	�,x���=��.%��Z|!��Z:@شwʪ��4os��qx}	��!�b9�%��Ӂ����pbn!�o�5kj��2�PU�����\�^kb�1$����J�2?���
w��� e����	�D�����JQPͰ����/��>9�QB��?�������qRV��m�''���K�3�{_��!w1��>vM,:�8:	��w.�`f�zZ���(�1'�@��߼����%|���i7�V
��l�:�/�>^3��<H���w�}����uaAAcڳdb0N��HT!N�j�����y���T�r��ۿD������3R]����P��	�vW�����t�}��x��HV��4�-��<G���B�dQ<��� C�T�ڌ���O�zF==��G�ԟ�֪��
c9�!T�i������_�����<~�Ͼz�����?����+��?���կ�4������K?�7��ͯ}ܶ�����ۼ<�~��ў>�q}��UY���+�zV=�v���#y��R۫�{%uFRb�.S|qPǩ���L�(���R�7x'EGo\�3��Ľ',)^��A�4������?��0#����'�><ę�j {��k�ZYJ�yTmK8G����#��_R�dO�s.ܓ��>v�vݝyE�&A�؝�a�͞�DCJ9�9� !B�ځցnSkuR�N�6�e�������g4�w*�1��:���s��FP�mP0��1B�?o��I�I_P�Ӗ�$t/�p���<�����;��);�r�ɀ�:	���>rYC��wN�S�0���d@���,C/��;�=䥵8f���N���������X*�3��QWq*b���hR"����r� U(�	�t�����g�j��7r��h3l�Nr�c�rf�ˆt�uLR�i�{�R��a�u�_��O2���	�d�p�5���Ƙ���h=2L����IQ���R�����$�QR
e��c��T�����>���_����/�?�����?���|�+);7����#� �ſ�����_�����O��/����^�w[9���>����+X	�W���b5̉5����������z#�7��~􂻇˪�GE��D�����1��~��vH�ה����<�^��=�r�w�E�!��$�
t��	K��N4"t�KAQ/|ӽl�!Mo_=R�� ��qs:�PC�h�fg�%�~�8���N��1H��r�y	3�-�ށ�['�ݢJ�A�*�l�h�!@CF��Sňt�q�7�g��
���& ��4�����������'�3�^����2��=�]�m�IRd�S�V<\|N�`ϑa�aIMݟ3��mSq�F���#��_��:ݿ�[߿�������Y�����[f���t��QjEe���8�1��
F����vl���z:�>,(�RC�qJ�L9��{�1�#苑
Ǻ1����9�#�	�߳=G�!��|G��K{�x���Π���.RǄPN�G����z6�}yQM?��68��I��� ?���ß{x��\�����?����s?�����!P|� _/��z�����	|�w��_���+�o�r+��=���w^��+t�@H�	mӺ!*��<mB��#��iCW5�[tp/��ţUo���A2��������U�����=?z�zI�T����9�Y�~�D=BG@�{2�8����k��c�D1��#:�< 7��6�x��X;}�1�P���L�]Q�x����`lL������v�ݻX5/x�hV��a�l��vJD��T� >�G�cIk�h��O�R <ߋ��d/Ϸr��}q�������^2F�Z�k�6�m��H�v>���=�4VJ���HE���b�tPPa��7�oQCA��Hόvɻ�à�\D�<>�Z��c�{����0��ϰ����;�\����E��pH���-�T|0P�`��������"��(��z�R�sJ��C���Ngи�X��71��ɩ��O�+��h�=Y���Vd�&��S����X��;��Y��H�I�(�lQ���=����јhSV���a=?��W����?��_����ӫ������F|�t�t�h�?�=?Uŵ5|���6�����>���~G�X�w���կĶ�d�C�LΛ�����:S٪� ����*�A׌����#�q[ݗr�A�q��T�z�."�D��������g{љ�`%77�! ��g*��@M�N1a2V.2o�ݴ��ˉD��p�V�V�A�d;A�nS�`����!��Z�_O{�y��c^j^�DFQ�H���2W7\�w�</����I����&m]�6��AA�^͂�;�TLn5�$�S! ��1�jjSqGGG�����ar�g��m�F%���D�><7+�w$��#���9
��@�wV�6�]@�ԛU�������耘�,�ؔ@�Iǉlx�*l���a�����(��{���ؚ4���iy)ʞ��^>���P�{	���QkHf�[�>.ڊt��Jݜ���Ή����h� ��S=���H�`3$���J�6�E ���U!?,#�iݰ�!ϒN�4��f�?κ�^ڎ���{~�^�A����(�?�t<�!r�g��R� m�Z�^�zBYΞ)٩Hb�D�E��@B����������|��_�G��~�7�r}�^��}�/��~���M|��}<��gN�����imu�=�#��U�\�a0*l�}�T���!��G�0Ըɡ���xV����S�%����g�i���}�����͓��&6���!�=�Y�� ���FPAǆ�q(��S4�����+� mP���Qu���tX�H@���M�S��^�/�qWF�T��k�6ѯ�.F��;;6���#�04��fp)˾�ɨ���)�|��� ]��"�ֽ`�L
铧̓gޢ?tLY$Uk%��*@&�R����U3P��$^�T¡�z�D�w��"	�EgErV��x��;�{oc�-��c�Pp_�r�A@��>nq�� �'C�O�r��6�3�f �d["I�:l����P���m��MD7G��r�sQ�X�{2zgÑ�P��Nʔ�E���\_�\o�z�A2�"h�H�1�Z@�T���t����`ش̲�.g+]�j�iT�q�Q �BNe�����6��Q?�U�F6�w�o6&�����nF/&�7������I��j2":�Bs$��#C�d���*�:�Ƞ��drp�����M�^���(�>�X��>>sy�3�S���4z�S��s?��O�N���������x��=��c�W��~����O���\��W���r�����y�j������
�
mH�ԃ3zuJ��F���3���guzg ��}��~^͕�Tޥ�0�;>Q�z"��X���z�ҧL�� ��3΂,��{��� ��I��	�n�P��5�<N�r��i�������Jґ[rJ�=Vrxw��dx.{�~�y?y��c�^��έ_�R�������hTk'gDa\!��;=�˳�Agi�K^�;d�Nt��h�`��뽧LmNw+�����)g��Ϯ�5 Z��Q��S�;�4�F���Ƶ���]^�������V�Qйo���:�����c�%Ekf8���:0�Z��UQj�
�@�@��6���v���zGa��m��X+T�M^�3;�KIG���ڼ��b�^Xs�ĬD�ǹدW~���@��ⵌ=$/��;!�x�ՑU��F�b]I��Ǜ�Z�r��j���>l�-2G�������3��������}"����o�������2�-�x|ϯ�!|��� ������WUdٸ�����#6Q��bסh}��	�ä\@� j4��͌�X�{0����ctH�����f�Q����i�C�@�(�N0��_��"t=ٷ�����;�����KE�� uQi,P#��37��(��n�tB(�Nc�q����a�윪���)O���Sۣ����@X�U������
��XUU��)�9�V�*���v ���1a�����r��1R���	��c6�#�^4�p}�Kk�N�Df���zWE��[��JD`�AHs�QM|�ji�@��@�����%'�@�cO4O�y�x��������I��M��ұ��]4�b�,�H>\J�_b�;--'�DQ����k  {�IDAT8�)�R�S#��Cl�+��ST���/��h�q�bOj����9ǥ�Ss�z"�'�4ޕϹ���7` �w4���8G�8�� �re;W�bRr&f�*��F/vV����N��<6������?�����k������mt�r�_��?@߮_xx�ST7��V�'��p䛍9Ǽ��R�%�bԆ��)⽩]�Ź�i_��z��W\�{���qϻ���a=K��6����@�"7:���1�wy�c�v�#���&�3��Wv�u/�Q�wQt	%�)���ب�B�J��ή}�qǺL`��JhΔv�&ϯ��cjRBw��U�*��x
%j(L2ܥ�<�Maμ_���@Wc ��0h2�S"�I�Q�%t/זb�t�EI�@��|qW��䱘c��ˆ9�mޓ����	�4t�
��$�ĊW���%�G�~��ü�H�O���/�GBn0^�,��|�
H��L�R��^�� r��·w=���_��@�	����G'��='�G.(������|P�U�;�S��hC���lNz��/�����ebv2�{Mg����%�ِ�8�i����^�(�=ݞ�@����J�U��4lV\H�-�DF�����j������������|u�����
������xz|�p��t�~͏�ķ$����6��/���/�g?�����&��j�簾)��,���
���c���b��4�0�+ȩ?4�Jx`��|w���<F�d���� �[{4u��߇�C�d;4q��q7帱�*Niy�yVA����ޕlֽ ],Ci̠3�AL���o����ۜԢ:_����d�W��*�{51[E�k���H�n%�J8~�
��ٽ�euF-���;<�SC�<�C���f7�6'R%�,|�k0.�r�i����������;<�q���A��=��\H�U���p��D���I��=:'���b��Ɂ����V�E��`C����隍�|��*����,�Ѱ�2F��ɽ����l��B�ڣE�@(5�A�Xo�9U�K1�7��Ҭ�X��f�
pq�ݲ��s�{Z{t���<�[��T~+Ծ���:�*��)z��0�]��<�G0���L����cׇ��	�щD�R*J9���@��zYD9�����[ey���������g������5����: h|ק��?�������"�A~�n0���
1:��; �������ӌ��Zl�o摂�{��+na������`�o�1U;�Ӝ���=e/Գj���A7�(#�.^d����o��
�(^�G> ]�Ό�f�}b�QL#��.0x�&�tvL�6�ca�U��W������{J�4��R�U":1�k�쎟&��8�e�͊����[�N�] ���3i9���F�` ;�y�q�#"�=�̕D��f85��ǘ�(���Qr�q�*J%&�IՊ�^|L��=�3�אq�7�ywgX�����p�a�c�8���E�����7f����,�WW����[9�/�ɼ{Q�;�;cp���D�y{�:�f����ާ*��]�Jo��r#V�JN�$-)[}��5а���IF�]�e܋��2q�8GGv��;�:˰��n�MQ����$"�`�0�׎.�;��ہDEJT��#���c�ƭOlF��+�<������?����/������2���;6���_���ÿ��g�y����/����/��� ��[���n���;�
)S���O�WOաMσ���S�ӵ$�o�ncX|
>�[�v����4���k�홆3��}�0�&�ɫ���A��D�M�)G�&��� � �^R6#���͍	[4�<r�0c� ���R�ESTu@�3����r[�*�m�@̎��E�J����/� ���{��S5�
�ym��z�X7�eSl�8�Elڔ�s�>�`�t�P��Lh
d�vvx��1�]~g������(��HQ�v'�H��{zN�Z3�9���c'�N�t+�$o�;����[b��YC�l
]!w|�o���Ao����Qp_OS�_P9�5's������*�'�5
̣�h�+�!�8�����hZ�:����#��Uw`C�H����츼q)�,�H�:���,�Z�@�	���������"ք�����HA�� ��i��ApG6��ɩO1p���/a�o���>��|�����F�μ�=:�����~�ٿF�0� �G�LՌy�Pf(��� �������x9�������������oů��t ���u��O�5�3�������|��������i�=]�������w�^�X+B����"om3�늫#��ywod��n����6�n>襛�`�1db��,U�}��w;�<[#x(�P�0�,������Z�`!RXn��qH|`��7��1����y�~������aW�E*��
M�k��(����S�,��o
��U} ��}�<�x�PW������]Ѥ�ڀ��X�b�ag��9ڔ����V�nF*����g%�:9�Fu,�L�0�2�~�4)�5�Cs��(��i�]i�<b�| ��UG@ҽ���p����;��m��~~U�����BLA�������X��n������	Zރ�����,}�M9|�������򏜴)�a��m���Q�����WdUQ/3�C��ԋ��za����R@��h�B)F�-�љ|��*qw��9��V]L�ȟ���%Qk�"�E�a��aTp�!}N� L;YO��|sDC�C2h��ٹGd��=��I�x"�ʌk��Ȁ�i�*o���T�����&tdgj������\�d�I�sDK�
*g���W����㯽y�������S?��ߚ޻��t ����I���/��_��^_}��U�~�_�����~-�3( @�%��P�[�3d�=g�\��3
�o�������s��O,��zs�[O	��{��0�?
����P��#<� 3�1(��p�`���I��X�&O���,D6Ioҝ��P�}�G��1m�]�
fk$�N��v��0��\��
q�|#�V��Q���5!Wx2�k��L9l,YQk���l�"�BCfW���5vG-��l�Ս(ᥢ���A��Ĩ@]�rXP0s�W������Bچ�6������98�Ű��M��DS�v��d|���U¹p4ϨO]n��6G/<SzG�4��	�6n�!��3��.X��9�r��y��9�Jٙ���s�����_�d�����LPf�m�n��$�N�n=r'���L�i�;�2�,�����PD�/�^�og������g}.�-��D�3u/�6 ��\�_�������8p��r�B8��s
4	�KB�\�����@��BkW|�=~%�_�A�����i�>>�z�~���ڷ�E*�hW�r|�C�p�[�l-]�S�4ra�M��%�� �����_��ѻ�'ŋJ��1G���hg2��pX�]�4a�-:+����d�[S���ם��G.6�;����fo�b��x�*�l4�4w|F N���1Q�qM#g�{Cv�i�9uq#u�a���Ju���s� �֦�4�&�8-+[�%MF�����9�4���`�{�d3���c�(����>�W�v��9��c��hh�d&��7��"5!IC��K&�Q�x��{�����WH_}���]�Ќ�(y$b͐g���
��Օ|����2Ҍv� ��?���O�i���|)Ĳs��u����ñ�~alw�{�|^8uq��z�y�u�̗��N4e�32(�w�sv]Y��������dp{q��T�Ӻ�3�)����n�C١g��s}  L�䨲�C���c��=��j=�=����3W���r�����hCگ��5i%O��,B�ji�@/�<UPY@��%�ğ�������?��}������Wl�����	�����u�ׇ?V��GD�?�}��RVXn�X����
g�S��@�����2�\a�1HV�1�b2�����f8e�!_��'/�F��3�/�r�����0�{��q�C:���+��tj�ϝ�$�1�{��V|r�PA��K�{���s-w��M��)��v(T��鵻H��7 �{�A\3���W1�T<�#�hB�n��*X{8#�7�7 p�0R�ժ��͝5F���Z��6�@La�$����|�Sq20z�w
K��x��/&��[B��Q0����:����E�w���A�
��q��������<:K�;hθ �������':���n�#�Y��Ζ�I����$RK������
=����qxtȧ�o���N�6!u4Г�+�>�<.x_�0���*�Y�>S�:�SD�:r� �3��u\�/F��pz�d�k\�����B �(�0���V�N㭺S�g��wQ񌀌b9�qu�`���X*��<��l�K)V��S(_jI>:/A�GC}SH���L�1�l��r�3���d�{��4q=e1����zz�7���w���*n+���ǯ�A����o�~��տ���U�?ޅ~-�P"��&�/hޝ�r������&43V4��!�՝�=�$�6yn���/F(�{��7��S�������!�IHTSk4�;���t}@v�?�Z`2�Sn��L���W�P��8Eͨ����ɘ'�8�k0I������&�0b����o����Ús�1�Ȯ�5+��lk�h�6�"�+�� K:�F���x�G�~�UCl;u&I����k�0)���0\�p ����0���㛭P����E�� +{��ۮ^���.9=�&�m6��2-|߅r9L$��fA��ơP T�T����؛���4�Y�u�L�q*�B8��i�fu����M L�_�C���ʜk�`,3���X��k���
P27-6��{����H^�y�F�Z�bC����v���G,���+1���{6DT\�u��=C[�st8���r�3Z
	�N.���ʭ�����M������K�D;��{/��C>]�a�r�	J6�	��i�+�h9	��_ZN��'*�&賟ů��Wՠ�����.�-��C�����(~����R�ђ��&��w̥���/���z�ɽ�c$"�㩴�@2�x���杇IJ<.9`�Y�)'�vR��0��#
�C$ޮ�0r�$�D-��3�N,b�U�H{4~�O�"�%�n4��Eq�\�q��~U��ppr�o}��aBe��?����؋+����(������ڰ�-&V��r1Gd)x��qk�W�ϝ���$�]��m�������}d��es}����!�{e�;9
���'��f�U���]G���b�c*�$=2��>�H��n�
�hv5ǈ�#^r�tΜ�J6�$`q�������~��ŴV��LeZ*����ϔ��\��>g�u������~�F��n��A� ˺T:zQHS�1�ǝʜe��<U`yx���3tk�ۆm���,��U]�D�&�B$�Hh�Y6�Ο�p�����0���a����i'>:㳃�x_d�_�{�{�a�{��Q}��x�?�ʲ���.��A/���߹���?\N�oן����oů��Wݠ���������Y��]P�$��D�?g�1M�a���8հ�.��{���J�lƬǴ��]KD�M�"��#e�	��1M�{����&%�Gh��w���(�1}���# .3�6��&s)Ōs�9݅&�k�H����gT�֬&DV.��.�E:-hq�B��P����Ǵ�4��k2T����fx=����鸏��4gu�$��m?} �	P�S�^g���	�W@�2�
+����=#�
����yDP�R
ά`w�p�3�	�GdtB��l�D���\���A���1�>R���ϕ:�jr��̋&�к4wX:������tt:�8���D�u��FDsxJ���ȏ��N�i`ҹ���D3�����!ս1pٍ�m��@���J�o �N1j-�`k���H=΃�cbdt�E�O7d=}L�����e2�2�"JE}�^�`���a]W�m��A���;�j�iL�.���6��C��G�2��LE�CC����ռM�t�3ՙ�{s�s����`�p̵N�3~T4�h����X��\+J=��
.%i����s� ��-���x�������~ ��R~��_u� �����������k��_����?�x�qR��k��Gi�*�2/�Dl�='�f��ȹ�\9kU
���{��vo66/<�1�2({
i��̚q�S&��( �)�3 ��Ǜ��W4 �h��52R��iE*��V�,��x�|����v�*CdC#�(^�U�bɫ�TT<�{��%��3m|��Ӄ|�Bw�aIX."]�[��k��R�F�!9U��*[YA��nX�׉!ڰu`�*��@��nO�������(�8~�Lv����פ�8-��2�Hh�ް@_�p�$��#X���L���hҊ���{��:��3�RW�:�^=K �v�`m�.��P�(*0s� 2N�
��6�� ���ZI ���/ � ��3P�"͇	�!DP-���Kq�:E��@]�~�#�:���Oy�TA8{���ADܐ�jB�����������9l�AM����m-�샙l��2N,�4�|ƹT@�*ضo`�Zh�X�:d�D���r��a���t��1|�����";*?f�a���49y�m��&v�Y&�<��0�k�0�i\��/o5 ��h�>Ӝ�*g�ogCP�,8�k���Љ�"P��]���������~��X: ����C���_�y�c�友�E;��唹F��� e��q1���DKC� �Vc�#~�a���|���O_E�FD��VJ�N��d�%Z��]W)�B?�4X�|��G�Qe�H����[F^Z::8�EYD�u�C�ڰ�����xd1R9�a�#q��Zs싺�{Qّ��P
7�.p�3�#k���X�>9zc���`��Fh�]���J�B|r.uW�$t�*������XQ����<H~Vb���
�m���;B�{��X����n�ۺO����A����ށ��n��)v w�B�
�qD���O��2�)1�����y�d�����`�(��4u��[.�-{�����{��i���	Q��A΢���>�&�;�x]�� -Y ��y�Ul��9�x
ʉp~�@ߜ �P"�z�Њ�4gtv�ޱ^�^ϗd�d,�ps�����)9����mi6DՈ�DB�vw�x�:`�ӵ���A��NS*��I��T��՟g����W��|�������[}�c3���G�o~[oW>=�;��O�<��.`�@ڲb��\\�,�I1
T
bXTl^���{�I��}�}�j�W<\�	uŉ>4+M��<�'�NcL�����[�����Üǁ	UESͶg��t�ϡ֘�dF����}F�k۰��E,LL���$�{��"��%z�^���zג�R��,��w���7�7F�7Ի#(��fQP�CiT��]
Val=R4
5u�ϙ��nl>%pF\c�S�hI�����A,5��&Y�:�w����g4�_rA���&��)c#
(j���~B�BnU �'}��+h�5�ϛ�C�=�h����8�2v[62a��됋H��C7�dv��|�;������t��}D�"á�b7�m�cFa�h�ʔ
`z����j�2��V=�T���S��a���l&K1��A�ay� }�F�$�e���
�*�&��l�~�!/K��3�я"w��J�o��_H@�df�AȊ8M'�H�x��dDȔ����`^��Xu;U�؋s>?QY��e9��'�y=��[�����͠������[���|��_��?����h򛣚�,�H&�y|�8�������mT9{!���a�^z����5�>
M�OR��ÃӃڑ0�4$� ��wJ�	���!��5����hD��������n�& !�ްiCG�
�P��h�
P�y@����[z쭝+@�e������N���~��P*�A�ɫ�cm�`E�5�����4��	:�D4��{�<�%���C�����m��@��;>���V|(�a����A{eA�3�'�'�L�b"r���ioZ�����!�{�F��i��qo�-}���_/����� l�p�>.�f�,mAP$q܍�X@.�RЉ�!�)b��О}��m���8lf%��sFn+F@�H��j{8ڨy�(�L1����pPF��B�` zoh���0�8���[CW-'�v�b��+zP��|^�u��8[qQ{�>,�;�������!�����R#����SR:Dn�sd�dx�z'ӝ�|9� "�2p��?�/��G�\O����p�ys��'����[�/�D���_y̻���x>�}�����|�+�+Z���B L�ژUt��L�����OPr�.�|�DD��c6�s�����D��y�!�Js.*%���V�^\6yʉ���3v/Sqe�0Y�Td-�/����sLe�v�N6{%:�����������=��ð�2��:�Oާ�̊0�b2�|�~?����1c�P��l]�|��(����1��i��S��O5;��Q��t��r�n8#��2��fx��9����-u/Y�]�����Um���~ؕ|�l�$1��C�Y	��nn��}�jv��\/���6��G�
ι�|���v�����ɨz?�,v5���-�߀9'>x�<�Ǿ�\�Y>��ǽ����f��^������3Mn8#_?��TQ,@�(ݣ\G���G!͌��	��n��;�Q����'uQl��m�W�$�(��Tf��<NAԋ��^�i �K^i����`6��{�(�& ��YS̓O�@*���{�x
�E&Ƽ, -P��ǝ��ᖿS��������o������oK���?v�N����i\���v~x�����.��$Ҡ�-g�N!�YU��b�ȹ�(�k�����!�����t��A�ȫ��j��T1���A�|`:�r����3^E�k���.����95#�(��n����Ѐ�=�ǀ��4/�i@o�l��t3Ӥ��+��PeT����Z���En�q�V��,�^5�mJW��������v9�a�
��veFA�O�o/�u[ �ص��W�(�Xv�R���N]�n��V�DL(T�(J`�1��=m�\X�S�^x����*���eT��
j�6�C�(h���u�O���Y�w���Wˡ���[)!��A��¹�1�ƴ���>�=�Z�M�M�֗)!�8;S�|�U�Wh�o9$�gG���丅�G^����"룎�}2��@+�,�
��7HkPQp	G�u�s�
��q�ܮ!	�X*N$t*���7x{�#u����N!�����{<��#'՘6�h@�����h�c��	.��֙�uǣŞK��}ܷ�Ǎ����l޹}���R߂�O=��}��	[�~[r��<�����#?U�?�����l�[A�G՛��Y��A@L��,֩Vй@�8k
AVC�Lw�N�&{�b��ｲ���D���}z���y��!ǎ�v�lv �Хa��U�F��Ū��U���A#���A��|bu~o"g5�@EA�>w36_}@��f4��K
��`�e84�:�Z_��G��'PTG@��%VQ`mT�O�v�(�4��U�u�7��u$7h0.t�&7���\��O�/���o���{��l��B�ʊ�4ǅ�>X��^N�I�$"��HC$R/�SD�ٹl��G����������k��bmˮ��9��{�s�[-�"�H�D�UC�ɆaAz�yȋ���!yH� ���(q�8�b;Aذ��U9��P��I�H�b'���朽ךs�<�1�Z��[
`K��<>�X��=g��ךk���#yj��$�$�@�:���z�A�·�ȑ�B�y�E{�k�ܷ%OpB�m@�w�.��F�o���p�V���3���	�պ��F�ͯO��٢k���S��v5f򜮨~>$g[#0����� $���D�}A���A���A>g�{���1VD�{~�x͊=�{�����܈b�8h=B����o�C�U`۬o_�~-����jΞ[�]o��X�y+����ސR�hO^���������`\���ɔ�8�Q�)�;��	H�o����{�ӧ�o��]���|St ��7����3 �oӜ�
R��H�(�S��Y�蕚�b� � ��T�+G�d�z�����=���V��z������jk�ppxԶ�0�ȫo��G��Ͻ������w@e�,3N����$�W�A�c��X���z��+��
ؼy�H��!�[En;&ɦ@��gߝ׼��X���#$�֚���RoTo# �@�R����t�����r���㄄Rp�ͨ�!�����w}u�n��:+�C9`H��f�k3C ��isŔ*v%!�l&��6�m���ka;4®`�yd]�����i��{����f5�lMW�Yĵ��lb�$�*6^9ۺ;)�xBZ���Pb2�%���#]��=���"���z�a�x{ UF��q��+t}���ovK���%qփ��f�0��QN�V���f*�O��x�{m���	�#�� ���
���~�����Gћ��=�f�(�h��RF��(�6^C�" mH�.*eE��K�ǹ�:^�E�y�<�=�/�ނ�̣R^�У�ϟE*]gk��)�g��j��P�:�ڈ�wAu���̄�9�~�j��kZ�,h�lmg�3BU�{��Ϙ=gkQD�He�i�\~���'�����w>�g�}��i���>�/��G@��w���P����.���z�S��Y����u=�H6�ΊX�0�vV\u�}����<?�e�w6^� �J�uz�6�z3\�Tp�`�����-3
���e[DK���n،��o0�/t��c,vX�C-؜-����0�����*�9��}ޣ!�P�t���(��F8�-�ko_�ń#���s]�k(UsS����r�ن��D��K]���_��[r�(9��q���ѥD�P����F�i�;z���|�*X[nVw{=�5Jg�~nܗǴP����9��nc+.,#>$��Q��d�&���0[�^��0�.����Z���z{�z$B7+���{?��}��v�z�o<�}�=FNx�����e�_���>�U�~v=��Y�Y��X��u��ݼ����
²4�f������V�Zdu�d�9��mޢ��kŸ*ԣ}ԍ醡O��̍��j��k@�w�U���ԪEs�߭׼?����w��FPO�l?��_�fx�{�������Y��\���v?��5���r�4��i`�sB�T���rE\����3��^A�w�,�i: ��=«_�,T��'�?)ҾhO[Q�چ,��7��g�<E�Y��U��C]�4vcn���l-��}}�R������(W�X�]��������;�y�ɍ|��y�U�4,*�;���O[�<���������V=��&���Ekn^-���H�ҲjcCoN���_,��ݾ0ڒ t�|D4ܪ�n�9v/�z���Y%�����Bk����o���I�T��T��^������HDP&h�=8B�q���=�%+JR��:�=i�д�Z�u}���Sg:c���\�՛ܬS=�����ޓ�C��{Y��Mz���6�³]裙�7_�����ڸXxT�,"▛�3?�ܘ	�@��Wj���q����^�g�7���5�H��;7��Y��lk_n@m�W�V�st���[��lv�8X�c�B�E� eF{M�JFJӴ�߿��m��*���<f,}~b�״{���o����.(�'���c�����v�G~�����V#���Z+�#\]5o�Lv�����o�O�<����Fa�����ϕ�U������a�y�C�'��G��l��c���x�\�8.)��!�ݟ���r�Dx����7�o� ��Kb�)�ť��B�M���KJ��b�m]25 ���=n��ᦛ<2%h�X;7�{����z�ga��p�ж2`�������g���o'M�}�\a���ϓV}O�uS%W�S�!�	��u�3?[�*
ۃ��{*`�OC4�_y����Ln�Kkr��Mα�m�Ms	SHm��,Xj���ൄ&��ӱ��0"��X�p=/ :��t�ߡ�5�	#wj��ke�v}�C���A���{c} �����%�b��}z�iW]\0����#x>���8YΝ�W����_�
uc̨�H��R�Y��RJ�G�W�
�q���n��|^-���5���Y-C_���nK����@��F�˳N�B�aw��~�i9a96��K���r��M�K��!�P�I̦��Ƙ"/2�բ-�V��Ix����MM�#������~zc♉��h��������g��r�#�����CΞ�.=@�3M����<LV߰F����)�a�t�"m�P.P.@��\�Ly��D�"��/~�L���s�~/���W..���|/(�����]��f�Y=���*��@#�8���	�=�)��B}�w���r�k�n|��}@ȣ}���gS�zhY�Ko66�����7ӋlN�{�je���N�Q��g>ސ/d5˔i��>�9<��_�{M�����u���h���m��!H���������W&_)J���$����1�<mk�r�f�������6,�۠ɼI"/ SZ7]d��Z?pv��3	_�{V7#���k��L]o�Y��_�.Ȅ��EX7G����K��u-'P��z�^�LxUIܖH�z�����t���=�n����m�����=�k����'^�@���0�G��|�v����������	*e�[�����E���H���њ��\��׼������X�_	�d��"�Z+겠-ER����,�ݣtM\�P��2_��l"�g_�\�>��Pd�c"q끎��nu���o���)o�k�M�M��`�������|�l�7j�!YtJ�s�f|vA�Jy�4�/���SϽ�C�����|�t ���_��G�A�����(�zഘ"\J�Ruo|-8�n3�(���77����c�<��^�&\���<~jͷ��Ϛ
�)������f�=yȳ���U]�%lg�w���ga%�l�=mb���j���3dcWW/�7勈��9��=���������3��[�g5:��7�����&�������P\����4����I�&�j��
[�Xl΃E:�0ڼ�-9@M#���X`sK*�0�i�R�z��PzT�_��d�w��7�n
v#�~�V�C���M�ϥ�V�<���C�쇆w$���<c�W[�q}:6�v/"�?�̣m
C��("hU�se���M�E�?���r�����A|�N��ͪ�a\oWjԺ
ed����3d�|6�EE��N�,f�]a������۸
_��kDz����D梣���@��'BK�^�]W�j�ٵy$}#�ؿ��n�i���3}ܬm���&�cݳ���g`Ѝ��Jgn�*�k����f�|m�I/R4�=G�NR��5ev�JY���1󟑺,x�xCt x��n�W��֝�_l�?B���Ԓ}�J�jT=d�'J�����x3e�B��V��|�&��_��^
�}H������i� ������"7s�����p-�9�|{��Z��Y%_J#�:z@�?$��0�����f����>�	�L��>Jz>���B���M��>�_�q�}
��ʞ�2�M��[n�}F^�?��@�!>DVA���6<8Uk�iu��矂{�m��Ms�uH�Zn�y�O�d1O!%7~�`Y��%�A�庯Q� ������#}6A/�qf��C��=��HX�Fī(�y�D���tow�3t���&lFC����Ev4fh���u��ߪ�m�3�?0�זM��Q=��~hml��8������0Z6ѡGX��7���)�G�k��v��+֐��>� N
i3>|t�̋�f9����Sf{����Jƴ+���n�c�įA����z�R��lv'���t8E��&����$o����u��{��u����M�v�e�Wt�@m��9�F��>vw�l����ꐽ#�[��7�Mjek��1�}
�$�dav�l9���ze.����OL��J}C�s�<��r�í8��+m��?���-�Ia���B6�O���ΐ�M��%��@h��5�|�w[�لf�-����X�HCLHc���o������r���s�Y��7� �'����������SF/��;��=�N}������-z��ՠ;*��%��9�6 ����6*N������~h�5���	��W�ԧV��GkU�a�+k�lc��#2� -�tif��x����z���!%F&��8�A03�ZaS�D�B�s6A��@MAd��T�\UܛOk��<�m�t�����J�m*s����2dh��h��6�:�B%{'�goS�T�*ZO>1-C�$s���5�	=F�%������6
�Z�Z)�SF˄�Pջ�� q�skuYX�ad���=q�#�	
~P�z��3b���:[���{;�y2��+Z�F��$���X�Ao��{]�� �vrJ�=�������z�5���x��x<b>�����+�8y�G��� �12��`=�b����5�2j~d�Dg��x��Nz���gz�C�i�fk���b�]������������筱�N������d�̉2ɟ儔
R�����"����o<��|����;Пx����_���~A��~��OQ*,O��U�BR>�F�@�!vb��	D �E���܆47��o���t�����ۙg?5o�0��C�����zcaZ�N�j_��H`ZC�}ZQ����=�&�<f}k���N���ڇ���TLrec���C��/����ԕ˺��zЯy��
^�`���x�����͙�ޅ��U@X@X�z�-�i��it�{���[x��'p���W_�7�/��M%7�T�z��4�HlmhW��hk����GPl�L;��k�m�%�s����d\�����c�;7s�7�)�����:"c=}3fx{=��;�{h*eU�+�k�0u��`�(�'CϿ7bHJ.����5��Eic8Co�Y���q���7��*{��z�;{�d��ߌv��H�l-z��GkЍo�����l3�N�������e�jg.�i���=/��`'3��b��p%QL%Ck#ےim���0��n�9=���y�wQ���=�M%r��O?����
���f��MQܸ�����{���#l���*Z���\0�(����iw�}Ⱦ�O+�ߎ/߿8<����F�� ���| ����g�_TF�K��!�4MUN@+X{
=t�d��zA�`���3o��{�#F�����d=T=�=���F�{l� l�@x�E�CD^#�	麐��&^�m����(���7���rֽ��N�,n��fL(�bX���ׁ�z��9�ǉv�m���u�m;�u��%ll���5������긯��Ud�[�j����iͼ�:�q-�)����	/��9|�ޅ{��z>���0��t̨}^u��~��nMVcbՕ�Ȕ�{�
u�YU���VX�f�?K�=�F�_�q��_������D��&xr�zJ^p�Ѵ9���u���:�!xb�iy���:&�	u�u��:�_�M���2���o���#i��g���腐�P��AX�[���	�m�7֪���0�Q�&��Q��8��pA�i��eF[��lW��g��(��
"Eʄ��F�21���*r����tkA�mRghc �_�GS�ۃp���p�t6��fG����it���/n`f�Ƽi�>nO��ɏ���ޒ�t�b�����wNy���@y��g��O���'��[߃E+�}���z���_~
ZT��A������x�Q�
4�9n��U�wk�&����dV*�-����8��G���x�`�/��w?�W\�eUA�}74ȨF�����t�Y�~5r� �������2�V�V���V5 �
�K��bu�B7�9�<w�#�:��6E�g`h�����	����^=�ؔ����j��^��@85�q!4u�X��	kH�H*�:���{����k���]3ж�-5`C�Z7�2�*�&x���\CQ۬��IHv=�m��-kps�b�_3�'�z�lDf��������g���}s뽒�>�+e�J��{�����R�{�j��ŕ��3*%T�ژ��کG䚎��z|�.����c����a,���9��YMVCDקWim�R��@a�x�W|[��M��B� ��6S�Li1�ͷhc��GJDP]��9L���vhˌ��R�s���Aٞ�B7X����u�G���q�Ekg��fxG��yx�-ճ��f����\����T<t�7�~D�3%8�l�R��3(O�����4���|�o_?�C==���{�F��o�Ї��_�9d0���禩�WJ���w/����n%r�m��H�~���J�����5�C��|�M��������}��S{�����џ_�L=L?���44,RQ��I3Fz�ݦ�<�m���S�=D�����2��k��l������::
6�a��<���ڶ��P�m�Mׇy��4�+�[*���Hl.UQxQW}ځnm�T�cePb$m�m�	��V=|�T|�׿���������H���	=�C˶^z��I��g-X�"&��k�u��]|�&1r1��Z+j]�JM���ȑ�����vM�������=rn���u	S�"B3��o5e7%���H+���U��q'+2��`�O�j�N�	���M]�Jb�)eԥA�j�^ϱ���<Ғt���t����p����X��mn��Fȹ�i��=� �E�"k1dJ�a?d^A ������󔐧r�[ſ�Y�����q�����P1����� #��#����������Cfd<N�K72S�Tv`&����/x��|�bv�5��^�{nz�ݠ����"M0�`�j�����c���34����Tn�O�<�-���?�7�7�@�����  ����駾������C�s���N)x���e�2R��̩�=�ښ4p^���V[���<M�[�*�y�f�g?��2��0V��x�iC�f:���E�s�.�L����)������@��w��{n�<��D�^K6�md�c�pcs��yN���I]�$�����i�!�����9�x��=���b��ko@�[��E�S��y�a1�F�bf���W|��	�64졻V�#���޵_���d���є\[���0�h��9N�	���N�!�2�}���2c��?�ߝ��
���{��HI��z$��W}����7S��o=�|ֶ�����]b4�3R. f$ʠ̠\@egJ��%�Ȼ=�T�4�h��]�8T7�1�j�{ȷ#�i���f^���=�d�w=ܲ
	�1Hg�|_��O�Zb#��cE-cm����>AXj��T M�Z�iF��3ي{o�GE�z�E�8c�v�7�n�6��e��I-����#qs��F{J��w`f,�y+ �׽S��=Ӵ���Í�����WV��H7h�!�kO��6վT�#��N�l�N�E��O�2��e9~-�����!�xS�U�׾�19��?W��NH�w�ȥ�"��x{a�p����Zĺn���|r�j������!,}��}cu��o�2�T�6�;�n���1tKY�&�!{��1��]�}zߺ�F��t�*���ER;�H�t����ǯ����z��d�a��x��iW��Hcx��-`�*c�&�b�ns�z$�o�g�{/E$\#>����ЅQ��HIM����+$'�4AZ2O~� ��yM]#�ߌxn���%���L�ځ��ہ�̣��c @�b^�l��1.��cch��}=��&4��ƒD+oB�#��G=t�b��O�Jid�m������>uʫ��C��i�&�T+n%+n圁��){4���g�$��J��kB����ͥ��V�ƃ;�:�J]]w��{�X�?�:�&���=��������O�m�j���*V�����*C�=,�!���*č{��UD��������ݣ��q�=M�\���58.ɚw�iY{���tG����U�-��~���7�O�o~�e���� �il0�C��Ъ��m-r�� {�sB*;P�~�S���� ����x��:П}�{���9 ���r~+��H�X��ԭ4���}�o�@j�#]�^�*$ [KR+�#��W���s�Ƭqtݱ��m�|�6�]�ݲ$�|zYh[=�=��{zQ���f`�{CX��]cX=
�եz�e��i* 5�¾Ag"$����LDA}L����vA��!�Vo��t�2vۤ�o����j���ĭ>�s�����Jk��\,fqO:5+�Y@�����`�083L��&1���e0+r��guU(ߚ=�/��N(d1���WG�1!� �wX��̽���z�ͷ�kߓ�XQ�d�:x����I�H#W޽Y#)���:M̢���t�܈+�$K�d�f�]��D&I^�h9��� M٢>�w-���ugQ��������[�˼`�ŵ��ͫ��}{{���F?n����%��m�4����>��	�s귕��WHպt K���S����TPe��Ċ�#�ہ�Z3!g��tlW}k�Մ,�c��xh^Dp��Hy�Ϙ�)\ER-Z'	@�>Q�ڣ5↳�BU��?��7�������a����^{3D��m#�2ڂ\�������$"�w��;��9�8A�
��r��\ (�N`ڻQ[@y��Ȼ?��?�7�����?�7Ձ �����_�9,K��n�JOr��ip��0���P��NԚ�x!ء�:*K{���G�������c����_���pc����YĲ	k�Yi�L��M�0i�>�O7�77������ɼ,�l{H�7�Q�L�F&��5ܷ�R��0�> �c}����5�%��� 6���m8�/�Nv�j�$~	��A]<a�:s#\WEU=������hJ��-R��y�x>�Ɋ���p�4N���*�f�kǆ��q�'�:G˩E⑏��5�QJ��E��k;������0<�/tv�ֲ�"�PuHޓ��i�l�����'���f�71�:�^��)!!�Y�F�i��^��̮�X.���R�.��*VX^�6�Zl�^X��t�Ϭ�$C}r�n�I-��g�����]��^�W����X�����ӫ\k`�f
p̌R\��>�4�h�v�UR��5ۏjkX*0�Z{V6�͕dG� �_�{���P�u9�I��E���5r3��#�Q���-b7�"]���=j�Q�d��^6��SF*djp�<d�X�4y�������t����w�Agq�����~��K���7~���NzE~�HY���h2�7���rZ=��a�]�o�2�����,k���m�cV9�߬�'76Y�hm.pϫ��Pݶ*�o`�y>���r��e%�y�͐t%� �V�:B�6�I|��9#�y���@N	3^T}x��i; ų�ÓD����5�{�!�l��彘,�^$�)2Ī�uV�M�M� r[<�A�J��`��ŕK������J������@�N	�^��
4��Sww��3�^[/���ӄ=�8��I���Z�:�����������>+�X�����:�^�u[���՝t�+�48�b�/��	>�N���SO�)�&9�5�~h+e0'��m��R�C1��ٌͨ0���z��A��g�y��������@"t��q���z�7�\\��Ū��Vḧ́�ך�_l{�=�$�ު���j\�J���r7������f`8@�V�	)OÐ�V��d3�ن�����u]�P<m)^i,zlp]��v��{Iלޮ�n�l��gA�m+���Kߺt��"������ϻ<��2��	x% R�(�<�ly#�I=�)!BJ�א��s����2�^���A��xS� P���o{���?��~�����|K%��M~W�̓���0��F�Эƞ�j��e{�����@�l��l����]e<�}'H.[�19{xh�gW�z_���
�0�y1��؄�Z�W�ZG����f.���X7��X3#b҂ H�$s�x�i&{���3k��!^?K�ٔi��@���u���:�6a��#^6�x[�sU y�V`n ��y�P������h��=�f���\�b���m��	˲@!�rBNdS����̣*��|�K��]$�W�����f׍y�z�c�S&�������خ_���[���ӱ��f=�����}� aW��e1/�<$��{�잒��!�Ecm�׾�\���@+�2��<	��$���,�v_�쨧��K�6�MX�/����ֵ�][�_;����@�/k�}���~��x�ǟ��vcٌ�_����o�=K e��6�~Y��� MpCI��n͢�Sbp���^Y,(@"F���ڈ��LP�H �)��M�3�،G�{(6?\1�q[�G�H��U�p��9ҿ�h�����8�8��=j�w����!�c��E� W��8O�#�8'(gP��T�<�R�0=��~2��+ǫ{�=���Q�y����~��﨟�9�����Ͽ��?�����"G4,X����C���IA ��۵J�ԇ���R�^/���O�6w��鮘�mB�:�D-�	�.�V>�sQ�Jzh+���R�2]�!�ILloߋglZP?_��IU��b��EO*�����t �4r��mU�g�{}�ȉ�h۞���?��26�5f�!Cү
�MR�Q�Rd�3��n��{���K2V�,��V\^6<)�L��Vۨ�ruh�S �U�d�3 ���խg�!e3D̨i,:��յ���޻�cܧ�g���ՙ��z�F�9��SztC��9z����~���M�A ͞̳�1r�������WkU�|4e@���zw�}-[�;�-���}
��]�2�Ț 9����ģX�0���y�\�|���q�����#i��n?-g��=6�k=��n�z��X��kU���4��"�%'L�	9%;�`�L
挤�T9	@�l�Fk�4r��CY��
z���M�B܈�\�H٣~�������zQ�p��������7�����zU�Yn����n���zU���{�*m�ל���@��(Д�����7�\��mJ{ ����ɟh��}���aqޤ�it"�~����Ư��q�����OO	��1�H��֦�^A����e�B�aH����#T�k�]M���C�7��ƚ�G��.[WF�yzŪ=�ݳ{�_�(Z��Z�V��Y�_���'Q�VJ�D��Z����3�0��t�6v�����"����)ﯕ֜��ٕ�n�9n����X�g�W�ۡ�s�.w+�:Q�M��s���e��+\���-S�n�qy!x��@� R=�n��j/SL)#1#�Aa�2RS�g��L4[;���抔3���L�\@<�6����h��q2���zR�b���M�j�7����Gd���{�CZe�EٚK6.b�֘�(2sF��BW[ߍ�
2�L�T��y���!����sF+tqt�.��y��@/�Z��wz�Q<�]O���zM����Y@���U6��d�{�Q�p��l�x3 s:o�!o����{�Z��li��~�4M`2�k��b�dbO�JV1�'�ͧ�l�*���*cؑ�v9EWEi���O���Q5�e��`|@�����ݯ�*�D7��X�vO��,cF�f�z=Ł�ߏܻ/w.�^�z:]�L}w6c���{p��yO{����0s��e������ `�(~���ެ�it CB�s�(�|]./~��<x����0��ݽ�q�k7�M!��湨����z��u������X���æ�lv�&44���%��t�9��#��4<�ѿO�屛��L�������y�Խi �40��v��`$O(��K��;�m�%v��IM>��=3*(�9�++	�������ٟ{� �:Q�W�JU���QEէn	�������Z�
hJ�1-G\��oy�Ɗ��ZQ[C�L���PB.�zf��y����&X��V@����ē`i���PJ��eƝ�~���W��&�9�f�mk�p�)*�zlN{t	MҪ7��w�Ev������aHٌoej���v;�a�r�l:�P�6��&���N;H���A@*;�i�@��'s�tq	=��.�8����Ji�n��a3�'7�ӣo�`$�\9��#���l���#2�kH�+���p�ѝ��Þ+��I�^���}�Wd��[=���m���b��n����N>��B�x��-��V/n�����G�9m���\�\zAl�
jd����å�>i�H�!��G��,����U~�������H�)Rqs�~�	�ŏk�EG�f��;@��kDJ��C��Ɣ����2퐦�T&�r���i�������S�����7���M�M}�w����s�(>����������K*�	Q����˧���9���e�ՕP��=r`�ʔ,TBCAZ�^�Yվ S?�W�����z�h-�R�ԳC
O���Gچ�\�]�F�����Ⱦ �(�a��B��@�)���j���[�	9�0Q�!gܚv��.pQ�8�=&-��9!��vJ�>'�Z��ۃ��d�ѣ��MW�z���am�{# *r�P�̌&�|D�'���l��{��	g���A����V.�Z��ǓU�i��3�
�Q���a���	mO(��e^���b��dnD*NMq���'2���t+cAc=�t1��}3|��^�E���t�Ve�*���E�x��;��}^wJ}F��NH��9���=\��&{b��кN�y<�i�`KM`�ВВ��!*�߃�'!w��g0JbdΞN�ϚR�y�<��7d��(�ի����U�&��[����Nڣ?�Ag uY0��=?SA��K��郡l*[�N�
�� M7��6�<��#�,H�L�`ڡ���&�,�V�'IR�tEj{��p<][$*O�i�z��CS,�tid�r;��?�z�9���"M�������[Ov�)�S�Z��E�v��6y�.��3aҸX#�}��+Fl_�}��
'���#�����-��:X��D�+�?��2A��\,���`���:�>ޖk��G����S�7�o��C�3�0n������^~��9ܯi��+𣤺K������|�%՞�@nM{ۅ􇗺����V����V�@�W��X���K��m����xo9a��Dmآ�E���ƿ�W;���	9��5�o]�@2#%�BJ�����[�`���T�����3i�e������%v(v%SvO P����=����U��>%�BA���H�_o�̬Tv�DBDJ�oӴS����'䴳��4�ݑ[���Z��¢�V�dJzJl=����`�k(�C��&�s<����&03��Ќ�)�J.���-|�Kh�Q���D6��� �	�+�d��'2�'�����б�������Ƴ�j����ѾǤ;����/xލa߽)����?�+T��n#]6�\lP���*H:���(B"�5���R&P�x�M�4�����m*����S�˧�r@&'�V��o&���5ZU��`���Ƭ AM�A�H9�%e&eb]�E[�*M�*n����������N|�����M�D���'�UIDIUHd�Jċܴ��}��.��0�X�R�)_�̱��� ��?y;��3)Ӕ��_@�p�X�()�	cވ�Z_����dެx�@�!���RaKM�}��M$��IU��u5�!d�(�5�;F��(���F��7������7�S'=`�=#��h��SA�%���r�;�:��ns�3���j�������\��|Ͽ�����?1�2: ����_�ٟ��˸������{�=��$���酪���k��+���q�����f�KI���ja\/"���zC8b�=4z��r{@������G����xiKtE'�zPTm85A�#�d�c����>)I�"��gMH�(^�iyfFJJ9`��\pk���t�|�|@!k� '$0)Zv�>�����������S#JU�-��DG"����> ½�t���!�'�{<pՓ�^K[qF������
9��*�*�T�lҞiwU���v��}-�:�'ngpR�Xt�@p�GiIN��2��e�t\x8N[D��v�D�����E#B*��pk���-­���.����yL��X r��k�ivD�2���MWA���vf����^�E���Y�U@�!��. d*����
��Ҿ��4%�\4��!�"������3v���O@�L��K��'�O�佧��̤��&�ĩ1s#BUEm�.�<SJs���r:��� >NJ�>щ���隠G �rﵓ��"h'-j�,`���W��(���p��C�])�n�����>�|	�U=�&��-mr)��փjۋ�I[+R[��L��$���"�T��HZPX�XG�\���).��)��@�KL��Φ�ժh�J��Ac�>TB����H��nl,��&P����=� �
�V�Aɮ��;�ױH����}���I5��u�g���)#�؝��*S�g���X�H��{��}�E)�K��7��v~��,�Q���w�9���G?���
~���=�f��˷ԁ ������+��q���_hy����m���<1��k�/Q�"%ki�&Hb�0i�N�:���*&X�ܛ��x=��hxI8������V7�U�C&`l �U`Q�PSA&��V�'�W ~�0)R�P�ȔL�L2�0�f1QA��r��i�;�ܙ�`���<!���VA[`�ښ��Y����T���<�Ӄ������5f�� }�2^d�<����h͉+���ݾ*s��n���ҔX.�����2��r��Sʍ�y.Rk���&�eB]
8=U�߯����wcW���������T�E�ITx�j���P�'n)�4/x���Ǚ�JΦ���	9eH3)K&����S�>+n���pkG�mFW"D���+����}��6̨��m�.o�J]ꛣ�^�lm�Ex���~��Z�.���. �Z�����	uf�(�H�V��݄S�q:	��)���gԚ���%��ٕJ�n/|�����S��#_3�Cb<,�����_�į xE��,*ߨN/��[.��[ޕ�)7�,�rc��D¹4"m��kd�e�&Mx7)�De�k�,�jEz�Qr��m�@��r}dL�y*iJ�K�Xu�mn	@Zj˵�,�%�9Km���V淋���R���|�H}mym~B��Vkˡ-ׅuIB�mAʌ�����q��i�����B�N��]ɸ�`\��КE2
d)�vB����hb:]��HPP]Еۈ H��u�Ż+]�����dE�"����Q�;��'�#u�BDS�;oM�{爌Z�q&�a>�@0{�>���>xe�R�#O{�2]q�-�������������R�9�-x�v���Ox���_�{��Oѯ�ҿ���A^�E�� -&�)&<Cb櫶il��R����D��dZ��\���lz�{��f����!���&N��@2AQA3�넂v���z�����+de
��M�1MH�=�N9{�3�JW�c���].pw�w����z*C9!��Ҥ�,Dt��&ί���Μ��S�\N�O	��*��9O'N��ʇ%]ޞ?�3?]�|��r��R3���֟Ih�J���n(������-���Vlr�js�L��'���������9\\�5��Y�q}��YQ�KD�[k���i>��c��[A*Y/��P8=��J��e��yλ]�23@���5��ä�ĉh_wD�/3������?����²]KοNە�9���D�`P���F�1Е�[�pV(�GE�B��:V��� �MՆt:i�_B�	����Δ���K�Zv;�ۇ��R�I��x�s�j��P%���y��SO�r��xI�o�i�Uʻ_W�/���
PK�%���VJie�qj<q�����7e��[,�"��y+��v��	�fc�T2���tЗ#�X��'kgj3P��5�S�L�z���Pv�L��Ί4�EZ�5H���P����"�a������u��Xj�3Z�2�_��m^^���h�۲�g��nk�����T��z(:CeA[ԥ�-���e9��#)���.�*{Bk��:5��m� ���־�D6��SS��' $Ӽ��l�J�#��vng�k)��0A��}��1 h����n<EYi7587"<%��Z,�;��R��xJ;K#��W����^*��J���.>��[�����-w��K���>���4�˸n����?$*���/u~{�si���fH�!��0���n۵b-�=�
�<�����L7��^ �ʱb���߱�l	�W�pya��������+�
����`E6jU��.�֐S�R2�2!sƄl����1+ Ta�
�|�C����%����gO�6����v�2	8w�_Ki����/�gSΟL)����IR�s޵��V=<�T��'>����z[3CiBK�' �g�y�o�z��W�
 �ZѤbYf���=�����^�ƽ|��5?|�Wi̜H[�Z+��L�-;�tGTo�����E�u߄wJ�������rI�3Cs��I�LXTY]S��'��Ki��T�%����z,,`�jR�["�*-��GA��L{�`�-�z/�C�T�R��fPv�RR�uG�}k=�ѓ�Px�&�U�[U�U����Y��ki���R[b�K[�R�)�:/u��~��ݾ�P3�ք_���|Yr������?�z�g����4?q[�p!�ť�|K ��}�SH�ۨ8y����l5����5���?���x~���  �IK���eF���!��m/����y��Nz���г�������;�����<�xWP��@��Y󤏧X�+d�RL�XeW��Rk*��tD=^��%��i����������R���f7�Y�t���A�0N��st���6C��P<r�3�X�\� `��X���/�6ʀ���ƞ���P&Fd��N6��],���H��i�������N����������Oķ� ���G��w��~	iaҧ����.˿�d����&�TZ;B<N*�y7��f�M���G�X��+?Yŧƞ]�.�^A�!�⣴�͏Tتe��ײ�ի������z}�Wu����
h"̲`>��Dؗɫ��r�dNإ	S*&/��g�j�(�w8L�qQ.q�p�������S�Ň��ʴ�r�ʧ	��=�_�����WN��i*{-��|���~���r�0��	���	w��^�w�RI8=8�x\p}\���}������Z�ڽ{�ݿ�w�S��,���=,�	��D��,hMH�uB�ɋM�D�o\1e��.�rb�2A�k�+Q����c�i��~�wW�ֻ���-�N��d�x޷$i�95��Ě�sK��wAV��&a�=0�o�{�M�7\!�*)TD�6�(�q�nr�n�r�ׯ<���8����^�_k�
�gk��.tw�6P��2��O��/t~�{��S�[O���3�[���ew@��HE��}�F��7z������~�+XN�X���f`>bz�I��5˼�\�$e��I�i�z�b�E}7P���4�ҔT�����j|k�C�j}�&�,G���ꅔq<U\_/&*����4pݴ��6�c�F}*�����T� �#&��Z�u��Zunqs[|C
ٍK�Q�H�����5�m��
ǽ��vS!T�^�m�ZJ�۾�T.>���.��?�����C�,���#o�R�'�[�@���/�P2�_��SU����j�ai�;[��&kaZ���R����pk5�9Ϗ�$x.�+m?��O���#޾����6�ի�{�+|���k�W���Ҁ�r�um�>�S�������*6PD�]���p�i��~qUP+ �q��;�{�$��}Wn_�zpk��������y7}\���~��_�}��اtwH�����l��t���^���Ջ#ꬸ���)�N`͠�P�x��5�EЈQ�RFk%��u�_b�9����6L��z���X��^~���p��C���ⷿ�{s�U��g>j��`��p�O?�=}j��km~?D_$�}����\?�;�F�|��x�,f8���"g�����Ԅ�i�i^��+�
���r��;>&�%&y\=�]�pm{��u-�+�P�yʜ���M�Ȥ/{�ڏ�o�~��P8%3+��J�B����bG)#s��8�\v���)���xˋ|���?5���Η>�1(	��5�O?��?�aY�����I����iE�I[��XߢV�0�}h�o�ӽ���X#U" �/���i�-��ke�"�
WU������#��W��'�bC)���QR���(�$L����!>�b`�&ȑӄ[��ؕ���jŔn#c�D	�/���~�ٯ=y��������n�����ҧ_���$4��sϾѷ4��B?�a���{
����an3Z[px�����{���%Ǉ/��J��K��Z�k���bAkC&��^�M	�
�B8͋�N'@��i3/W�Zsx�����F%\�I���+���'�9#%B���d����)���pLލB��Z�l#Y}��	 2��4ٰ�4������k9��J�WA����>���8��-��7�������@�/|�ؽ�i\��h�G�y�����^�N��wf�ߩ�h�����Ui{�Z �Td��^��G��7mܫ��#��f���a�
}������J׆������,*�#� jC|��I��WhRQ�u�K���%d6�f���i���U����\���w��;O�}�c��̻>��/}�ݓ�s����p���7�6A ��_�E �VA�3�y��镯���t�.>Ȍ�6ײ���{ҖI*�r�2� ���s�>m�P���ٔ7��@��xS����]�>�
U�b5�UKIu�����e�i�GǞ�2��qA�x��y+RE`���{ΩW��(/�r?O��r��/Q��H��r��;���/E����=�;��O���`y������SO�vz[m�gAx*ߣ��Է�ջ"� �C2IUXUX��h��d5�㒮��R���Ůq4%+a����{�}�EM`B\���� �����MLPb7MP.>�E-4�4�\�����������������O��,������e���[Z��?��O �^�����>�j~��[o� <xG=]�u��
�>��{���і;m^��T8^�Z5u����54��mmV5�&�'o
�v�k�z#�����3!�U���(q#2��ܵ!o(��p�˔�g��I�.�,̩��2_'N��k����?���?���^�� ��}��F���t~��[��?�ҳ��P��׸x�S}����[h�Ro�N"����P}Z���[*8a�������խ����c_q��
���7�.?IB�,�m��*����>�0��וf�����m���5-˂��Jɨb�1S.Z�W%O��������px�s���/�{�ٷ�-�<�����o�� �g�ԧ���x�|��� rxn�,�����6�<S8�J�U��o"z��o�N�Ts���(��yO
�jz6O���"������
�6C����ܭ-nk�$))aۤ>�i�2"��2%%NB����J�f%>�
����K�ӗ�����qY꧙���F�^|I_��R�L�Uo{���ѷﷄfw�/|�v�j5��@� /����#K]�&�h�Y[M�IRQ6�g"�邈n�-�iOL;UL
ͤH`Ndc���X��J�d�G�*T�`�FB��5���B}�+��De�8-3��#�*�2�~�'�V�J�����<����������O������/�u�4��|��ѷ"�JT�}�8�M����p��~�N��p:ͻZka���:�D�ۙ���������nI�Q�h�k�y^��T91133)"�b��f��@�Y�Z�\r΀���W��X))1	@ں�-�1QQc�
�
�3���9�gN���U��N���,���>+���S�S^��N������¯��'�
�����w?�Y�؏��}�� � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ��1�Ӓ������   %tEXtdate:create 2019-08-11T01:25:28+00:00�d�B   %tEXtdate:modify 2019-07-26T05:04:57+00:00�_�X    IEND�B`�PK
     ^�[d��   �   /   images/a262aa33-74c4-460b-b0ad-c746896f6744.png�PNG

   IHDR   d   d   p�T   gAMA  ���a   	pHYs     ��   %tEXtdate:create 2019-08-11T01:25:28+00:00�d�B   %tEXtdate:modify 2019-07-26T05:04:57+00:00�_�X  �IDATx��{y���u׹���Z�j��ez�����L�b'������2�eH$BaJ�@�dC��`�@��![G6NlϒqO{2��=��RU]{��ۿ�����1�'��n�u�{�[�=�s~�w��ʥ��1d���1@�lL �1d���1@�lL �1d���1@�lL �1d���1@�lL �1d���1@�lL �1d���1@�lL �1d���1@�lL �1d���1@�l�c@�a�z��Ti�R��)�|�H)����]ǧ0�Vg�¸K�F�Z���=:0��y��8L^a�&����4�"ϨH32ʐv4������>Y��6����=�n� ��w�H��)�~�����t�g��!�<T~V�Yz`�����j����ר�����Z�:@N�NF�ޢ���,S�ޠ��NY<�Zk��J��� m
& ̡T�nW���]����{}*f��>s���m�ݽ㯐[����u��)h~�����>�����R����h_�М�NݴC͠���ޘ�g>�?���g�~��P�R8葉ڤ+�T�O�8�,�`�UZ�	!�n�6�a���y6O"ǭVk��D o�D9~G��[�m���^�u�'^"�[^���O�N����+ DF�u
��v�����/M2�P���&���8\��
\��w�z��V�K3�K3���h㇟|������~ݟ����W���f�ȉCD�M"�!Y֕�.���n�Sf�	ch��G�&�q�H5���*o/��%�ݼIj��KI�Z����.J[�(�\ׇGk2�j�4���X:
A�tԿ�M?�Yg����K_����pkC通K�23�*0o�g3�$����0�v�g~�/+�W7��|��ּ�,un_����� I;���\��u��_},�~�n@"��-ob+b�v��X�I��f�L]�Һ^��U�8�E'?vV�x�C�k�;���M�}$�DLi�S����mQ�Ņ�:��(_Ug�����F�����	��ġ`VcrDqf*��q
4SU�NLm&U^�������G��i�8�3�.�۩.tؙ9|fp�[�D����W)�lSg}�����ѡ��0���%�]���pa�[���>PD���~󧢵�� �v���ԡ�����?�j�UZ��ε��@��_
��e���,�=McB�'�pt�&���.���
{^�K�zst���t��I��#���\N������r���4a�8&:��i�M����fS޻�0�*N�� ��%
V^��'B�%���w�1�@��Yuh$L�wQ&�0�3��	B8f��e�wA���Hi��%�?�p-,$|M^�0$ln���ÃN��'���S���;u���}���~g�| ��eP�>Gӧ>�����)3���I�+Q$d���򼴍�*ձ�aѣ�x�M�"D�ܤ,=E��Cdẝ��HKb�=~���kur��0!�-�)���!��D��)�px0D!�`����!��YҞ+sU9��x�T�J�,�OR@do6v�"�J��:������gB�K���E�����Ԡ?±��� ����s�Kh���+��7^mn����&]
wV�:{���i��u�Z�|�I��'��&��=�{��֠}m�r�<�r � ��c%ED��*�	���8k�0�Z��5�׃S�w����i@�g�ׅ�âz��w[�D'��I�Ar<��a�L*�އ\M����G�+�+��߰s[�����
��T�l1�z��=��.� �v+r�v��[�D�KO��c�	�K�N����[_|���S\�m#$ł��y��s��~)�oR�"�qm�ߵU�/�ԃpw��
"��U��2��Nڦ�<���w]B�^�X�U�F�ozZ�3d��(w�m����&�ҳɂ�d^J��)$��D� ]��X0�*\KIy,`Z�S�oا\G�څ��k�ԫ����G(4ED�+�i8���\r;Y_�Fa�bn���V�`���܉'�n��z �}G����#7��{�B���/ga�`:��v!{�%Z�A�q�P�w���~CYT�UM@u�C�D&�����m�O���KY`��Cs5�e@Q�f�\Z�m��-�%*$4�H`ٟ�i2WD�L]VCq�)�~�dQE�:�)IX˵喝
��O=E>U�)��:[[��Bβ�saȜF3�`H)E1��>>CN�?оs������=��;k�.�$�ҩ��x�~���p��_Α7�p�&q�@NTNu����	yф���ά�K���	]�WQ�6���p^S7����N�z��7e�WY��G�95�F��+�ÁBሚ�t�D�,UX�/��p $o�T(M{5�ր�2�gBrNa��r����
�7_׃s̟z���S��\!3X#߳�7��0��p�3��<��D4��Y���b4~�:��˝�7^�H,P��J�ܰ�K핛tv�y��'�w���y�����a2UNQ��8���/#z��!X�4Ee�w�.���9��� �ޙш���.U�5rI?��H�>��!���~�
S%6Y!
F��[ͪJ�亢�"PNтĚ�Ҿ��\�*Ȫ"�윬c�*#��%j��}���y�����﵌r+���Q����5��#w�<� o`Nٰ]M�꿞=��3������i#$�z,�Sm��}ݕ��}�{���ޑ(P���̄ZP^U<P��7�E�)s��p� �Jg�"L��s���8=�8�&Q&	�A@����d��U��Z%p@ e�w�C�� jT���xbn�[惟^��.�ӶxmhI�R�8��X[;��Dn�E~�^��WR# j.�5�RX�_�r�+��]�ʜ-��"���^�t늬դ^��G� x�s�⿸���ԉ?��Q���:�o��� j���g㝫���8��/�(���E�a���r��j�Tܻa/k8S�PY$����I:9s��;��1�M��0RE��<�Rھ��DR�y�2���D�*��$�ETdF�(�8*4�uD)1{6G�����@]-��=F���r��q����0��؜(y�s����@onm/;1�y�&�'����YH��.�KT]xP���SY2�A9qE���	r��������������έ����{>�����@S��/�c��eu��ʘ���	9%�Qڪ��x�"�4a�$ۡN�o��t���"��Z�m�O�ȉ�/SmΞ���%���b[�Ap�����29?gi�IH+�� p"��� xH_�\U�#�8 �=���� �Ʈ��Π�P|9�G�ex����)ݥT�$��5����)L��H��=�c-9Q��3�C���"��BS��4�=w9Z~j;�~����i�ě�}Ű"a��$�ڝ{<��X�1x;"g U.�*Y-���$�0��=��FG*��wi�f���zK�l^���~M��!t`����E�ޗ��5@���R�3�7(T�rl��<��T��;D5�PD��ѹ���d����\�p�!ё�I�#&��Hn=�Afa������[�M�����ox(�}��jߑ5*8�ҷ��D]�kduƵX���E��e��g���s5��w: +�KaS��q��0Y*rc�dZR��+J�*�G�Zc���"4A30��7���ޯ�Q�/�޸D���xs��D�p���.a����6�9%�3ա��XYn�"L[�˭"� �� 1��MR��(a�F��Pcs�6���w�UD#�ƴ�k�:&g�ɻ��P����]^[U��գ�W�s�%���@X���f�S�?��:	���.�B�r8�魐��57�ڛ'�G�͢�k�$�\.�Ӳ3�������|�R�|�|�܁�ڴ���P-���ץ�+Qhlo�)�^��˹!;�S��1C'�aT����Uz+�t�$½�;j�9�d(t��x����m�0H�Հ�"�Yi��BT������5���8R��/6�̽L�FKn�M_r;4��<�\�؊K�E~�%ut���ص;�2��e�@4�����*kY4S���X/���9������
�Y
p=���8�8,Xp��ͽʶ,�{F�>Q�H�Q�Ĩ�SCsnF���g���T���胁őX���}d�$PJR�_Ξ)�
���֠�hGh[���j����'M1��'�>�Hd�D5��8R��,
k"�Y!���C��\Ŕ�AqY�(7��=�b�H�Kr6���e�Nو+_2Kc�����]9ڪ�£���a�Y)@+[3N���?�u@Y�I��2�a^I
��a�|&R��e/Ki�Y����������<}8���$i��{{*2m��"��ZjF�R9\ c�YZ���V�#�j)y�*j�Pj�T))6�����Q�Ƥq��(؟���Z�K�כ�ό��bЃ�l%"w6�s9j�k^\	�m��J� ą�|�(�MҜ[_$9��.e�h5e��ؾ�eJ�F�M0>ߵ�����C���W��4n�&8A�{�^�U,|^x[]��~{�/ۓ��S���r�*��VM:�Ibh*,J2�{`PY��-s�&BU�S��!b%f6zx�"(���u��_NM��ϯ�]	p���[ِ�������C(A��ʚ�&V�%n��Ҳ��m��XZ)�77�lH>�~X���w>�ⴇ�P8Y��e�z��>�!,�S�}%�[��˕�P$+!g�0��Qd�F��-¬��X5�@�iPE�vٟa�T�r7����hޅme���-�a�����Ɣ��;GМ��`��?��{��~�ɿ��'�������C�r.r��Hf@�޾�ѹ���J�ƲЛ�J8����1��� B.N0���=6ۈ3ei��0����E+<÷�V�sI���ϋ{=)�[Q�����#�Ap$�r��q�a(�`�FQО�Y��jî1��X�~�ʍ����C��V!��e���z�3�r�[)W�`�'��?�%��_x���gg�~�Gk�7l>�UH��E�ǡ.J!�dv��:�Ք&�6N���&�1�Ri3צ��=#*�!>�
�mI��P�{�0$j����쵲�ABf�Y֒#����j�����K+GDA�iy_dv�Q��M��T�b���xm.��P�vű|����g�e�X:�JP�W�})B����qQ���H��=���t{��?;�U2�1�	���`���'�~?l.���!Q�w+gD��w��<F��8� ��#$�I�G^�Aa)�un��-O!
c�	����ԋ
�	i(6;��R��	�����|#M�RJd�sRa��
VO^'ANL��Y�k���PY��6��Z��<mMf7�4�t&{,E)�*v�t$F[��1!,�Y�y�s������}2;7YW�����c�q�u�x��T_,.y�}?}�y��,�Ӱc���Z��团�`����)&��|,Q�%�3�Z�T���OD�R����M�όy����|DJ�s�<���O(]��Yx�L�|��X�ǀ�ANY�ؘ 2��H0/n]��z�̍�s�B$+D���"Ys3�T�
Z9?�`NY�h$�(ͲQj�cIQe�_�)��T�~.�t�̳�z�U:�����!�����(��+/�����_s���n�E}��P�{o�����\P���r���J*@S)GG����Ae!ȋ�G\^���P4l�ݞO��+�;�,�}!<��F�R�L���=T`��v������[C�����8/QV�I��@�[�%���-s"� d����uH2��<�P1��:h��gI>�b��I�ѯ�Ch5�������7���st�]��\�v�~7-_x�K��c����YtH��O�-��:�F�"iK�\Ŀ�׏���4�ϐ�x��
�d���Y���Oi+���V���!���h�w�e
 Ң)�;�YِR;@nom��@O���#&���V��UBq���ͯE�.E��4�΂+�5YO�{�F��`d�mp_>��A�Q/���t���h�(��;�_�Ï�|���|����k����W�n�u�1��H꿡������H1��;�^�[��dQ!G��Ȇ2�@qN��A!)�k�ҶVE�V��u2��f�u�k$xn��(0p��]6�F�DSFF!^���+
��l��?W�yn��\Ԡ)v(�6�r�u$��k�
PEO!���$c��'�,]
�Q=�st�t�\���ׇ^�������yo����G����!�v@fg��k/����?���������S�ҡbЅ��e�~i+e%BVG��b�f�n��Cb,�N�w���Ƚ �T�k\�K��'���V��h���]�B�� ^�>]�����lM+�wJ�2u������5)Ly�2�MR�UI5�}��L��k1����k�	oN9Vy�߇�#Y1a;T�&�.����í�~��c������c��i���?0��e|�)�u�T���[itď��FC��'�Oūx��i�\�s����3Μ�-���'���*��jו�6$���-��4��"k����z��J�Z��sը�Pvo]B5��\Q�{߳5�[%g��ٽ)8�eC��0�,~F�_�J��@t�4U�*(�R��#��>�M-�hQ�3�܀�t�m�e�l�a=^s��������~�wx�̇�w�������K��|�vV.��}�?���?b��;����"�e��=�f/.��kT_���En��u:��!j֏H����V��|W;^�K���MD���*��4���AUy���Ss)�f������|��#;���.�u ɎHw���.!��#К��BZG�����8�%��N5O�zGSY�u'�}����O\B� ��Ȯ�H�N���a�'.j�.Ҝ�g)�#p+Ti-Qe��E����a{c��n.�������ճF��w6�S'�������:���H�}R�sn)���>���z�&�3�Uϣ�?M3�����Go�V�3����W_s+��&��N/�G�+���Q���Yz���k۝f�f�����@{��㙄�"����Ju��9�r�i�v������������X��� �:��LT��N{�/)<L����l߭;�f�y�5����ߗ{�<r����.��y/��^"�@�ZI=�F?s �<8^0��U�s���t�s;���H�}oJ��y�V_y�q�����d�����~�v>��n�%G GS+]A1��4��x*�������D�ۊW�=W��k�>��/]�򯷛G���	��P�_'�*�.kqgv{��RoQ7�d�*qR
}EQ��0�і���|�>9Bൕ�e2�-�i��,�bؕ=>'K�w6h8�KG��� `<PRvP<�)���y���?�ɠw��G%�:��=SSt�0Eu�婙�H�Z��S�z��M�yם��?[�N����s�<E5�X�����w3���}ȁG�CwΝ�J����is��*4������V��6}���ȼ���T+�����ڌ)	w�9�_����W~��W.�C��%ZlP-h������}/^�L?N/|�b`|P��֚l�nܜ��U�y�ؗ��ڇ2�[��}�[����<t9`@K���w:�W_���BՇ�{典H�o�4�f��2-��_���[�p�C��
��9.'u!\1���tz�5|�|��>t���W�9��D<����Auߙ'�~�s�"�?�7i��D�����G~��_{)�]D�D��.
ɵΦ��j[Mz��ץg�͆t����q����r�N<�m�W.~���CTi�݋�%�W�ƉluKu�P����FS��5����� ~i�~��wt�?�}�w�����O��O���wf��c�W�c6&��٘ 2fcȘ�	 c6&��٘ 2fcȘ�	 c6&��٘ 2fcȘ�	 c6&��٘ 2fcȘ�	 c6&��٘ 2fcȘ�	 c6&��٘ 2fcȘ�	 c6&��٘ 2fcȘ�	 c6&��٘ 2f�D�{��w��    IEND�B`�PK
     ^�[�c��f  �f  /   images/c88b2895-5e8b-4a57-9f9a-b80dd50058b1.png�PNG

   IHDR  �  �   ��ߊ  TiCCPICC Profile  x�c``RI,(�aa``��+)
rwR���R`����b
����>@%0|����/��:%5�I�^��b��Ջ�D������d ��S��JS�l����):
Ȟb�C�@�$�XMH�3�}�VH�H�����IBOGbC�n��ₜ�J� c���Ԋ�_PY���Q���Tϼd=#CsP�CT�%���X�}�����ߍ�������k'BLÂ�A�����΂ĢD�33��10|Z����� |�'�8��,������z����j��N��������.j���p  !e�2���   	pHYs  %  %IR$�   xeXIfII*            (           J       R   i�    Z       %     %      �    o  �           a���  �zTXtRaw profile type icc  x��S[n�0��)z^�8~$R��b;^eW�J�ё"�@`H�n-|DI�D��@ȴ�v=L�"�	�s,`�ۮ��z����"H����pz����3�ͬ,9&�h'�tN9#���(���d>CQ�h�|q�k��R�R����mOi�q�6�Z�ܶ=���C�>hrK$>���U`�͚t3�s;����%�S�T�c��\���~�y§b�_"%�G"a=}J�H����|)�Ni����2��yl�c���r�E��|�7$��8��s���.PJ����
��wq�8��P'��j����[ܞ�c2����g�+��|����RM�=�c2gҥl��ϞauTh���҈�\�z���줡㜥   %tEXtdate:create 2020-01-31T21:31:09+00:00��y{   %tEXtdate:modify 2020-01-31T21:31:00+00:00	�   tEXtexif:ExifOffset 90Y�ޛ   tEXtexif:PixelXDimension 1391c�   tEXtexif:PixelYDimension 800�요   (tEXticc:copyright Copyright Apple Inc., 2017���   tEXticc:description Display P3�y��  a�IDATx���|SU���M�M��ޣ {��Dq�����~�V*�~���(���(�"{�Q6-�-�M�{�'I�M������K��{onn���cU{�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!@��-[a츱�aC�5?�q8�^ݺ"���0�
�"���l�a���>C��p���Oo��vn����"��mE�9F�1\���?ۛ�����(:���c�X���_wlP(�ʔ{���=��|+��#}�Y��mo�w��k��]�o�������?�O�0�?���'�Q���W?s��3��"Sڶo�dՊ�}�I���i�f����gf^�t8Z������^d�g`���>�n�q�0K���k|=Ϗ���5�1��}���I0�p]�y��U��'3r��~'_{���G���ߢ��h������1o��v�#�����޵{�I��z�}Պ�ged��x0'""��!;;�߁�������t8�ADDDՎ��4���N����E�l4"""��L�����QQ���ԿTP�UK���	���sn������BDDDՓ}����{�������H/�=��|!'""�c�4a��sh׮ݔ�#F���u�}�?_+.q��p8PPP��o�O���m+�p���DDDG�}ǎ툯0;+k����C���PA܉��\��+z��I#<r䑓�\y���O5�Q�?�^D��R]�]R<�5k����q֦=11Q�s�*Yǖ�Ull,���0�C�Y6'"�`V|֠g�HKKS�o����T���Ύr���������GXd$���(T�:����=3+Y*��D�~2+3K��H�h#"���sx���_����`:͈�����O��;r��"""
f����6.��p�)�ggg��oDDD�����R�7Mgx�'�����"""
n�Cii����p:M{�'��]��QP3��SSѼE�8���,�3�:gOݟ�F��:�������y�
�DDD���";+;ơzI2�kff&���(��j����H�4�L��at""�`&��:���K@/3�^�a�Љ����nC����E��J膻��0���(���*w�^���(@VV���(���*����:��D^^>���(����p�Yo`� ��;w@/;�����FDDD�Mr�0��mPP�ϵЉ����iB��'ԭiՆ.������Q�V�%""�Qt/w���^J�&�΀NDD����m6È𶁴�{+�Qp�/^�T���t""��g߾m�*���6�Q𲧤�H������]��1�'���i��*w""��g����m*`��r���/��Ä�m�����NDD���3��G@g�;Q�S%�Æ����˝��(��3�����G����ΐNDD�Lس23��i�I��S��)U�ge���'{�3{NN�
����%�;Ճ������zdDD�i��K�DDDA�T=&&Ff��Н*�;Y�NDD�L{xD�t�S�:M�~Q��l6;|T�;�&L�Љ����=L��*w�Su"""
^v�a�ax�&�܉�����0�QN	�U�DDDA�T�\J�׉e���U�DDD��.K�|tV�3�|�i�̽t�U�DDDA��%���F��8tV��rK��U�DDDǀ�����t�K���˝��(���K�z���X���(��E�{	��7���t�,��ʝ��(�ٝO	�:��:űʝ��(hI����4�r��YB'""
fv��a�iz	�n?7�)���(�ٝ�sm��NDD��r���SQ�n��^�n��GDD�쐕�L��T07Љ����)U�J8|�r�Nq�DDDA�n+/�K�g@����<����@=?""�F��0;�*��乸ҵ033ii��k�.$'�@jj*>�����9	�QQ��S�ѨQC4k��6���\���1%>�|��%rpq��+�*3��?V�Y�?���Eb��-طo/<���<W�C=��,|��\`�!6&u��C�V�ЫWO0 }��A�&�f�1�Qȑ��i[�I@���p�{�W�܌���X�z5���;�:��V�ޯJ��(��Q�w�{�>)ͧ�Ė���/s0i�$t8�#�=�\|���ܹ��v��D$<�����pU���Ʉi7`��r��s�C��\�U�^�x1�����n�n٬��E�ۆ�)����`�E���Oq��W���GR���yv"��\�g.~��w|��g���;п_?�i`7нN��¹�}�\�-[�b����Gcǎ�p�W�����=轢������i�O��P\p���������O���u����拓�'�S��o�T!����>���2>�͘����3������_��p���T�Y���tf������ذq#��nԉ�cP'��'������ix뭷�|�2]�Y�^�z���'��2���V�{!�Pz^�0���*RS�µ��Gݷg��g'a��Mw���������{���#R�۟���#G���x䑇Ѡ~}u"
Zy���7o&��f͚���8��yHo���;�1��&��ޔ�y~&M�\�f��`�
���hܸZ�h�:�E˖z8Z�*UGGG#7'�z8ۆ�n�:lݲU�TU�[�Z�QV�a����HOKǨQ#� 1�A������K�,��߁�����Qi�tn��lC�C�����g�><����!??�oF׵kԸ1����3���&M��v�ڈ�{o���b�ʕ�a�:�~�:w���Gf ?/~�$��'�@LT�:�Ca�^��,���eʐ�0���or�gf��_�G*��`���9Q'>�>n��V=��v�Z�ϖ�|/C:�5i�H?�~n��L�<S>�\��S�5��s���[h׮n��z�~Y�(�2+&K�"��n�f9U��W\�Á�U	x���s���Űa�p�9�v\-�_+Ƴ�L�׭Kg�;��|2��֮�ù�J������ѱc�ؿ?K�DD!Nt�s����!�{Μ_���~�2�M�!����#г[7�_+O���/�	u�b��aX�l)�36�6��ѥK�� "�P�c�i7���*w]-̀^�n�ꫯb�d�z��L����p�Wb���hռy�Kƞ��u�@����~�H޶�����{�	�_xK�DD!ɕ�۝�i���q����0��)���_Q����p�����FTI0/N�}�Yg�����ǟ@���(�/3p�@*�y�m�4` ��cP'"
9�����rg��#���,F�9Y�.;ѵ[�G�M�VG%p��,2����/�L񲕁?���?���%]""
I�L�곛�k�Ԛ]B����i_c�jo��L������ރ^=z�R�'�N݃~�os�o�X��3��0s�L�{�DFDT��y�"X�X���x�����X]��:Ne��.��� ״������͞�}���[8�2{�u@|�ٸ��K�ɲ'8�w�{���O��������m=�c���xbP�p�ٟrss�����f��u&"B=�ߞ��y�v����y���Cn^���OV}���a+���N�[�8r��!�1�(ǲ��V�Nq�|����EFxȹʵ)p�>[u�rm��ץ���u}]�����OC��:����9�?���"��\}��ˌ���^��Пc�{�hU��)}>޶�R�5RT�y�s�C~J�@~�V�,�[9C�����57"��_@��U�?ϙ��+V�ۭ%cͯ��zԍ�?�7�/&:�^v	�M��C�0���-lطo�-_���Y"v���X�vV�Y��6`��]f��S�P�,�B�Z�ШQ#�n��:u�q�uD�����JZF233��]ۺ		:�*�>��)�f���X�x֩��s�N�I�##"�{hѲ:v�^�{����k�}^ŏ�r�*,Z�k�5۵k���t@����36o��{�@��]о];Ԋ�����u�8��W�3K��t�	�H��r��!���Q�X������u���lչ5m��}ջW/���u�9��a��5X�p�>Ύ;�q$C�����M�4E��ѭ[7$%��k U��{2��3-=[�l�K!�9n۶�))�����C��(�OL�3A��E�ΝѦMk�V���~�:��.�����MIJ�)���+T���6mB�>y��zK�D��f͛��,�u���㐘X��ZT��gVvv���}<p����_�X�����)�T��21g�(��t���k�8t�(���S_om�&���O<�R�>}�]}�������֊����m����ޭ{w�P��螛�J|���f̘����[�nEzz�����u^��t ���x�s�98��S�P%���w���x���٧��U8r%���5l�/��2ڵiS���C�o������
+T�g��>އ�";4h����õ�^�A�����8;U��n�����/�l�2���w/�k����(u�p�)����N>�$�R�ؑ^�/���<iR��r]d��_��*Hz����ᇙ��/�x�b��>>_�͎z�����5�\�s�g[O��J��`��F�ܰdrd�$���q�#T�T�9���u�	�$xUU��\�M���5�'���X�d����Hp�uT�.�6P�]O�ё"��*�W6�{�U�~1#G�ҁ�0��j�L�#�<Rbd�<������ս>Uw�MNNF���zoR����Z�.�1�sp��#�}{���� ���'��o��H׌2*��ґ��,X6�����?��v��#����.�С�)��^��C�`�l�R������;�ޱ�A.ǭ���*�4h�=z�K1�tP���>��U�ɫ3U[����{����z�g����t��.��c�JXd:ܛo�Y�ʮ'� ��%�ϕ�X��$�9[�
y���N��r��z�8�ޭ2�|��~��^v)U�gR�ve�]�b���ٳ����:���q�*w{�6|���0�Ǚ�Zɇ�J�͎��T%���_��u���<�+�ȿ����_�sGvv�_�+�lʾ��5�����y��ǟxݺv-���I�����B��Z�'_�.w�ځi_}�9?��ŗ\��{I����'g�k�|���z9ϕ+W�i���-�����nՏg�T���p�������KGb�*����?�{���K���Uk���̾R�����'[[��>'�dIAa����G��o֙)��L��M�����Z[j�֬^�u��T&��ge�ԯ���(g�pKU0߽[� �=�%~�q�I�������5�گ�GZ����[=�m؀�^{��9N;{$�6%������/�E]�r�Z����5�m��֩��,ǘz� ^U��7����}(���\�;=���}lٲ�����]J������7'��^��=�ܯ��5sm�?5o���ά���:v���)푆V*4u��p����N����|���f�?c�u�!�_L�[�n����|��"�>� /���]ŏ��VJx�n�\��cǢo�^��r&�9�UeXe�sU�-//��<{s][ɠIFsŊ�駟�裏�_����2��-�S�-��⟩��]x��gT@��&��̊ٵ�̮Z��?���H,���>��I����6��x���r�#����D�Х�2���>���:wB��m�Ӗ���[*J>�9*Q{z���믿�^�)��2�J(2���ч�R�J�H<�!C�v'T�%���'�x����d�k����~����@?���B����3�{5j��4dee��2?E�q80��oUf-�Ox�<�$�*�9
o��ffT�|ſ���Gzo�3�up��8���J�/�_R���>������O���$}�+S%57�F���Ƕ-��f�x��r��0��iذ~=�}�\tᅺ�_�SXO���/�£�<Zl�)��m[6]��������۶n�NjA@�����:lM.��t�t�2[�зO�׉�:�\jf���C����໻����m���WJ�Y��d��bX�w��_�h!��^�����_���*ڋ�	Z�1�w����a�B^���t|߁�'U
�4q�Q��-,���1a�J�=U�9�����NJ��= �r]���1��W0��	�ζʼ�������yx�����K/�Nco��^;i(��?��@���u�ȑ#�h�#!����F����9�[f��zH��������|���ū��s��z�
���zg㪫�
�gYڌ�3K�b�c���+�������Ǚ?⥗�cܸ�������eR:����ǝ�Tk��g��Ѝ�bz͹xť��`Ϟ�^����B�.]t5o(]!OR4��Y:t6o� ��ê ^�~��8ӻw4k�u���UT�h��]z���˖��]	��=gö����Ï�k{�E��T�ק�~��%���#"Ѵi3�B]Su���7';�R��Ҕ�n���VS�JЎ||�ɧ8���|�
_/�]	hLl��h��m�"11QG����uo�;v�;�Yg|�T�H��E_�.�W����=u�4LU%9W{y���D�=M�4Vץ�>o�$��RSS�a�l޴I��[_W�2L�:_r�
��0�L0w]���u�4G����u��n2�Jz��]�V]�dx_�X����(��N8�_�������ȑ��v� ���N��B��I��K�.�3�����Qڵ7oެ۶�'|��C�.Fq6=���=�;�^�I�$��t�2L�<����\ރ|O۴i�{�K�HG�C��r�򹦧�y9w��LӁ��}s���c��A>�G���}��/��\=�7mܨ�[�d��%�ף�t�S�֭[6+��)s���2>�����ak2�H!�ک��H 5��_�|9�?5��`�Db���T%�W^y��#פtu���ԗW��M�:����k�Nx�;�oÓO<�F�h�8Ce�Ru tu�+
�R��ۯ/���J�v�ih�����̈;)q�P�9����oM�R�1�f�Ϟ{n֫���]7�
�u0��3p�:N�޽Ѥq#=��s9���6�k\�����}{���#Ìf��:��^��"�>R�s�v.
�a*A�ޣ7�P���[�j�;W���W�dΤcۤI�����e�	�34t�x̘�طgRS���v":�N9�\}�U�qӦMu	�s]dH�֭��ݷ�����W`���"C�O���}zW����3�ǘ����yp'��o�駝����,���!�1�S��߅�����Y�,2K�s�{]VN����y"����}��ΕΠի� g�u&.��b=�q�ƺ7���zA~>RTfm��%�����H�Qِ�o�}�]�pB=����m곸��{p�-7���]���;u������gj��Q#1��u?�Lɐİ��?��kf@�R�+���D6Х�P������*p_Ub'�|*~�a�q�@Ĩ���'9��x��W�������6g�l��X��mX�z%�W	�۪�Ѩa�J't�P�\��T%���;q뭷��JPQ�L�p))�҅<������>V��t�Q%�����[���x��Gq�E��P��8R"�ݳ�w�'��?��*SeyUR��N�m\�а�8T`�*�G��"�*�ȃ�Եi�Jp�+c�\��-[��u-q�
�R��
�e��B�u��l�kޢ�=4LW97�_��K�jת���ҹ���N�ñ��?��IUb���{�͚4���^֬߀ѣ�ww����'�n��s�mh�2c��:��&������Izʿ8�E/�(ٰr�r�S�O|�Mԫ�P�{]�냅�Q������O�Ї���멈s�m�y2��|�q��aʔ)5r�:�����$C�j�9��nE�Bf��Gq��Յ���2����4��>A�I	��zg�'�q��ϬH�Zž�b���u���1}��qc�}˻C<��&g<�[��c�=�i_M��8B�)�|�ɧx���T�V�6j�Q�G��7�Ꜽ���R%����믿�vxz���T��^��K�DwZ�VaoǑ`0d�`]���۱g�.��lܸIWG׫�$.֊�K|ݺ��8����I����[Ǥ$<���X�n}���H&�ƽ8�{��1ͅ-���?U�1c���nƖ�-�c`��d=#�t���a�ĉX��[�թJ��1b�H]����ɞ�V_]O�II��V�	V��3f`�*9ߦ2��Q��J��u�_��T�3�9?o��!�Ho��]Z��~oSKK��|��:��^��X锸��Zzj|j^�9bz.w��멚�)N:rI��+�['P2�HL%&�6�i�ܵ��.2K5�u7p� =L+�]�#z�����J��t5���H{�|�ǨK/��\gW{�C���]����ݯl'��I�ᤷ�*wk�.=��`^ѡ���:^t�:�D�g=6X�z�J�+��;�w�q��ů"ץW������1F�t}��H�[O<�.8�����{��N��T`�>��C�aݺu8EmW���]���-��V�e��O>����+0��g���L{����t�{�+6��hˬ��z(��g֥〥)�|��a�葅����h*�I��K/�K�,յVs�H��c��	�N���Ց]���g��m�vM_d�p/SfVWs~��ŋ�[0�j��숃���V�ǞxLw[�'�([)�l~��ttx�� u��8��tӍ�ڸ��A�L�������mE��ύ7݄s�����9IIpР���O�x���1t�=iK'��֝�RʖL�ۓ�Fj�>x���J\~�e>k,���*�O�4��C("7JG+����S�#S�Ju�Ν�U���|�M�A�n+̋�Ƌ/�Pw}a����$C}��1�����Nt�p�Zb���W^#�j�G�)S�m�U��y�f�?p $k,��Ͱ�۳�&��KG���l[�V��P�i)��~��7�Y��~i�'�T.��SN�|;�����}�}�a���k�������s7�p�n���qM=%�u�]W���:w�&M���`��G'Z�l��.��2:$�~b}��f���A]�&"#�����)�Oj�V�Z�:�y�xm�>C�u�Ǒ���w�5)P����蒤�NS�*	����2��:wŭ�ݪ�D��.���o���f��.�+K��e:��^�\���0��$��a�k׮���B�{��]��Cꚻ:�ѱbJ��M&a.GMkC�_:Qe����B�+�ۄ�y���$\q���L��OI�.��=��?�:�X�b��5hr�9�<����uĀJ�엨J;�u@_�u�SO;�U��� �p��z���L��U-��V�[a���+���ؼE/S|��s��ǣg��*�JB����m�uQ��^�s��Uj+�2�aa�ͼC��z\�ަuk�{޹z� ��ҿ�.�M���[�5h�Hw@�L�kO@�*yw��	�M�n����̬��б�>k��]/�jb�db��[J�6�`�=D���3�:�[�
h��Kz��w�y�c�UU����0�!�^}UB)=g+P"UF�a��^����r�#��.N����72C��- �>=z�@�J���u��$��ye�лO�J��/���KH��uY�C:�z��(���3o�<����^v��F���,u��x�	i�8p &�5�G��ۇ*�"�Kf�c����(�;YAN'���*s��"1tL�v���u9�����M�>f��ܵL�*�W�L�b���:2ɔ���B�F�4i}�7\�c,XY�K�}9���B:]�t��{��_�׶BSO��1 �Ԇ���qb�>/A+�g��IV�mV�5�ef�U������U+Cw2S׿V-�m��zQ_v�ك��Vx}�k�nh߾j�Hr7M<����J&ϑ9�s�n��^r�ש�������"B���VMcNgH��Ւ����yU��n��sTt�ϭ$G*������٧�`)Î��z�Y���j��ڷw���n٪�l.=����� �+KWT��{�ԓ�4k��e�����H:�1u"ݮ]�J��}]t3���A�?�l��%ǩlgTڶ�ː@���;�`0���I����K[7o�|�y�w53+���m�Fe
7O�d�$3lU�.�Ռot4�_˫r����$ш�Yb1��4W�Ȕ���ɬ�i�u}TsV��]R�����<�b�0��;v�eJ��(qq�t'�ʒ�k�')=���y?�u*�픡��&ޛD\%t9Ve�U��쨌M�7##����=\��[Uj�_��d`�e|v�ڭgᓀ~dLDFE�q��Nz%�*ڼ-��b��/�$t���g���3�I�!���*s�I[]%�Ƃ��͝��Y��4C��I�oU�	��!+�Ig$�6:�t����W+N=j��IЊ�=�Z��k\�V2TU-Zer�t��*S)&	�nݢ�}�H&j��=���_�HaS��L�*�Y��?x�S�W�8��A�@L:TD������YCg&~U���JJ2��M�����۷O�U�w��`���4�eɼ޲�CU/BӴi]��(�8��;��[��.�?G��X�(U:�N�H���Q��H�������܇�}޷G��YO�����Ǐ�믿T�o��ѽ��z�����d�1�F��(8I	�^4o�L��]KJ����MWz]=��i�suj);�7�����/�yJ�99e�2�:Oα2w�T�JG��&�;F5J�$�v42 R"=��M��R�&��x#�k2��q6e�&5��؏�d����j�k�#�\m�5�m�Q�ƈ�]���:�i{�w��`&��[�M�*>
U��1���Idsr+7,�nS�+�����]M��W���e<���X�����z�Uѩ��jH	���n����dLm�zu�o���.;�Ɂ������O���V��G��*@Ib���C���l5s��J.�J�*��<�f"W]HG���e��@u�*��d�;Y����r{��jh@o�X퓒�F�3^�kv$Y6P��7o�3e5o��u�`>?��>�P`��+\��U���Q�*��SNUC�1G9��qk%�Nӽ�0���pk���a��򎥚�gϞ�V�;���˗/׳N�`��ʒ�F^}�5|��7�бz��޽{��%�KOfo3_IU��`)�hf��0HR��g=9�!c��5>�'
��L���C�v�\�3G�f3u���@T1�Yn���5��^*�K`?�a=fu��eض-�:f��#%g�/%EO��c�6����l��ZĐ�3z��K/����)�N�p"	��(�H�`)�W5�s����OT͝Oǎs��
M�?��$&�?f��:U0��8ӟznC�u:N�n[`��(�mHNކ�9�]�]��7�B<�*=Ʒmݬ���ڷo�zi����A�p~PzȘ*�gdT}�_��Z+�و���Ы��`^+�{'O�0J�\h�8��TT�Mu�H�ʽRU}'�zY����?���_�e��]	؇���%����t򓕮�ԫ[O�Ѷ��(��Ν;u�۪v�59���v��1̍f63�٤������Y����mT�:1������]޵Ls������U���v���_�d�R8�rF[�nÌ߫�J�̭>RS�v*���� Q�������*K:ffe!.6�J����]�N�L*Svq9������m�2��Uږ����۷��~�]���R����ft���;�-^��k���Æ�;vbʔ/зO�c6C��gb����|�z���#q֠Az-i�O�^�zhּ6m�^�e�Mz�}\_s-������6��u2;�$x�����BNN�I�d�����K.�Z�%yd^�#��n�Ն^3'��%k�r�U)}���^��u��]vN9i�Q�b��yr2>��s���d6�����mZ���O�܇gq����1��_,�"��u�֣e��
[�n�ƍ��mXY�֭u��(ڨ�^�nv�*��|#d	S�z������H���.���R� 'AIa�������������t�m6\~�e��/�q�:��ٰ=y^z�%t萄���G�)�L@1y��X��?�7��s���0{;�������`�1�Х��Qe
N+LtE�i�쟱{��>���٫�^~��ߊ �y���T@�a񬁕+WaŊ�8픓z\��������s�~��*cQ6@�&MФqc�h���:�����N~3u�	[yU�5��]�}�Νqɥ�`��qz&'+�&M������ȣ�e�i�l���{((��L&�hּ��'A��9���[q۱}�f�*���]wމvm����ٻ3�NG>���ckšO�����}'R �=$�����s����>uON�2����.\�_���Ԕ�أ�d/:��]�>�p�'�se6s����巽BL��:/l�
�W]}��6�[��e����+HHH��s"�ë얔m�*�?�̳ػ�[�z"��.��{�*w�R��ۯ�;��f����0u�T64`S�����|K/���ŤI��úw>ё����3�w��S8�����^ݗ�^���k ��r�ÙY���U0���;��2�UI=�S]�h�����z�I�YN�l2����~�m�a�S��p���؟��}N_��o����W�|�^�/��,^���dNt��7�|�.e�:ݎ^��?�|UZ����&m�'N���N9�J�/9�e+V���^Cf�� ({+JO�s�=͛5�B
$��ڧo�4�GX�1�=9/�8mޜ����W|e�Q���o�nW;g�uV��i��ЭÏ4�y�d����Ə:sJ"\݀7� ��*O��+/��6]���O�^<p?ڵi��	D ����3Ĩ��x��`����E�.]�>�Yg���y�υU_��[6���c�L%rmZ�:���j߇^��*�[�V�hѪ.��|]�
���O��UW_�y��!+Ӻs܌�CR�x��'sd�Lxz��^�cǎՙ~o��N���5ADd�^��j1���<�Kܒ%�ωe@p�v�����ª���n�{�X6d��a�oa��ŸM��SZ������6�I]6mقw�yWW��L���NJ�W_}���
�۞eY
��oT���*�;�����J4�0t�0�ya:�kW�DN��c�.<��p|�ŗ��l�$,,�^{-�w��`NU��s��_���V�z~~�|��G������n|���ҫ�ɧ��?{�j�v��|��hP�~���ccbi�?��}���3rM����t�SB7ٖQ��XRU7��0l�CؽSz�Z}A}����O=���'�����y��'�u�V��c^r9��,lܸ�~����5V�Ҭ����X�W<s }����}���~��3>��S��e%��_���}��GqҀ�^�&��Zi..Z�J*���7��/�p��	'���E�������{J��}��WGw��.:s�����q�
�����"G%_��Q����g��Y::{�ٺ�����w����<k�̾t�����z�T��n_���N�e�U�Zn	ݕ蒇L6q�嗫l�	��jއ��Ds~�	���;Z�j�~���G�����84i�1��:�K)\������{�`ٲ�X�d�.�oS9��Y�|��LO��1ϣm����}݄x�Y�իWc��%�J䤏��ٳ�f�\}�5�����!)Ig ��N:mڼ	ӿ��>�[6m.�WYN�l��?��^�`NUi����{���#��]z���eMM����q���~-[�@���}f��`��ǧ�->��l\���8ѵ{<��Cz\zM����j�ɢ֭�z���];q�}`��i�ԩ���9����ߥ�q�1��+�ak�r���6`�ZD����_�uz���F`�~�+odC��v�����٧vĨĠN|��)�H@�ǲT@Vw�����}�߳|�I'�ŗơO�^���ӫWO�5��s�^��[-Į�;0�����T/5+��e<�L#����g��)Y�p!�'o��᫆����`��0���@T��b-*(�y�ر};�y�/C@��z���xRe�'O���w��4j�	ut'���=m�r����زe�*I�.��{�F���SO���WMIg�}Ʃz+U��s�^�ru2���4���as��2q�i������G��T@/�#�蚢*\����$��z��c\r�˗-��Jg�[��d!�Çӽl��J���0���{�y1�Yt��9 7�9C�F���裏b��M�ԥ��k�v��~�=�UxD�c����<��Ư��M�5�SÇ��T����hеR*0H&2?� ���C�v�m�#遽i�z���˯��uהφ������3#��y�&x��q�X���d������u2
���X|�\������{�a���HP����z�Q^���ß�Rsx��e�^�6mZc��Q�q��ɖ��\+o�:W�L�ÿ��[q��w�I�FKdH��a�����ß��E���^)z����I���ʕ[�ҵ�J܆�63���&%ntlɽ�X}wF??J��ߞ�6�I/k�Mi�W��*�+�[^F���mݦ-�����
�\�����G��X����f
�))ػo��Ŧj�
��k����={b�ĉ��������H�|=�ze��W��SO;��s7�W���$��;g�^Fv�8���-2����U�9�s��:�	���K����ݺu�Čp�3���^��:�=��Ӻ���W^����aZ� X�E�ʻ���=22��q�}�����DU�]N_�#�=���{?v�H��A����HNN>f+\)���ˣ�����?��ުґCf�[�j5������G���!O�[OO[y�5W��s��OH�۽kL��:��x������,l.�H�M���O���O9�]w�^�F&�����^!N����5Z��W�������@�S�Z4���q��^��z�Ksp�	�>����*�e���G~y]lt4n��z=c�dοV���7��~?3��C���
�Q1�ر��Tw���6jРR���Ɏ�{��^�Z���bu<��qD��Is�|��F��}\(oi���9nӦ��=Opv�A�Н�����Ti����õ�K�L���m.���lݲUw�������HH�G�vmq�	'b��A�ӻ7��M�[�*Ty_҃]ޓ�������3�`�?ر}������К�fG�
�mU�\f�2dN:i �={+}��^�[�e�v:�zᜰ��Wmʾ���t�ֽ�LWr��I�V�!5r���֭[�kWu���Ǒ��S�Jur��=�d�%�v��!`��ʔ��{�,�w9���� ̋.׿Es�믎Ӷm�A�Hy�:��2r�sz����9?��ʕ+�����ɽe\
Oa���Eb�D����w.NS%r����Vi�٣�
n9% ��e��/=���tb릮yZڡ��/Sjk���W�\i^�fK��|���i�Oزy3���c��B��Zj3dTP||�����K����]],�J���մNG�s��gC�t�8�3t�;v"y{�^&TƖ������Y���HH�ڵ�PO���5k�\y�W]�fw���[�9��&w���ur�v�Y�F�N�e��Y%#=]�Ws�$*�j��^f��ر:w�W��#d����׫�	Z2���$�뮻���V"""W��+�I���>����QQQ~�ŕ��qϊ]�#>@���S�/�r�p��}e�#������-7�d��|b��+}lԵ�N����6m�ڵk�z��}�����lnn���bս.�=˒��ڵC'��v�{�Z�Z�
��s;��S��w�-kO�\�����S�|��/-�%� _��C�:�����Sqݮ

�����~%'�:u�ѨQC4i�T��1�2�S�
Ԭr�"�W݌�*ˣg����ِ\���5���@$��A)J%J2�Qj�����_��%�o��>�]� C��2w�zߒ ��� ��Ë����}�u�Dӓp�:�ʪ���qU{�o�VD�=��������"�LU}��qq�Q��)�/�I���&=ⳳ���ס�}��$�(:yHf˰�O�H/����r�;P�7��aUu<O�Tc��Q�9��k������΀^)f�K)C�\����b?�w,��#��L�im/��;�hݥ��8��|��8ގ)�ňp�z�����<��58��0K���0�~L��6�@;�\{u�yy�PM����Ni��f7����YB'""
f�S\�[y:�Q�ѝ8�)������^����3�-ӯ6�|v�#""
b���������(�ٝN��ֈ���7=S\�[�,HN�Љ������W~	]�9:����T:v���3M�r'"":�����,�Tn�7+�O"""
�K�ݯ8-%tFt""��d��m�::QPR1����DDDAKW��UBg�8""��e��˝Et""��U�:#:QP���U��8t""�`&U�~lU�?"""
F��ΈNDD�̊��3�)݆ι܉���;��~e/w""�����,�NDD�L��YB'""
jXm�m�DDD��"���������r�z�DDD՞S�r�5""����U*�}�k�r'""
ZR���VN�f,'""
fz�5?7eX'""
V�ߋ�0�'��,�U{�˧2�5?�r�܉�����m�r'""
b��U��DDDA��Nq�����(��~W�Q�b�;Q�Ǚ∈�B g�#""
~�C�˧2�+��^��DDDA���2DDD�ʏ�\�L��NDD���ΨNDD�����*w""���*w""�`�ʝ��(p�8""����kb=S+'�܉��B ;�U\m������K�p.w""�����\�DDD���X�U�DDDA��Q��LqDDD!����,DDD�*�˝m�DDDA�ɉe�������CgX'""
R�
T�Q�͉e���B��m�&�܉������6t"""
F�U��Gk��DDD����܉����
t�#""�`���WЉ����Dh�m��(񃈈���aT$��UBw8�HKK�!�p���� �`PS
Q���c�=�l����j���둓��ז�n��0l�C��Wæ�5�������]8
�������p����*�&6���e��-�8\yS~U��^�t1����h2�g�.��6��sDDDt�I��f4��&��� ""��JJ�:�烈���+UB7��͖n:�� ""��Hfsأ��ege�U;6�-3:::�^�n��������{�g��0=""�I&������K���;w$�Өqӻ<�t^^^/�4cTD��u�ƪ�3*8���c:1ϑ��g�#|���g��OF��x���$�����jժ�y�����W�<l��k�ŧ�O����;v����LP�F��]mn�G���E��l6�&m�v��0�æ�`ap�4�����rd��ϫXf��Ta���
�+����ſ�F�_JoWl����l�	�Q�k1׉x����󇢿B�8*�g�J����b{/���}����(:f��Qxn(���.u��{�`[�~���0T�.b�ҥ�{v�
/���G���NC�&M�T�^n7TWr�֬Y����[f�������=��ILl�o�Nɟ�f��MX�<[Q��}y�~����1�\4%�Y�wϮ�����,�{������vW��3K���yxv�c?%�l�Kb�R��\��W���)|q9��,q%��[����ĮK��}���n�a���{��_�]�r)�'�z_/)���N�l�b+��(�-6-�Y�b����J�-��ڨ�9��G�}{ΧԖ����t��pJ�e���%���-:�b�G�J�JM����.rџ�ݠ��:IϹ��\�������0̘�hg|BvIIs�����Saw���ʇ���G4�΅�Ϡ ?W?j"�gY"P������Ӑ@�p��ÐB�l�S�t8W pr�����T$u:�Õ��p?����w���&���\]$�b��$�o�^ܙ���kѾ����m6�����u�]o�ٽ�ً\t�Ÿ��[Bnn�;z��͸�λt"Q���N���on���'�<�������OOL�<O�EyUw�g��&�%�f�L������õ�Y�I�?\���u����hY<u���	S�,�;u):/��s�]6
ӛb�r�����
_��G���R�����̰�^����kc��4�ͦs�6Wy��-5�0�\�����6�]^cs[�e�._�CA��o��0RB�zHٿo��>�S?�� O�l٪UH��7�

���Vtx�is8t��4��J4�m�j��m�w��/�(5�_�O!_ega2�J%J��#��X�]<�g�إ{�i�'6�^�٧�Lexb�Y��Z�;�'���|��������Jl��2y�.�-�܌Ȉ��Zu#WD ��x���\���j�ژ��~̯s~Y߿}���E���[_a��p�2�mW|�ҥ�R��(�P�F�s+��(��/��(]�*��2�M��x�k�9��?ós�t�<�t�B�{��#�?=�Og^�{Tx6�k��F��'�����ܙ��r����w��=��M\�C���x�y0e[��|�}������vU��2��pU"R��Ɂ�
��c8�Զ��r���گ�S������r�Jt�ܹ�ug����e�,���o��� ����W;����"�#

�eF���e���سgZ6o�/S�T婌���o�c��-]:�mҬ�ks�u���'`��u���+AD,Щ���T<�$$$����J��ʬWr[�l���kt@�`.�;���*CS���f�^��?�>��t��6��{�Q0a@�2ڷh�ǞxR�����v��V&����a�?�`��A�>������_<��sػG��R���Jn߱ø���vh�] "
F�d�q�&�ݧw�_|�^�ڵ����������:��m;����x�駱j�
������f͚���/s�~y��6�w�� "
6�d)-��p|n���V���]*�J[�j5�nۊݺ�:ҝ���1f��y�l�i80ԫW��O>��/��Lꐄ�cǂ�(1���N�#:&f�
�y*�G��¦;�-Y��������λ����(�	N����h׾ݘO?�$%'�0���:Y�6�6m�ʔ���#���5*�M^n6����\s"��Q����{���K���@��0�=�Q��o��}�'�?�fM��;�"�`ŀN�.��b\{��6�#""|Wf��Ȫ/���K����^�jӎ.�bي�1b$��މ��\�����g��w�;��>�Y'>�G<"�`ƀN^����۴9�����U��Uv[�n����t@�$������ѣ�d�b�	�JtTTr��-�L�655/;DD�:y����`r�ڴi�Ff�*;ͫ��b�e8���Q���㭉1��o`5���W��k�.���� �n��O?"�`ǀN^}�~.����j���s�yyQ��q8�p�"���"*22��g��oLx��ٰ*�׊��ѭG��Np�����޻o���:`@'��M�ݺ�@TT�&e~^nS�v�U+Wb_J
Z4k�`�i75r����`��y���ϛ�����C��޻Љ��`@'��z�\vŕ��Ď�QQ۳27-���m۶bÆ�A�u��~w��b�vs�ݞݰA��+W,[8��G�Գ;n��jU��S߾}p�ק�<{�Z〭�%�:tK�.����`$����˒�����|�)�ߓ���mxi� "�N�ɧ����
���e�Ͷ��뻗�t`ѢE��ɑ�AՎ.'+��'�h7���]ٮ}����-c��� "���ɧ_�͚�D�:�W���g��^�j;iG߻oZ�h�`�״����p���n7���hܴ�����)_}��K�aԨ "�n�ɧ��.B�=l˚ի����Xt��۱~���	��SRS1z��^Ǜ6�,����\�պ�k0�|���K "��Щ\	uиq�ݪ�%=-�M�-����y��y�5�fϓv�I����v��:uz��/�ʱ���)�����b@�ru��I��9�U�a�Q�c�t`������Flt�1oG�v�7&L���[��#���7o�r�/?��y���ؽsN?�tUW�T.w�8�{�^�򚣠� �j�U+Wa�޽hӪ��x�#Gc��vsy6���s�͜�����O��3O���:c@�r͚5]��@|B����������e���ؾ�֭?f��<�`�E���_{�����/���w'OQuǀN�:��q�7�t:��/]�+++�n٭����v��:��(���y�EtL̎�mڌ�����0 ��Qv;"����_�z����/��?x�`�mLӡ�S���BlL�QoG�����7����`n���7i������3#����`ND!���Ҹi�rӍ��:���l��]y�e���ػwڴnu��MB�Ju\�j߻w,�����P��'�<��AC�1۶m��oL Q�`@'�<��Ø��iG_�J�9y+�Ihݹs'�o�p��������`���n��]�v�g�������q��_3�QHa@'�HǸ�I���Y����J,�v�e˖��AgU�9I0�/(��＋iS�I�?����#�7i����[2���ѳ[Q#��ÀN~��q=��t"۵�߅�2�3,�V3��ѳ��sƣ�4�g���k��΄U����s/�`J��]�v�Z<x߽ "
5���m����n94��S��`5��X�z��KA�U3�g��u6�y�w��˪vUX��]��Ν;��釙Y���� "
E����Cҹ�ٳW��av�� ?�2��x�M7VY@��JO�ر�������n�ڢeˑsf��)�a��_����Q(b@'�=8t(>��+ԩS{UDDxFA~^�	f��Ұt�2�y��*9��~�?|���0M'���e6���Mz��W�r�x���0⹧AD���o���Z�i���M��ѻ�23�Xm�׽*�G����ܹxy����̀uU���s���Mxz�3�5�[��ND!���ֿ�?^Ƥ����/������m�5�Wc_J
Z6o��K0߲u+F��m[7���m�ڷ����{�r���_���?Q(c@�
9����1))�s�n+m6���Hޖ�M�6,�K0����K/��彩�-�����4m�t��?��9���дi\q� "
u�T!��ɨ];			K#""rsrr"�n�jG_�l�vj@��0M|��g���>���U��a��~�ĩ���K/3���1�Y��Q���N2��3q�"22r}dT�����&V������%K�������J������k>^�"2��[���ۻ��*�<��?�����n4$kBGMk׭�bv�r�s'k7��f�v�Y�j^Rlk�Uh3#l[��dE!0�&"��*'8��e7��s�[�<|?3g8����w��9���L����ܶ�3� ���~�>*J���k������%��8m�F�Y�Dz򃴘מ���5k��\���G�|}[Ǎ�� ���T�|~�3y��' ���~�6�f��ҥm�3�t��_`�Kjj���ٳ
����Z:;e}F��������zWxDĎ�~����
� ?_�n� �pB��oK�zJ[`ƞp�m%��e����A�%-�-RRR"���;�jQ��y_v��]v�����	:���cGW@@���1��v:��Ç%.>ABCCK||}�m6k�����V)*:!]6�x�}:��W���Xa��MY+��f�����	�����Z�N��M*{��:�m������gŠ7T;v��J{{���_�|%M�&�w����74HRR��*+�^Q���ᆌ=|��W^����አc@�B�d��Sr?ʭ���0�Ӹ��*����	z_h1���ƍ�$���<��
�?w�?����/�k� W29�$��ϲ.%��*�~���p3J�su^ZZ*�Ϝ��s�ݷW�l�"6�U<͛�Un���o�ަ��RXX(��� �pE�1 ?��DG��M�'����X-���q6[�?^$֧�b4��禥�Dq�$'�H���t�����=>�Ճ���; �.\���x�ጠc@���f�~��������k�X:�=]Mk����-�q];��,)�k�d�	����N'QQQ{�WO�?c��v����+ �;��������L1u�
�k/{�$?w��������&[�n�?�#�}��Z!�!E3�e���hjn�m��  A� ����c�>bޙ�uZ���{ڨ���(��e2c�t���ҝ��'37HW�7ڢ�r�K�Z~:yrʮ���t�3R[^..  A� DDE�,0��_�Sl��~�����(/���EEb�Q����{W���%yM����Iϭv7��Fo׍��;�צ~x�;��Ȋ�� �_6w�,���Hxxx�ȑ#-�W�~�o�����XZ��亠����F6��Jj�:���/�Ӽ���ZdT�;�ߙ�>����%9�� �w:L�"uz\����-��dn�����R[S��o����)ٻ����i��%A����3��^{�g5���*� �C�1`�G����>Ѿ^��Ω����t��_� {��S�Iz}O���]��.�X����s����s�bc7�d��ߕ�P�1���y� ��:eF|��
h	)3��6���8m]��۷K��Y2g�,�8wN��$u_�WK/��i���_�Т7W�|�.�,~H  �"���ks��y��t����ߔNj��%=-]���$c}�=rD<=��]�GFF��=gv�ƍ�N����
 �cP^߲E��#gΜ)�;엺�����򤪲J*����Ԗ�u?o8j��֙�fnX���g�!�>yR  �t��%�n�Nʻ�|\z��t~�)�'��MR�e���i�L�]���훶lq���ɯ�<)  �:�d2ɒ����������ں��tz�~���w'L�X}Ͻ��ݺu���ݻD�d;A��tZ��J�:m��/>q����ā��%�GZܽ s�����j��u�̝@t�'��˧G���;�x�iʦ���X�V����`0J\|\ުU�v,8䊈���� �aC��?��{\Ǝ���?���b}�.�K��`4��W�Ǜ��j����pF�1$��^��:f츎�G������q���>��K:�n[xT��i�ؤ���[� �Cf�Ν��ޮm�r�������T����C�i�+��<�����-�  ����2˖,��/���s�J�ط���w���-���*<!!��]wߕ|������� }G�1���ِ������l�X��m�I=��������3>m�^9��ŕ���*/���  ���cH͙3Gv��-oeeɁ��"_�$�ݑ�]�Qn���z�;f�y��g�9��ӈ9 Aǐ[�x��d2���D����t:&8�UN���|�����`4�1��Eǋ���ʤ��V  C��8UZ*:�QBCB�'LL375�X::��lA:�����'wtp��u��wZ,�z�j1M�$ ��!���86ih��^��������dn�:V: `�:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
�O��Ր���    IEND�B`�PK
     ^�[��EM  M  /   images/d3694a2e-5bba-40c3-8069-8db85c4c9209.png�PNG

   IHDR   d   d   p�T  TiCCPICC Profile  x�c``RI,(�aa``��+)
rwR���R`����b
����>@%0|����/��:%5�I�^��b��Ջ�D������d ��S��JS�l����):
Ȟb�C�@�$�XMH�3�}�VH�H�����IBOGbC�n��ₜ�J� c���Ԋ�_PY���Q���Tϼd=#CsP�CT�%���X�}�����ߍ�������k'BLÂ�A�����΂ĢD�33��10|Z����� |�'�8��,������z����j��N��������.j���p  !e�2���   	pHYs  %  %IR$�   xeXIfII*            (           J       R   i�    Z       %     %      �    o  �           a���  �zTXtRaw profile type icc  x��S[n�0��)z^�8~$R��b;^eW�J�ё"�@`H�n-|DI�D��@ȴ�v=L�"�	�s,`�ۮ��z����"H����pz����3�ͬ,9&�h'�tN9#���(���d>CQ�h�|q�k��R�R����mOi�q�6�Z�ܶ=���C�>hrK$>���U`�͚t3�s;����%�S�T�c��\���~�y§b�_"%�G"a=}J�H����|)�Ni����2��yl�c���r�E��|�7$��8��s���.PJ����
��wq�8��P'��j����[ܞ�c2����g�+��|����RM�=�c2gҥl��ϞauTh���҈�\�z���줡㜥   %tEXtdate:create 2020-01-31T21:31:09+00:00��y{   %tEXtdate:modify 2020-01-31T21:31:00+00:00	�   tEXtexif:ExifOffset 90Y�ޛ   tEXtexif:PixelXDimension 1391c�   tEXtexif:PixelYDimension 800�요   (tEXticc:copyright Copyright Apple Inc., 2017���   tEXticc:description Display P3�y��  cIDATx��]	xLW~��d�(%�J"��}�%(�Z���B��_[y~R�R[u�E[[����J����ҿZ��j��B)��'s��;��Ĉ����>���=��s�s��-�37:�PTB��A%DaP	QTB��A%DaP	QTB��A%DaP	QTB��A%DaP	QTB��AW÷&��z\I���7�)I*�Ev�Z�:d;iJ�3mtRɲ�������V�$IY6��"a[�d��$}/����~�l���99��t.��$u0Z��d�M��(��5D��a�}0�*�
��?���h��dY~�`ȫq+��L��yY���@���[���������ƍ����0��`�Aк�C��"�|<B&�������r����t�PQ:�;w'N�{˧����a)y���3�t>���ʂ
E@fB\yyP� �f�3b�1�(p�3!�<ÃY=��䫄(�d���?0��&1A3vH�JIi�	�YCd��c,�p?��0���g�Ж���lqtws���%b�G��ɒ�2d'jaxR�v�Zl߈s��S�����_C���2Js;�i���8�f�ɒM>�Q.]�����С�x�g/�5J<����зO̚=�g����f6.:6lX�t]������B��5�D��;ѽ[7���s�p�0g�,�n�=_x��(���E��~/���u{���F�m�6�2�h��!����v����;����dX�i5�7�}�����ٿ�2~޳?��#n������1p�@xV�$��u˖�Ѳe��H�zi��|��u��,�Ν'�����ԩ3�/�5PP��7o���,�_���C�޽ѵK���ǚ5k�t�:>�,^|q 4�XȺ����7!&&�+{�_�~��d��ǎ	SԥkW�o؀������A��n��B�p2�7n����Na��>$3��ARLN�G��&����~�� �����QQ��wq�������Тe+xU�ºu_ lQ������͐�լ�K�.����ԙK�.��9����(�QN4|���X�p&M|�����5�OLLDu��x�"�.Y�9o��&�l7ww7�b�rD�c�)��?��޽E��jO����[���a�0�?B��ۿr6n����o�Y�}��E�E�:uh@lAZZ*�i`5]�ر�u�9Ǻ��<s�4�V���ի۽��1�Q�n�:AƢ����D�?O�F�g:b����a� i4puuÑ�#������W��u� ̜�iL8^<H�Ȏ��ʕ+Bui������®�v�u�zS����u>l�ФΝ�P�U�@.��+��������^M�5c�L�L��S��nW",�Y��e��'""#�|���'B�B�FMТœ8���	�R��ӓC��w��t�b�_G�R׿ƛG߭~=L�6U��?���קў��ݻ[��Z���\�rLd0�q�	��o@Ey.D<kI��
2^U��~�zB�!C^65V�E�6m�W���$!-^�j� ��溃��������͂�٤������m׮j׮����{��l"��e����G�fg�AQ�%{ΫbM�6��F�흚6m"�.\@�ƍD���]P��	��g�ΕG���e?h�V��\��ӊ�����ٳq"m���`1i.�[8c:fd��Y����<P��6���׻�2�sq�{dDG2kd'j	h�͛��)2;U�jW��%�=z|j���)�b~b����!JcӁ�L��+$3�i��ߪ[�Fc�8����2�F����~~���dG��?��%\�9���ɡ���3lw[wGDD���Ç�6�V�Z8AQ?��6U_"���YԢq�0��$��_M�i������W[P��@�nns+�F*Z��@'����!����ǤI��`�<a�CI�>��p������<*T�[�Cɩ�1K�,>�>}�/�h�M�vhD�*��89�-�aq�֭�M0m�t�jQt������5k?C��M�ۻ�Mk5���Z�e����ZSVY'�����L���������'����F����g(4�Ŷ��P�^G�>|<(��p������_�R�VUDK</`9rr��WhI�6��E^��9��~��΁�ʧ(��K�c��K�^���}Ѭis<���b�s���J�efp �e
���,���5��<�5o۶oD��h���%.�sab��F��%a�ȑ4I܍��u�Ȗ-�!00�==̤?�9@���������A��"���K�T����J��2
�������r�̋h���C�Шn+���\�t	�i~`�'t�dA�����Ӄ|�'���GEDCQ��z�5{zP�gA`�@��?�h����\�h*��5���]�r^^^pbb(��1��[ޒbo�ػ^8�s4�叽|�4�@����4}�#0(h�my
?A�#����Mg�<��7��?�il���_ �2Eto�����"����j�37-N^��4g��)�8����&��'�*JBCLQ�JH�C���=d��,���}X5D�2`�����0��g窆(&Q#,���!�.o���e�TF��[���9ʲIQ�[�<l�M�V��|/="D�xOR���vG�_G�3˚��7��aj�gE��s�6��ˋk�Q'I����܊�GBEiB���j���QCG�h4Z�D�$ݢY�-R��By%�V+i�T���I|3����4����ĉؙ}���2r����)���Om�fk\]�zH�|�R�iO�l�Mۗ�I6_dْϜf4G��Fk-匷�ݥe�k�\𛍶���V���_�3���X:�-�b(ڴ#ݾ���KĤ����h$�v!VI~}��+s�^����xg��p�h4"�E@�Ӈ$^N������1���	�����ǁ=j��������o��qbZW�?��i�1��wI�t�G��v��e��^3�x޹���k+�t�w��`-;q<3��rJ�r�##���Κr$55G��޶;�a�±c_�ٿΜ�V�{J9�Ԕd��=�(B���}�\�.1�7����׭w�^v�.\�[��"{x<����̣������{�"o���]�|ҵ�"#��[v��n�ٻoޚ>�Mۢ�̛;[�A���(Ks�#�����@�V�s��I������׸��������gn�fV��8\��@�*e	%F��#�n�����8v� �2�Ǎƙ3�2+yV{<6���ܜ����#d9�¡��ȏ ""�z�ז-_�M���^nzjJ�QNk��i�܇��#��~_�Z(_��?���&��2�G9��ɡ�=�gge|�yx�fY$�Q�/R~�'������ll���<����� ~�N�z�����t
s�PVQ��<^�q�s��mOrrJ@�=�t-���K		粲24x6�;�;�%JHJJ
*�|D��-KKMN!p5�olI�x��ݺ�Ge�F��kǏ�H�"A�ռ!i\�xzz�/_�<�R�u�7�u�����U�F��K0��N�rx����̬L�(B���^b���x:y9��}���E������k��%u����QTB��A%DaP	QTB��A%DaP	QTB��A%DaP	QTB��A%DaP	QTB����Blg���    IEND�B`�PK 
     ^�[;�9:�  :�                   cirkitFile.jsonPK 
     ^�[                        g�  jsons/PK 
     ^�[B�@\�'  �'               ��  jsons/user_defined.jsonPK 
     ^�[                        z�  images/PK 
     ^�[�:��� �� /             ��  images/c7631ad6-ed21-46e6-964c-e953ba5165ac.pngPK 
     ^�[�AWv�'  �'  /             �� images/97fe1122-b934-4e82-b9ff-450ac31bc7af.pngPK 
     ^�[x^��_� _� /             � images/d5d3b89f-59ab-4c38-95f7-2948dd30f8f5.pngPK 
     ^�[/�i�$  �$  /             +r images/60da03ea-f7cc-456a-983c-41a209708cd9.pngPK 
     ^�[��
�G2  G2  /             � images/ee130f24-d674-430f-bd58-6b2b8a983a65.pngPK 
     ^�[��Vt�  �  /             �� images/193bec7f-e59d-4bcf-b15c-6ea8617b7acc.pngPK 
     ^�[	��} } /             �� images/bbfae99c-8036-4c5e-89fd-a87441410720.pngPK 
     ^�[d��   �   /             "` images/a262aa33-74c4-460b-b0ad-c746896f6744.pngPK 
     ^�[�c��f  �f  /             �� images/c88b2895-5e8b-4a57-9f9a-b80dd50058b1.pngPK 
     ^�[��EM  M  /             (� images/d3694a2e-5bba-40c3-8069-8db85c4c9209.pngPK      �  ��   