PK
     8p�[_6c�  c�     cirkitFile.json{"raven_core_version":15,"hardware_version":0,"pin_to_graph":{"pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_0_0":[],"pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_1_0":["pin-type-component_18c68858-ce98-4365-aa62-ff9cecd47749_2","pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_0_15"],"pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_0_1":[],"pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_1_1":["pin-type-component_18c68858-ce98-4365-aa62-ff9cecd47749_1","pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_0_16"],"pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_0_2":[],"pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_1_2":["pin-type-component_18c68858-ce98-4365-aa62-ff9cecd47749_0","pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_6"],"pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_0_3":[],"pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_1_3":[],"pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_0_4":[],"pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_1_4":[],"pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_0_5":[],"pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_1_5":[],"pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_0_6":[],"pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_1_6":[],"pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_0_7":[],"pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_1_7":[],"pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_0_8":[],"pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_1_8":[],"pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_0_9":[],"pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_1_9":[],"pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_0_10":[],"pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_1_10":[],"pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_0_11":[],"pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_1_11":[],"pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_0_12":[],"pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_1_12":[],"pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_0_13":[],"pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_1_13":[],"pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_0_14":[],"pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_1_14":["pin-type-component_19abf22e-c985-43dc-b307-bec227e65f21_0","pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_5"],"pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_0_15":["pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_38","pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_1_16","pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_1_0"],"pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_1_15":["pin-type-component_19abf22e-c985-43dc-b307-bec227e65f21_1","pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_0_16"],"pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_0_16":["pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_37","pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_1_1","pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_1_15"],"pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_1_16":["pin-type-component_19abf22e-c985-43dc-b307-bec227e65f21_2","pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_0_15"],"pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_0":[],"pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_1":[],"pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_2":[],"pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_3":[],"pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_4":[],"pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_5":["pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_1_14"],"pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_6":["pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_1_2"],"pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_7":[],"pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_8":[],"pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_10":[],"pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_11":[],"pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_12":[],"pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_13":[],"pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_14":[],"pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_16":[],"pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_18":[],"pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_19":[],"pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_20":[],"pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_21":[],"pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_22":[],"pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_23":[],"pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_24":[],"pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_25":[],"pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_27":[],"pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_28":[],"pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_29":[],"pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_30":[],"pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_31":[],"pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_32":[],"pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_33":[],"pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_34":[],"pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_35":[],"pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_36":[],"pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_37":["pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_0_16"],"pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_38":["pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_0_15"],"pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_39":[],"pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_40":[],"pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_41":[],"pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_15":[],"pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_17":[],"pin-type-component_19abf22e-c985-43dc-b307-bec227e65f21_0":["pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_1_14"],"pin-type-component_19abf22e-c985-43dc-b307-bec227e65f21_1":["pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_1_15"],"pin-type-component_19abf22e-c985-43dc-b307-bec227e65f21_2":["pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_1_16"],"pin-type-component_18c68858-ce98-4365-aa62-ff9cecd47749_0":["pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_1_2"],"pin-type-component_18c68858-ce98-4365-aa62-ff9cecd47749_1":["pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_1_1"],"pin-type-component_18c68858-ce98-4365-aa62-ff9cecd47749_2":["pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_1_0"]},"pin_to_color":{"pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_0_0":"#000000","pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_1_0":"#9929bd","pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_0_1":"#000000","pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_1_1":"#000000","pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_0_2":"#000000","pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_1_2":"#e32400","pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_0_3":"#000000","pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_1_3":"#000000","pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_0_4":"#000000","pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_1_4":"#000000","pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_0_5":"#000000","pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_1_5":"#000000","pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_0_6":"#000000","pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_1_6":"#000000","pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_0_7":"#000000","pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_1_7":"#000000","pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_0_8":"#000000","pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_1_8":"#000000","pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_0_9":"#000000","pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_1_9":"#000000","pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_0_10":"#000000","pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_1_10":"#000000","pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_0_11":"#000000","pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_1_11":"#000000","pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_0_12":"#000000","pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_1_12":"#000000","pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_0_13":"#000000","pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_1_13":"#000000","pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_0_14":"#000000","pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_1_14":"#ff9300","pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_0_15":"#9929bd","pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_1_15":"#000000","pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_0_16":"#000000","pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_1_16":"#9929bd","pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_0":"#000000","pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_1":"#000000","pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_2":"#000000","pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_3":"#000000","pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_4":"#000000","pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_5":"#ff9300","pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_6":"#e32400","pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_7":"#000000","pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_8":"#000000","pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_10":"#000000","pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_11":"#000000","pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_12":"#000000","pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_13":"#000000","pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_14":"#000000","pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_16":"#000000","pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_18":"#000000","pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_19":"#000000","pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_20":"#000000","pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_21":"#000000","pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_22":"#000000","pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_23":"#000000","pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_24":"#000000","pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_25":"#000000","pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_27":"#000000","pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_28":"#000000","pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_29":"#000000","pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_30":"#000000","pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_31":"#000000","pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_32":"#000000","pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_33":"#000000","pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_34":"#000000","pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_35":"#000000","pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_36":"#000000","pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_37":"#000000","pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_38":"#9929bd","pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_39":"#000000","pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_40":"#000000","pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_41":"#000000","pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_15":"#000000","pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_17":"#000000","pin-type-component_19abf22e-c985-43dc-b307-bec227e65f21_0":"#ff9300","pin-type-component_19abf22e-c985-43dc-b307-bec227e65f21_1":"#000000","pin-type-component_19abf22e-c985-43dc-b307-bec227e65f21_2":"#9929bd","pin-type-component_18c68858-ce98-4365-aa62-ff9cecd47749_0":"#e32400","pin-type-component_18c68858-ce98-4365-aa62-ff9cecd47749_1":"#000000","pin-type-component_18c68858-ce98-4365-aa62-ff9cecd47749_2":"#9929bd"},"pin_to_state":{"pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_0_0":"neutral","pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_1_0":"neutral","pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_0_1":"neutral","pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_1_1":"neutral","pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_0_2":"neutral","pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_1_2":"neutral","pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_0_3":"neutral","pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_1_3":"neutral","pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_0_4":"neutral","pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_1_4":"neutral","pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_0_5":"neutral","pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_1_5":"neutral","pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_0_6":"neutral","pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_1_6":"neutral","pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_0_7":"neutral","pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_1_7":"neutral","pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_0_8":"neutral","pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_1_8":"neutral","pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_0_9":"neutral","pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_1_9":"neutral","pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_0_10":"neutral","pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_1_10":"neutral","pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_0_11":"neutral","pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_1_11":"neutral","pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_0_12":"neutral","pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_1_12":"neutral","pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_0_13":"neutral","pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_1_13":"neutral","pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_0_14":"neutral","pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_1_14":"neutral","pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_0_15":"neutral","pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_1_15":"neutral","pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_0_16":"neutral","pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_1_16":"neutral","pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_0":"neutral","pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_1":"neutral","pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_2":"neutral","pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_3":"neutral","pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_4":"neutral","pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_5":"neutral","pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_6":"neutral","pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_7":"neutral","pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_8":"neutral","pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_10":"neutral","pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_11":"neutral","pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_12":"neutral","pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_13":"neutral","pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_14":"neutral","pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_16":"neutral","pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_18":"neutral","pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_19":"neutral","pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_20":"neutral","pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_21":"neutral","pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_22":"neutral","pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_23":"neutral","pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_24":"neutral","pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_25":"neutral","pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_27":"neutral","pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_28":"neutral","pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_29":"neutral","pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_30":"neutral","pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_31":"neutral","pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_32":"neutral","pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_33":"neutral","pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_34":"neutral","pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_35":"neutral","pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_36":"neutral","pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_37":"neutral","pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_38":"neutral","pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_39":"neutral","pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_40":"neutral","pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_41":"neutral","pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_15":"neutral","pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_17":"neutral","pin-type-component_19abf22e-c985-43dc-b307-bec227e65f21_0":"neutral","pin-type-component_19abf22e-c985-43dc-b307-bec227e65f21_1":"neutral","pin-type-component_19abf22e-c985-43dc-b307-bec227e65f21_2":"neutral","pin-type-component_18c68858-ce98-4365-aa62-ff9cecd47749_0":"neutral","pin-type-component_18c68858-ce98-4365-aa62-ff9cecd47749_1":"neutral","pin-type-component_18c68858-ce98-4365-aa62-ff9cecd47749_2":"neutral"},"next_color_idx":9,"wires_placed_in_order":[["pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_38","pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_0_15"],["pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_37","pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_0_16"],["pin-type-component_19abf22e-c985-43dc-b307-bec227e65f21_2","pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_1_16"],["pin-type-component_19abf22e-c985-43dc-b307-bec227e65f21_1","pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_1_15"],["pin-type-component_19abf22e-c985-43dc-b307-bec227e65f21_0","pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_1_14"],["pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_0_15","pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_1_16"],["pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_0_15","pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_1_16"],["pin-type-component_18c68858-ce98-4365-aa62-ff9cecd47749_2","pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_1_0"],["pin-type-component_18c68858-ce98-4365-aa62-ff9cecd47749_1","pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_1_1"],["pin-type-component_18c68858-ce98-4365-aa62-ff9cecd47749_0","pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_1_2"],["pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_0_15","pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_1_0"],["pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_0_16","pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_1_1"],["pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_0_16","pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_1_15"],["pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_1_14","pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_5"],["pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_1_2","pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_6"]],"wires_removed_and_placed_in_order":[[[],[["pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_38","pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_0_15"]]],[[],[["pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_37","pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_0_16"]]],[[],[["pin-type-component_19abf22e-c985-43dc-b307-bec227e65f21_2","pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_1_16"]]],[[],[["pin-type-component_19abf22e-c985-43dc-b307-bec227e65f21_1","pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_1_15"]]],[[],[["pin-type-component_19abf22e-c985-43dc-b307-bec227e65f21_0","pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_1_14"]]],[[],[["pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_0_15","pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_1_16"]]],[[["pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_0_15","pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_1_16"]],[]],[[],[["pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_0_15","pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_1_16"]]],[[],[["pin-type-component_18c68858-ce98-4365-aa62-ff9cecd47749_2","pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_1_0"]]],[[],[["pin-type-component_18c68858-ce98-4365-aa62-ff9cecd47749_1","pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_1_1"]]],[[],[["pin-type-component_18c68858-ce98-4365-aa62-ff9cecd47749_0","pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_1_2"]]],[[],[["pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_0_15","pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_1_0"]]],[[],[["pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_0_16","pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_1_1"]]],[[],[["pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_0_16","pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_1_15"]]],[[],[["pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_1_14","pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_5"]]],[[],[["pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_1_2","pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_6"]]]],"arduino_state":"arduino_off","pin_to_uid":{"pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_0_0":"_","pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_1_0":"0000000000000000","pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_0_1":"_","pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_1_1":"0000000000000001","pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_0_2":"_","pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_1_2":"0000000000000006","pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_0_3":"_","pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_1_3":"_","pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_0_4":"_","pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_1_4":"_","pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_0_5":"_","pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_1_5":"_","pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_0_6":"_","pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_1_6":"_","pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_0_7":"_","pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_1_7":"_","pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_0_8":"_","pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_1_8":"_","pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_0_9":"_","pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_1_9":"_","pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_0_10":"_","pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_1_10":"_","pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_0_11":"_","pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_1_11":"_","pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_0_12":"_","pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_1_12":"_","pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_0_13":"_","pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_1_13":"_","pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_0_14":"_","pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_1_14":"0000000000000004","pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_0_15":"0000000000000000","pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_1_15":"0000000000000001","pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_0_16":"0000000000000001","pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_1_16":"0000000000000000","pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_0":"_","pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_1":"_","pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_2":"_","pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_3":"_","pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_4":"_","pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_5":"0000000000000004","pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_6":"0000000000000006","pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_7":"_","pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_8":"_","pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_10":"_","pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_11":"_","pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_12":"_","pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_13":"_","pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_14":"_","pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_16":"_","pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_18":"_","pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_19":"_","pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_20":"_","pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_21":"_","pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_22":"_","pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_23":"_","pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_24":"_","pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_25":"_","pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_27":"_","pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_28":"_","pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_29":"_","pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_30":"_","pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_31":"_","pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_32":"_","pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_33":"_","pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_34":"_","pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_35":"_","pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_36":"_","pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_37":"0000000000000001","pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_38":"0000000000000000","pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_39":"_","pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_40":"_","pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_41":"_","pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_15":"_","pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_17":"_","pin-type-component_19abf22e-c985-43dc-b307-bec227e65f21_0":"0000000000000004","pin-type-component_19abf22e-c985-43dc-b307-bec227e65f21_1":"0000000000000001","pin-type-component_19abf22e-c985-43dc-b307-bec227e65f21_2":"0000000000000000","pin-type-component_18c68858-ce98-4365-aa62-ff9cecd47749_0":"0000000000000006","pin-type-component_18c68858-ce98-4365-aa62-ff9cecd47749_1":"0000000000000001","pin-type-component_18c68858-ce98-4365-aa62-ff9cecd47749_2":"0000000000000000"},"component_id_to_pins":{"9ed9f913-4687-4140-b5ca-f53cf9998566":["0","1","2","3","4","5","6","7","8","10","11","12","13","14","16","18","19","20","21","22","23","24","25","27","28","29","30","31","32","33","34","35","36","37","38","39","40","41","15","17"],"19abf22e-c985-43dc-b307-bec227e65f21":["0","1","2"],"18c68858-ce98-4365-aa62-ff9cecd47749":["0","1","2"],"9d530ea4-6449-4e29-a81e-6c2c23ffcdbe":[]},"uid_to_net":{"_":[],"0000000000000000":["pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_0_15","pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_1_0","pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_1_16","pin-type-component_18c68858-ce98-4365-aa62-ff9cecd47749_2","pin-type-component_19abf22e-c985-43dc-b307-bec227e65f21_2","pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_38"],"0000000000000001":["pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_0_16","pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_1_1","pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_1_15","pin-type-component_18c68858-ce98-4365-aa62-ff9cecd47749_1","pin-type-component_19abf22e-c985-43dc-b307-bec227e65f21_1","pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_37"],"0000000000000004":["pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_1_14","pin-type-component_19abf22e-c985-43dc-b307-bec227e65f21_0","pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_5"],"0000000000000006":["pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_1_2","pin-type-component_18c68858-ce98-4365-aa62-ff9cecd47749_0","pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_6"]},"uid_to_text_label":{"0000000000000000":"Net 0","0000000000000001":"Net 1","0000000000000004":"Net 4","0000000000000006":"Net 6"},"all_breadboard_info_list":["37073b3b-134f-45d6-97fb-5c4c86637137_17_2_False_663.0000000000002_348.0000000000002_right"],"breadboard_info_list":["37073b3b-134f-45d6-97fb-5c4c86637137_17_2_False_663.0000000000002_348.0000000000002_right"],"componentsData":[{"compProperties":{"mpn":{"version":2,"id":"mpn","label":"mpn","description":"","units":"","type":"string","value":"RPI3-MODB-16GB-NOOBS","displayFormat":"input","showOnComp":false,"isVisibleToUser":false,"name":"mpn","unit":"","userVisible":false,"required":true},"manufacturer":{"version":2,"id":"manufacturer","label":"manufacturer","description":"","units":"","type":"string","value":"Raspberry Pi","displayFormat":"input","showOnComp":false,"isVisibleToUser":false,"name":"manufacturer","unit":"","userVisible":false,"required":true}},"position":[1199.31025,375.44717],"typeId":"b739cbaf-bacb-4ee2-abf3-78459baee6db","componentVersion":1,"instanceId":"9ed9f913-4687-4140-b5ca-f53cf9998566","orientation":"up","circleData":[[992.5,230.00000000000003],[1007.5,230.00000000000003],[1022.5,230.00000000000003],[1037.5,230.00000000000003],[1052.5,230.00000000000003],[1067.5,230.00000000000003],[1082.5,230.00000000000003],[1097.5,230.00000000000003],[1112.5,230.00000000000003],[1142.5,230.00000000000003],[1157.5,230.00000000000003],[1172.5,230.00000000000003],[1187.5,230.00000000000003],[1202.5,230.00000000000003],[1232.5,230.00000000000003],[1262.5,230.00000000000003],[1277.5,230.00000000000003],[1277.5,215.00000000000003],[1262.5,215.00000000000003],[1247.5,215.00000000000003],[1232.5,215.00000000000003],[1217.5,215.00000000000003],[1202.5,215.00000000000003],[1172.5,215.00000000000003],[1157.5,215.00000000000003],[1142.5,215.00000000000003],[1127.5,215.00000000000003],[1112.5,215.00000000000003],[1097.5,215.00000000000003],[1082.5,215.00000000000003],[1067.5,215.00000000000003],[1052.5,215.00000000000003],[1037.5,215.00000000000003],[1022.5,215.00000000000003],[1007.5,215.00000000000003],[992.5,215.00000000000003],[1127.5,230.00000000000003],[1187.5,215.00000000000003],[1217.5,230.00000000000003],[1247.5,230.00000000000003]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[749.078923,885.6579214999999],"typeId":"905c0666-7ddd-4192-a785-7e454e84ab15","componentVersion":1,"instanceId":"19abf22e-c985-43dc-b307-bec227e65f21","orientation":"down","circleData":[[767.5,755],[745,755],[722.5,755]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[899.0789229999999,885.6579214999999],"typeId":"905c0666-7ddd-4192-a785-7e454e84ab15","componentVersion":1,"instanceId":"18c68858-ce98-4365-aa62-ff9cecd47749","orientation":"down","circleData":[[917.5,755],[895,755],[872.5,755]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"Comment":{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"IR sensor pins:\n  GND - GND\n  VCC - 5V\n  OUT(right)=GPIO17, \n  OUT(left)=GPIO27\n\n Instead of connecting GND, VCC to each of IR sensors individually, \n connect only a single GND, VCC from RPi to breadboard then \n distribute from there to IR sensors which are also connected to breadboard","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"backgroundColor":{"version":2,"id":"backgroundColor","label":"Background Color","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"backgroundOpacity":{"version":2,"id":"backgroundOpacity","label":"Background Opacity","description":"","units":"","type":"decimal","value":"1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"textColor":{"version":2,"id":"textColor","label":"Text Color","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"fontSize":{"version":2,"id":"fontSize","label":"Font Size","description":"","units":"","type":"integer","value":"12","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"font":{"version":2,"id":"font","label":"Font","description":"","units":"","type":"string","value":"Arial","displayFormat":"input","showOnComp":false,"isVisibleToUser":true}},"position":[1247.3264341267043,683.0797772307837],"typeId":"9a5a4baa-44d4-4aa0-8d82-488487322b20","componentVersion":1,"instanceId":"9d530ea4-6449-4e29-a81e-6c2c23ffcdbe","orientation":"up","circleData":[],"cirkitStudioVersion":"1.3.3"}],"bounds":{"top":"194.26042","left":"583.00000","width":"891.03542","height":"841.32290","x":"583.00000","y":"194.26042"},"cachedBreadboardPrettyViewWires":["{\"color\":\"#9929bd\",\"startPinId\":\"pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_0_15\",\"endPinId\":\"pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_38\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_37073b3b-134f-45d6-97fb-5c4c86637137_0_15_0\",\"rawEndPinId\":\"pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_38\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"602.5000000000_395.0000000000\\\",\\\"602.5000000000_185.0000000000\\\",\\\"1007.5000000000_185.0000000000\\\",\\\"1007.5000000000_215.0000000000\\\"]}\"}","{\"color\":\"#9929bd\",\"startPinId\":\"pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_1_16\",\"endPinId\":\"pin-type-component_19abf22e-c985-43dc-b307-bec227e65f21_2\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_37073b3b-134f-45d6-97fb-5c4c86637137_1_16_4\",\"rawEndPinId\":\"pin-type-component_19abf22e-c985-43dc-b307-bec227e65f21_2\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"587.5000000000_560.0000000000\\\",\\\"587.5000000000_680.0000000000\\\",\\\"722.5000000000_680.0000000000\\\",\\\"722.5000000000_755.0000000000\\\"]}\"}","{\"color\":\"#9929bd\",\"startPinId\":\"pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_0_15\",\"endPinId\":\"pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_1_16\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_37073b3b-134f-45d6-97fb-5c4c86637137_0_15_2\",\"rawEndPinId\":\"pin-type-breadboard-sub-pin_37073b3b-134f-45d6-97fb-5c4c86637137_1_16_3\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"602.5000000000_425.0000000000\\\",\\\"602.5000000000_485.0000000000\\\",\\\"587.5000000000_485.0000000000\\\",\\\"587.5000000000_545.0000000000\\\"]}\"}","{\"color\":\"#9929bd\",\"startPinId\":\"pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_1_0\",\"endPinId\":\"pin-type-component_18c68858-ce98-4365-aa62-ff9cecd47749_2\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_37073b3b-134f-45d6-97fb-5c4c86637137_1_0_4\",\"rawEndPinId\":\"pin-type-component_18c68858-ce98-4365-aa62-ff9cecd47749_2\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"827.5000000000_560.0000000000\\\",\\\"872.5000000000_560.0000000000\\\",\\\"872.5000000000_755.0000000000\\\"]}\"}","{\"color\":\"#9929bd\",\"startPinId\":\"pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_1_0\",\"endPinId\":\"pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_0_15\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_37073b3b-134f-45d6-97fb-5c4c86637137_1_0_3\",\"rawEndPinId\":\"pin-type-breadboard-sub-pin_37073b3b-134f-45d6-97fb-5c4c86637137_0_15_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"827.5000000000_545.0000000000\\\",\\\"827.5000000000_410.0000000000\\\",\\\"602.5000000000_410.0000000000\\\"]}\"}","{\"color\":\"#000000\",\"startPinId\":\"pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_0_16\",\"endPinId\":\"pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_37\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_37073b3b-134f-45d6-97fb-5c4c86637137_0_16_0\",\"rawEndPinId\":\"pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_37\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"587.5000000000_395.0000000000\\\",\\\"587.5000000000_170.0000000000\\\",\\\"1022.5000000000_170.0000000000\\\",\\\"1022.5000000000_215.0000000000\\\"]}\"}","{\"color\":\"#000000\",\"startPinId\":\"pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_1_1\",\"endPinId\":\"pin-type-component_18c68858-ce98-4365-aa62-ff9cecd47749_1\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_37073b3b-134f-45d6-97fb-5c4c86637137_1_1_4\",\"rawEndPinId\":\"pin-type-component_18c68858-ce98-4365-aa62-ff9cecd47749_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"812.5000000000_560.0000000000\\\",\\\"812.5000000000_725.0000000000\\\",\\\"895.0000000000_725.0000000000\\\",\\\"895.0000000000_755.0000000000\\\"]}\"}","{\"color\":\"#000000\",\"startPinId\":\"pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_1_1\",\"endPinId\":\"pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_0_16\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_37073b3b-134f-45d6-97fb-5c4c86637137_1_1_3\",\"rawEndPinId\":\"pin-type-breadboard-sub-pin_37073b3b-134f-45d6-97fb-5c4c86637137_0_16_2\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"812.5000000000_545.0000000000\\\",\\\"812.5000000000_470.0000000000\\\",\\\"587.5000000000_470.0000000000\\\",\\\"587.5000000000_425.0000000000\\\"]}\"}","{\"color\":\"#000000\",\"startPinId\":\"pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_1_15\",\"endPinId\":\"pin-type-component_19abf22e-c985-43dc-b307-bec227e65f21_1\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_37073b3b-134f-45d6-97fb-5c4c86637137_1_15_4\",\"rawEndPinId\":\"pin-type-component_19abf22e-c985-43dc-b307-bec227e65f21_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"602.5000000000_560.0000000000\\\",\\\"602.5000000000_665.0000000000\\\",\\\"745.0000000000_665.0000000000\\\",\\\"745.0000000000_755.0000000000\\\"]}\"}","{\"color\":\"#000000\",\"startPinId\":\"pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_1_15\",\"endPinId\":\"pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_0_16\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_37073b3b-134f-45d6-97fb-5c4c86637137_1_15_3\",\"rawEndPinId\":\"pin-type-breadboard-sub-pin_37073b3b-134f-45d6-97fb-5c4c86637137_0_16_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"602.5000000000_545.0000000000\\\",\\\"550.0000000000_545.0000000000\\\",\\\"550.0000000000_410.0000000000\\\",\\\"587.5000000000_410.0000000000\\\"]}\"}","{\"color\":\"#ff9300\",\"startPinId\":\"pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_1_14\",\"endPinId\":\"pin-type-component_19abf22e-c985-43dc-b307-bec227e65f21_0\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_37073b3b-134f-45d6-97fb-5c4c86637137_1_14_4\",\"rawEndPinId\":\"pin-type-component_19abf22e-c985-43dc-b307-bec227e65f21_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"617.5000000000_560.0000000000\\\",\\\"617.5000000000_650.0000000000\\\",\\\"767.5000000000_650.0000000000\\\",\\\"767.5000000000_755.0000000000\\\"]}\"}","{\"color\":\"#ff9300\",\"startPinId\":\"pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_1_14\",\"endPinId\":\"pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_5\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_37073b3b-134f-45d6-97fb-5c4c86637137_1_14_3\",\"rawEndPinId\":\"pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_5\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"617.5000000000_545.0000000000\\\",\\\"617.5000000000_260.0000000000\\\",\\\"1067.5000000000_260.0000000000\\\",\\\"1067.5000000000_230.0000000000\\\"]}\"}","{\"color\":\"#e32400\",\"startPinId\":\"pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_1_2\",\"endPinId\":\"pin-type-component_18c68858-ce98-4365-aa62-ff9cecd47749_0\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_37073b3b-134f-45d6-97fb-5c4c86637137_1_2_4\",\"rawEndPinId\":\"pin-type-component_18c68858-ce98-4365-aa62-ff9cecd47749_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"797.5000000000_560.0000000000\\\",\\\"797.5000000000_702.5000000000\\\",\\\"917.5000000000_702.5000000000\\\",\\\"917.5000000000_755.0000000000\\\"]}\"}","{\"color\":\"#e32400\",\"startPinId\":\"pin-type-breadboard_37073b3b-134f-45d6-97fb-5c4c86637137_1_2\",\"endPinId\":\"pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_6\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_37073b3b-134f-45d6-97fb-5c4c86637137_1_2_3\",\"rawEndPinId\":\"pin-type-component_9ed9f913-4687-4140-b5ca-f53cf9998566_6\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"797.5000000000_545.0000000000\\\",\\\"797.5000000000_320.0000000000\\\",\\\"1082.5000000000_320.0000000000\\\",\\\"1082.5000000000_230.0000000000\\\"]}\"}"],"projectDescription":""}PK
     8p�[               jsons/PK
     8p�[��LQ  Q     jsons/user_defined.json{"type":"user_defined","version":"0.0.1","subtypes":[{"subtypeName":"Raspberry Pi 3B","category":["User Defined"],"userDefined":true,"id":"b739cbaf-bacb-4ee2-abf3-78459baee6db","subtypeDescription":"","subtypePic":"8a866263-8c14-4821-a3ed-cf7b88c4ff1b.png","pinInfo":{"numDisplayCols":"34.16220","numDisplayRows":"22.82490","pins":[{"uniquePinIdString":"0","positionMil":"329.37500,2110.89280","isAnchorPin":true,"label":"1"},{"uniquePinIdString":"1","positionMil":"429.37500,2110.89280","isAnchorPin":false,"label":"3"},{"uniquePinIdString":"2","positionMil":"529.37500,2110.89280","isAnchorPin":false,"label":"5"},{"uniquePinIdString":"3","positionMil":"629.37500,2110.89280","isAnchorPin":false,"label":"7"},{"uniquePinIdString":"4","positionMil":"729.37500,2110.89280","isAnchorPin":false,"label":"9"},{"uniquePinIdString":"5","positionMil":"829.37500,2110.89280","isAnchorPin":false,"label":"11"},{"uniquePinIdString":"6","positionMil":"929.37500,2110.89280","isAnchorPin":false,"label":"13"},{"uniquePinIdString":"7","positionMil":"1029.37500,2110.89280","isAnchorPin":false,"label":"15"},{"uniquePinIdString":"8","positionMil":"1129.37500,2110.89280","isAnchorPin":false,"label":"17"},{"uniquePinIdString":"10","positionMil":"1329.37500,2110.89280","isAnchorPin":false,"label":"21"},{"uniquePinIdString":"11","positionMil":"1429.37500,2110.89280","isAnchorPin":false,"label":"23"},{"uniquePinIdString":"12","positionMil":"1529.37500,2110.89280","isAnchorPin":false,"label":"25"},{"uniquePinIdString":"13","positionMil":"1629.37500,2110.89280","isAnchorPin":false,"label":"27"},{"uniquePinIdString":"14","positionMil":"1729.37500,2110.89280","isAnchorPin":false,"label":"29"},{"uniquePinIdString":"16","positionMil":"1929.37500,2110.89280","isAnchorPin":false,"label":"33"},{"uniquePinIdString":"18","positionMil":"2129.37500,2110.89280","isAnchorPin":false,"label":"37"},{"uniquePinIdString":"19","positionMil":"2229.37500,2110.89280","isAnchorPin":false,"label":"39"},{"uniquePinIdString":"20","positionMil":"2229.37500,2210.89280","isAnchorPin":false,"label":"40"},{"uniquePinIdString":"21","positionMil":"2129.37500,2210.89280","isAnchorPin":false,"label":"38"},{"uniquePinIdString":"22","positionMil":"2029.37500,2210.89280","isAnchorPin":false,"label":"36"},{"uniquePinIdString":"23","positionMil":"1929.37500,2210.89280","isAnchorPin":false,"label":"34"},{"uniquePinIdString":"24","positionMil":"1829.37500,2210.89280","isAnchorPin":false,"label":"32"},{"uniquePinIdString":"25","positionMil":"1729.37500,2210.89280","isAnchorPin":false,"label":"30"},{"uniquePinIdString":"27","positionMil":"1529.37500,2210.89280","isAnchorPin":false,"label":"26"},{"uniquePinIdString":"28","positionMil":"1429.37500,2210.89280","isAnchorPin":false,"label":"24"},{"uniquePinIdString":"29","positionMil":"1329.37500,2210.89280","isAnchorPin":false,"label":"22"},{"uniquePinIdString":"30","positionMil":"1229.37500,2210.89280","isAnchorPin":false,"label":"20"},{"uniquePinIdString":"31","positionMil":"1129.37500,2210.89280","isAnchorPin":false,"label":"18"},{"uniquePinIdString":"32","positionMil":"1029.37500,2210.89280","isAnchorPin":false,"label":"16"},{"uniquePinIdString":"33","positionMil":"929.37500,2210.89280","isAnchorPin":false,"label":"14"},{"uniquePinIdString":"34","positionMil":"829.37500,2210.89280","isAnchorPin":false,"label":"12"},{"uniquePinIdString":"35","positionMil":"729.37500,2210.89280","isAnchorPin":false,"label":"10"},{"uniquePinIdString":"36","positionMil":"629.37500,2210.89280","isAnchorPin":false,"label":"8"},{"uniquePinIdString":"37","positionMil":"529.37500,2210.89280","isAnchorPin":false,"label":"6"},{"uniquePinIdString":"38","positionMil":"429.37500,2210.89280","isAnchorPin":false,"label":"4"},{"uniquePinIdString":"39","positionMil":"329.37500,2210.89280","isAnchorPin":false,"label":"2(5V)"},{"uniquePinIdString":"40","positionMil":"1229.37500,2110.89280","isAnchorPin":false,"label":"19"},{"uniquePinIdString":"41","positionMil":"1629.37500,2210.89280","isAnchorPin":false,"label":"28"},{"uniquePinIdString":"15","positionMil":"1829.37500,2110.89280","isAnchorPin":false,"label":"31"},{"uniquePinIdString":"17","positionMil":"2029.37500,2110.89280","isAnchorPin":false,"label":"35"}],"pinType":"wired"},"properties":[{"type":"string","name":"mpn","value":"RPI3-MODB-16GB-NOOBS","unit":"","showOnComp":false,"userVisible":false,"required":true},{"type":"string","name":"manufacturer","value":"Raspberry Pi","unit":"","showOnComp":false,"userVisible":false,"required":true}],"iconPic":"b53b2c7c-bb6b-4047-8ddd-b279832d777a.png","componentVersion":1,"imageLocation":"local_cache","hasComponentImageSvg":false,"componentImageSvgUrl":""},{"subtypeName":"ir sensor ","category":["User Defined"],"id":"905c0666-7ddd-4192-a785-7e454e84ab15","componentVersion":1,"userDefined":true,"subtypeDescription":"","subtypePic":"8f771a2d-db90-4bfd-8b3e-8d66edcda07a.png","iconPic":"0c7fd013-2f4e-47d0-a46e-2d19cc1fd6f6.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"6.66667","numDisplayRows":"18.65672","pins":[{"uniquePinIdString":"0","positionMil":"210.52632,61.78319","isAnchorPin":true,"label":"out"},{"uniquePinIdString":"1","positionMil":"360.52632,61.78319","isAnchorPin":false,"label":"gnd"},{"uniquePinIdString":"2","positionMil":"510.52632,61.78319","isAnchorPin":false,"label":"vcc"}],"pinType":"wired"},"properties":[],"hasComponentImageSvg":false,"componentImageSvgUrl":""},{"subtypeName":"ir sensor ","category":["User Defined"],"id":"905c0666-7ddd-4192-a785-7e454e84ab15","componentVersion":1,"userDefined":true,"subtypeDescription":"","subtypePic":"8f771a2d-db90-4bfd-8b3e-8d66edcda07a.png","iconPic":"0c7fd013-2f4e-47d0-a46e-2d19cc1fd6f6.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"6.66667","numDisplayRows":"18.65672","pins":[{"uniquePinIdString":"0","positionMil":"210.52632,61.78319","isAnchorPin":true,"label":"out"},{"uniquePinIdString":"1","positionMil":"360.52632,61.78319","isAnchorPin":false,"label":"gnd"},{"uniquePinIdString":"2","positionMil":"510.52632,61.78319","isAnchorPin":false,"label":"vcc"}],"pinType":"wired"},"properties":[],"hasComponentImageSvg":false,"componentImageSvgUrl":""},{"subtypeName":"Comment V2","category":["User Defined"],"componentClass":"textbox","userDefined":true,"id":"9a5a4baa-44d4-4aa0-8d82-488487322b20","subtypeDescription":"","subtypePic":"c88b2895-5e8b-4a57-9f9a-b80dd50058b1.png","pinInfo":{"numPins":"0","polarity":[],"pinType":"movable"},"properties":[{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"text box (click to edit)","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"backgroundColor","label":"Background Color","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"backgroundOpacity","label":"Background Opacity","description":"","units":"","type":"decimal","value":"1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"textColor","label":"Text Color","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"fontSize","label":"Font Size","description":"","units":"","type":"integer","value":"10","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"font","label":"Font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true}],"iconPic":"d3694a2e-5bba-40c3-8069-8db85c4c9209.png","componentVersion":1,"imageLocation":"local_cache","propertiesV2":[],"hasComponentImageSvg":false,"componentImageSvgUrl":""}]}PK
     8p�[               images/PK
     8p�[����^� ^� /   images/8a866263-8c14-4821-a3ed-cf7b88c4ff1b.png�PNG

   IHDR  �  �   vEj�   	pHYs  �  ���R/   �eXIfII*            (           V       ^   1 
   f   i�    p       �     �     ezgif.com  �       �    �  �    �      �w��  �iTXtXML:com.adobe.xmp     <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="XMP Core 6.0.0">
   <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#">
      <rdf:Description rdf:about=""
            xmlns:tiff="http://ns.adobe.com/tiff/1.0/"
            xmlns:xmp="http://ns.adobe.com/xap/1.0/">
         <tiff:Orientation>1</tiff:Orientation>
         <xmp:CreatorTool>ezgif.com</xmp:CreatorTool>
      </rdf:Description>
   </rdf:RDF>
</x:xmpmeta>
�[n  ��IDATx���	|]gy�����w�ڭ}�-/��@B��B�Z��RJJ��a銁N�$$��t���@[�a�RJ
ek�eŉ�Œ-/�"˖Y�,k�s�׉IKbk��9�����J�%ٺ����<�'Q�z�T����g(K!�ُ���l	έ���                      ��	hI˺��{WԜ�Ҵ�'��mJ�:���gp=�b��L �E�(A��{5�V���˜'�|�v�s��ޞQ��d`��o�                       ���O�?+�m��v���lS7ކt�y{���#Z�Qe�$�2@l�êtv�έM�.����_��Q�ݩ?W�n                       ��fk��g3���=�y�иs�����񧝷���l�Դ DA1�d����Q������p7)�����ʻ�9��                       ���l�v�7�	�m��8��;�>���9�[�� �A1~���T�6;;�;;��5�lR�s�z LH                        �U��v�� ��p^�;�_!�@Yڭ���5#(�OL0L��ԲM�2�0Ζ@                        ��Rg�K!g3f��������?(K�کeX1�b��A�*�W8���l�tv�)7ҵ                        �!K&!�l��5�)=�o+�ojI_ӧ5! 7EP��<�$g��
g��Fgg��#U                       ���V��[��?��9����}UOhP ~A1^�SA��Ev�O;)rn                       �A���*`��k����_VH_�c:  A1n��p���|��ى                       �]�B�����7Bc�=���A1n�*Ի4��wޫ                        ı�1f{H�S@�ղ��'tU@�!(�v*��z�s�g��&g��                       �\�ἾCA}F;�E���Q=% NHK;T��ޭ��yo�                        p+9�����m�~����2�E�Ԭ #(&�g'�s�g�w                        �F�
9ی��C��J�'��N	�!BJ�'��u��sy�s�.                        \r����_�}�y������A1��S�����C��,                        DJ����l�j��NA}J��{|���Hy@I��;5��v�+                        �%�lwk����ۿ���mFPL��tv��S
�:��	                        �Ћ����}S��=��<���py6 fF���                         7y���fc���Փ<���pxX�׌>���                        7{��է����}ZGx A1���c
�.                       �+���6%�MzH�D��ь #(f->�\������^�i	)�IJw�e'�)˹���no'���1R�IJ^�;�;�-jqyɾyiN�PHˡe�.]�3o��hzqV3�Wu�y{i����В                 x��`��q75�ٶ�ݹ���)	I
8/���s�	JM��n����P@���`߿�4�n���U�vnyA�LM����g�׸/��W5��       DT�z�����ǔ�?�N-p!�bVc���������{E%U�����<��>��9��:ϵ'�	1��f�����]�����漽v��m�^ԅ��                �G0TAr֍�v��G�s� T3�4��uq�Θ��g��O_���W/����g�`U      ��Fg�]ֻ��ޯ��o\����ڡm�џ*�������BUg��n%�L+TAr����(=1�ni���&����s::{FG��v�I��Թk�                p���1u�j3K�׹���يRsb6��VR�Ub��<)���|1�dc�\�����gj�Ok����      �RH]
��ڡ�jI֧uQ�Ks+*M	�7�_wދM��G$�Ԙ�Q-���(��0�i��=Y�V��i�}fS���8{����I�|J��㚘;/                @�A;�5�Ru�<�DU�EJ	��5��엥���v�����Ҽ�͞���I�]��Хq;0u9�,      �R��P����W��+\�������в>����������2�fW�-�J���߻Tvb�:sk����5z��/�����I͇                ���d�f���Ը?�e&�)^�:�MY�vS���]]������>f�c����U     ��8ۗ�C����	1��7�a�hAײ~�y/(X����:u�5�#�J����3a:�74�͘_^���I�>�=����S
9/                ��1�N;r�m�{gN��Ӌ�p3&L�-��n�rhYG�L���#�s��_:��e��     <����;�CU�>��Z��g;�j-��P����"m�kҖ�Zu�T+1� �]r0��?���/ץ�Y{B}��1�������                ��JS�%��n]y�JKH����e����e/��Q/�k�������=+      ܐ�l�֌^����N	�2�b��^�(Isn}���6B�$�wmhЋ6�h[^��3���NJ�mv{�B�9���G��s��P               ��K{N�n/hUW^��R��1�Q�����W���)�]8��Oi�ҸB�      �J-iP��)}A@c|@-J�_:�6+%�-�Nw���JO$Q=����r��_�r�ݩ}��~�:%                �UE���SwmV~r��iv{���t��%}����{vPC3�
��     q-W!��v�u��_�검(������{���{¹��8ՒU����e���W�|O�L/�}�/�۳�1�>�O'��mGڔ>˾��hը�3��W�7��D�pk�2/i�jD~t^:F;���,�\(�@݀�R��W�g�Uz�T��sy�tx�a�U�R�:v(�nn)aI���i1qQ~U{�V���'�Nh�pB~�>����mb�ح�'��麧���o5iV�,E�+q���.�\�_���~�^���i�5\;,?�4�I)���R@�ҕ�+��bUNV
�v>�����W�ˉ�tp���[.k�~�'�˯�OW��\�pkE:QxB~�:���C�
���-$.h_�>���cMʾ�-�ڑ�G4���59Wr�x��sO+`�CuC�3�<�v-M��@ ���aͤ�ȯ��;��	֗+1�=�ъQ�Up9��C�J\��r�[����K�omC��
��+n�t�i/9. L8��m���S��w�O��K{�v�ڴ���0�1      ��J��zX��S�w�W�~M�Z��QH�SՐ������[�*g�M��ṡ1/��7N�ѷ���ܒ~�.�G6+�r��2��k_�>_6�L�}��"�ʘ�P�T=����Ƅ�t��V�<E�+�3ԣ=-{4�:+�)�,W�	|W*c"CII��J^LV�@�����������ݾl�3��&D
+�4ޤĥD_[�c�m��l!6n��mܮ��>_6�m:�ɆObe���`�/��6\�`����w%̾!�@��l~R~c֗]]J�F@�Jmڦ�M{5��f���e�8�}���sO���ߘ�s�)e� ���>�C��i.��|u��Tq�BX�5��~*6�ۻ����L��J�6p�v���b�A��:�?M@�J�i���&��T�s9G�#�vm�[{v}���/?��R�l��2[l��b��W�`BbL`5�˕1����d;��o��r����U��VK�/kLi��jae�P3(f�̿A�p���L�DA�^[����
Srn�Ƙa��8�����..�7�     �&jҿ�!���c��A1�f��2�8�LT�&���K�sj�DxWC�F5�߭wռJ�9;������e�s�=�t)�
�T�a�X�f��AM������B*�N�L�-��S3�Tkc�㻆���e�f����G!�ڔ�-����/�4gۨ�D��j�`?6�c��sŢ�zu�N����Ѳ���m;�M��:�a��zzl����b!]=���v�M�h�`R~q#���}%�o����/!]�ud��5�ӅL�4�An��)<_��P�j���g�̱P�b|^�\+��0����~ͦ����ҵ��������g���mUB�sO�a�{�;�˶�ZL�OX!�k���6�cɓ'����M֕�����>�)_���2�24k5lm��M�����F5�7�oX������� S�`֗&H+g������i�����ɿ�T�*'*��3�ъ����h娀H0��͹������f%X�{�h��կ�;�^�����3O�熵��5o     �HV@�j�^�DݯOjZ@�_��C�OK�������EzmI��,�Tf"��~���j/��md愾1ٯ�ݯ�K�B����|cm�֙�3�:�9��i�3�~��G!����-�[|3��Ę���	o,9WbS~h�c����h�k��l����Z���!1kUu��>_.�����+96�4`�RR�;Ыݭ�h�#�t��:��X�Ԙ(�~X�	!m9�"��9Oc&���x�������|#�����`�{�D�jN�E�D\�O3_�b�z	�Y+�.7A�{Z��b�{��fO��\�5�c�mÄ���ٷ��e�n�'z�Z2!���p���Ƌ��u����ٷ��hw�nϯ/m��VN��6j-n©�T���B�>~�C�����eo�^ͤ{����x���B�V&��<_�T����,��x�^S�Mũ�����l��d��s�O������S      V�Z�n=�7�	
���
����^��(���ڲ�tO����k��𿦬r�=P���ٽ�ʉ��5ưvR��)�n=ܪ��M�{���B��0��z�zl��WQH7&�7x���B���C3Ӝ��6�z���L�Ϳ�/��9�������^n�˙��惄Ĭ�	��>�]��vy:,�L͘%�t���5�f��'�U�ѻ�X��>���w�W��vk9��	�����9n�4�I�u����n3_��jUOT��f���T{^���	.mX�ޖ��I�n�	�+:Wĵ�u�C3!�ᑸ������ާ��9yն�mʺ�%�O͉��:VrL^Eix�ϥ{~}ij����c�����H���/©:U��	BH����:�/[���4Ay&��a�lmÁ�׃�3�[�@ix�N��ǔ	֣6�Dw���ś�`?JR���Uw��ʗ���ЗO|_��O
      N4*�j�ީ��agX?���q<�&�2��/-��[�nWuz���S���^������X3
�¯�h�-�8Y��#Ӝ�+�j����f�M棐*�Lv��N�h*�{�|R�������^��τ)���������6���f���q��6`���Ի�z��|��&�B~u'���x�qy��3�x�Q��3���f>BH��<߶��i�vؓ�|'T6Y&��������m��Ya��:}���mګ��/o����/7�B^&x�{����5�콠bBz��p0ǐ�'��}�p�ay!��e֗��oW_G���
*6!���e�B�!]�S�����1�����Bxd�f{v!��e��7�l���A8���W�B����Z`��
��pGA��g�����Ӯ�
�B     �Lg���g���)o]��k���AuiI_sn�ȇL0ȫ���-�/VAr� ���X+
�"��X���AO5�I�f�3�˄��6t�v���L3�-���#�i��P�mИ��NX�T�a��<�4��,<�̷et�m�Bx�f>�}��;�|E��z�U/s?0E�{��xf�;!��a���N�)i9I�7z���|�\�'��2k����e�.�4�Bf��z��6@M�{��τG�)��i���Ҟ�=򊌹gBH	�	+;�}d��5x������b3!��a���D�ͦz#,Ƭ/���~-]�ت<]i���+!������F������m��mv�Wӱ&{]�D�	y�9�d�?!��8ǜ���a}f�a��&�j*�;���FF��u�v��Ƨ�
CP�Bڲ*��z��^���N��7'��|�k     �52��ߧ5�Cz��w��Z���~P�QP_rne�g��m8�ݥە��,��<{2�Е	}�ط�����#:(��</5�1�9�R��ئ�����n
�lHӶ"¬�ڏ�kxiX��r;Ә�?M!U����4��\�Q�H'�:�f���.e�f
�Qx�P���h�+>_��#Ls��`'���k6���|��F^�D��f�2�7�BYII�>�݆������IMG���ɂ�r;,W8U��2B2�2�����>�7�e]ɲ�BH#���v�뉩�7�@��˹Bd�f��7멆��v�6��a����mh�L���LH�Y�ͧ	�Q1Ya�9�T������2�������|��,y)�^kM\�w�[,՝��ǒ^��8ި�g	!��}p����\_�@id���mcm�֙�3r;BH#+o&�s�p]I�D��x��V��'���aT�Q���߭�W�T_8�]���~-��     �c�Ւ~��.}R����W�w����g�ƴ����G��ߡ�D&2c��3J���{u`愾p�;�!�1xS��3H!U4�f>-K����4��H]HU��^WO棐*JBR˱��7Q���﶐j�B�H�B3�)�3����,S����&�ۧ9��1��W3����d>S��0���!����!wO~'�4:�c��t�4Z5*��;^��3Bd���7�B=�l�x�{��i�ax6D�9���f��+96���9��Cm��T�{�b!���K��o�#�4:�mޢ�M{5��ΰBH��t����ʭ!��l�|�;ח�6D�9��A8-G[T4U��2�L`���d�fhہm��;"��Z���s|��m �4:� ��o���@�^Zԡ{+^���<+U���_����G���|RK!ww      �A�����ޠG��"������>����HjB��.ݮ{�oWf"Ӳ�v�Y���z��.����KO]toA��Ls����<S4Q9Yi��G+���g����SH%���4��js��w��oCb(�����&%��4^�f>
�����|Ls�.sh��5��f>;�y�[i�X�F��'�-W�8Ӝ�ń������{5��f>�9G�Ʃ�v�|��ܦ�x��ϔ��l3__{����&��v��V%�����5�X�X�1�!����f���|�l'$&J�y��#�^�d��܆��rs3_��2B��0����lվ�}��鮠bs�<�%/$�a���C����B]&x�\��o��l����Mm�	�'�4z� s�>V6&�!�4�� T��A8��FYHj:�d�%O���B]YW�욾�ٽ�p��������W�,5_�Z���}�w�m�/�O|��     �g����a��>��Xum�T�f���=�`�޸q��)�C�I�¥5�R���s�{qL~������<
�bg�ٍ�He�jDn�r�E������$�����ݮ��G!U���Qh9��%��]��y�B�h��|�=v���f>3͹�H�]���m�Mõ�:�wFn`B*z�z�z-U�.�̷ux��lqOXLթ*�L��e��l�SOi:kZn�4��)�*Qp1���!�E��fO���6��׽�[����MqG3!��a�!�OV+a1A���NHLl���������*�($�k�!s��nCH��6Gi������ذA�#���~�.�#,���)�P���N=���������e�̰�=-{4���e�\�m�7�=昽�t�]_�V�g���0nn��3����m���c�|�x�{�B����@�v7�a1�'��6����*O+.ũ�60�'7ަύKߛ     �e*����O����*k>�]��Ћ���􋵯Ui*�9[r봹�V�?7������3D���m�F�X*�*��kc�B��2�1{�z��uO�'�QH[�ز�d����t�,��|���ʘ��*VL��[��L�w�f!6̾��p��4��f>;�y�G��Ls����l�c��V}�Z��Bl��ͣ��O~ϊm3!��Wt�H	c	�_�?�?��+:Wd��}��o��|��Ɩ9������o���o��2�E9�s��pS3_��"�ib��X����4^�f>c� !���7�/[b��W5Q��S��Ɗ9n0׉�5�;ӟń�vt��g����<N�ds샊��4��!��bY�u"s_�I����bkL)!11�q�A8ձ�c�5�^�b�M�pL�KǡBHc��D��7+9ӟÆ�:ǐi�!�����m�6�j��A8����R���ujϮ)��������	���o8o�3|      LL��!U�q}D�*����#�ӂ������I�j^����`S��Գ�Q_>�}}���4r��D���|��7(�P���v���g $��KAmܦ����5�QH�f2��=������3��=l3��v[P�f��g6��x�{MG�����'b���4����6�
�e�-mXL'�՟�W�$Ӝc�6�n�`���rb��g{Ms)�:��1߆=��T�~��ȟΧ�/����G�{l<�L3_U��LxQ��L!�l3�3a��j�+>_l�{5�kZ�xIl+L��i�KYHb+}.]���}c��gHM)bˬ/���4\;�3ygb�3B��W��ux��l�]X!��Xh���mګ��ج/��di��V֗.Pz�T	K	����`�!e]�b��ў�=�K����`CH�Bk���d��7�j!��r-�FP1a1��!9K�U�L�)ު`�냈��r=���֙}��#���     �+}X;�׏9o��~P��U���sk�<.+1M�U�Lo(���9b"%�t�N�6��c�Կ�yZ�PH��9�O��u�v��Ƨ������.�N~�o�ו�+Q��R��)�2a1fj�Het��(�r���g���wk>1��|&A�=����E����i΄ĸ�	�1Ŗ}m}Q/�4�Q&D
�`���i�nXgr����4g�ɝɍ��wBH�%��|���O�T�m����7vQL��	!�;��&����/��|&��a��}�K��C��:�Ƌv3���߭�EBb�sl���:���nPqÉ�M�	�`��GZ�����~oBH�'{6[]�]�Ӷ'�߻�`��/B�f��	j�׸O2/D�{S��>E�<�@}��B�.f}i���[�5��A8����9��<]i��c���cC�{�<�,�C�|�z�_#�� DNb Aw����/Wz"�u}�9�΢N�8�E_9���     ?��v([Y���ܸ%o�<�
�M疧�ۛPs�˕�HC.b� 9[7�Y�*ڢ�>�w�=+��	��߅�f���G!�;�b�m�io�^ͤG���B*�*=[j�T���c��{�f���6�1�ٽl3�r�o�N3�i3M!fwI�O��^&H*Za1&X�p��F���|�[�P����i�˘Ͱǭ���b&�wu���/j��4m�^���F3_�>]ȊN3_�t�����)<_���v�E��τ��}Qڵ4�]̔�h7�B�^&��K��E��/y)ٮaY_��	�����f���z��%$�uBR��&{,y��dT�%!��9���!g�м��E�!�D�ۘkU�F6i_���̉��2&_��	�q!���|p��jx**�Ϭ/���~�R�yvΞ�=�M����?��H�ܧb�A8U���l�vw1�3�bW�.�b|d��&���u*M�k�	�v(��;�G����     �#�ь��S?�l�d�My�
��~&$�NV�^�4�Q�Y�fSN��p�/�'�M����yN�2SP�4gw3�|�Ѳ��?���4�d\���6���d>
�ܯd��T�F���i���f���u�8���*&��ϲt�<�a1f��9n0žp�ԅԨM�k;�f��9lp)��w�IZ�&
#�4g�3���n���E����@�2�B�V����&�|3!��Wp�@���z���~��t�Af�0�)��|U��T3Q#��9'h�bl3_ed��L����NH�{��Q�@�#�O����2���Y_�Xñ{>r�x<�߇R�K��n}���"T�et�rfrw2�&�g�nPS�S�^�7��P;�/],�RnT�����64�d����ro�^ͤEvN��r[� �*�*��k#�}X_�_�bҍ��ɑ]_"�r�2����΢Nn�1m�>�v��75h��N/\     �Oܫ%�ݧ��/��WJT����s˳#�	zsًt�˔�����W�)�C/.h���[�>"x�)�"$���dEt2�-�`��ܘ�����RyG��u�uh���|}�9{G4���~���n渮r��[�V�F�{�i�[��*!DH��Ec2���<�4g/hoRR(I�E�i�c��w��x���B�H5�uw��N��]_�f��AM�E��τ�6�7�7��f>s|j֗�Lsv�h4�U��V��j��Jϖ��U"��S�Sm�!��gB��8���]k�k9ܢ��E
XS�]͉�o8Vr,"_�R�0��IEj}�5ܥ�YBH�Μ�nk�p��䝉��0��G[��� B:Э�BH���ު���t�tD�G�D�jNB�f�@{�=b�p���k���#�n�w�;ԫ=�{4�٠bD�mzo����.���}uKn�����7&�
�     ��(K�ک�9[d'
ó�w��C*ג�)�ĴfW��oTez� �(K��'�ΞD�ӣ����k�7�B�#Ry����s �a1���43��;�d���L棐�{�/�G���i[�c��)������|�Y�SLs���g7�f����N~ϸ�4g���d>Bb���x���o�c�����ys��B:ح�9BH��<nۏ�k�y	w3!��c��Lד-a^_.%�I�IKI�7���-�[��i�f2»��?^��3��zI�T�		w3_�|�%2�3�	K	�ZB[؛�:v(�R>�<�C�Я��.?֯�3���	��ԅT��jw��wu����oh=ܪ��M�O��k�/V�f�;� ��k�km!��c���s����©>U��j�;� ���N=��tX�.!��\
j��6���Gl¯85W﫿[�r9���LL��ۗvء�'��	     �ެ��s���:[d���Ӽ�������?9�<�՜���wU�J�/��d&����K�y�o��V}
�F!�w���ۆn�S;���G!�wݘ�W7�3��i�3ET��
�c���C!�w���p7�iQ�9�9{Q�T�m����c��w�c���iߣ�Ĺ�|�m�۔5�%xˍf��.O3Ӝ����6�/�wi1��f>c֗��R�	)��|��zW�l�=n0���`BHͤwBb��N~��f���Fj	�1�|c�_�?,_/c.î)��s��k�K{Z����φ�^"��k���r�Ҟs���4!��:��� s��I�j���B�C�]#�ԋ��6�cɓ'�����c�x�2AO�C��ݾ[�a�O5!���C.��\W�<ة��M�gNÉ�Mzv�`\˛�km�]_1���r�K�����~Ep/s�����ʗ+5�CxӦ����_��:�/��S?T�\     ��ӌ�[����+�P�s���V�<�1�Lnz����x]aJ�>�v���������4��i���g6��x��])�Rl�-�ZGXӜ���d���7�QH�}&,�6i��Y��1��=�=4�xX8�����}�
�>�n�o�#�r�:G:)��0d���[�5���f>S��y5S�&��w��珕���kB�}II�>�݆�����4��&�����L3_�b�N�X��!���LP��i޽���6�t���������r�EESE�/=,�b~X����d����z�9o�=�m�3i�*�2�E939�w� �x�Y��!������;�k��^'`�1�X�Rok8֠�bP�K���딟-W�x��]���~g}ٶ�چgBH�ynxTHj;�f�L�o}ij�L����v֗-�[_�@�m��2�3�ý�{5��A8���L�h|���x�	:zO�k՛ߤGG��s�.	     ��ީ�4���~�፫��U��Oέ-�Ӕ�ƍ����W)1@�4��΢N5dn�'G�����B��(�,W�	
�� u!U��{mA�Z�����#��O棐�?2�2�=ح���55�1��?LsƦ����n�.�-,�i��Qp�@���z���5�}s?0�A��x߳���:��Ls��R��t��*&+lc�Z�����&,�6���|���lH��n�,�u'���Z��!��}p�������g�mH�2�?</�|�:�?M��f�u���\���̈́��@`9�-�[��i�f2����5ܥ�YBH��t�Ԯk���	!�s�����iߣ�Ĺ��}�~�3أ��d���N�)i9I�7^�߯:U�����L��m�iW�.-W_�@��s��G�5�4�ɂ�5}s�P|����dϮo�K���pl�SOi:kZp����w+;�k���9���-������3�_      ����C��>*���yPi
��έnyLQJ�>��S�ȩ�W���������_���B��1U}�Z�'��0a/�agW��&�SH�Of2��������QH�?&�e-�|�L��shӚ��LQ]��\�?�f����W0]���v�?L�	�Y�d>c� ����(9[b�/TX��c����f���1d{ߪ������3У�E��N�ʘ���6��B�YBb��<�Ǹ	�Z���Y�nڪ���b=�|6�t�R?1a1��r_kߪ�^�L������#��od��5�Ӆ����P���?
��}�]u��{���GB�f}i�!���k6e�A�f}i�\,2��O*&*�s�X�ت�^��jUOT�a��{���z!�>�Z���k�>�r�E��m��ɹ��ΑN�!}�/l�|}}���A8��`��U�J���W�_e&��ךߪ�3���c_�ե��      p���C����� �?(&����y{�<掂6���ne&�X�K$�ʗ�=�J����]�$�F�ZUNT
�c�%{��ڂ���[_�����jN���c%�V��R��m��^l��f>�m��)�k;ܦUV���u�K�W���G���B�7�����4�#-���v2���luRR	*9Wb��+k�c������4��Rs�IH�?����R�J]HU�@�v�����4�o&�ԗ���G����j��LXP��v��|��lҾ�}��s�f>B�/Ӯq�܏
.�s�SO7>���'�Կ�uHT��e�fSW���!1K����y�8]a�9�V����ԟ�W�d��?�nח�5�x��BH���X�*/Z� BH�k��p6\ڠ�C�/}��N7�n�`���rV7�ӘY�7�Ee�����E�jˮ�#��WC�V7�     �UzD��煸����z�y�3��@�~��.��x��x�9�V����_G���W7)
�W�^�g(��3���;ԫ=�{4���ŖR��)��>Y���.���w
��/u~e�|Ls�?�oXi3Ӝ�/�J�����7o�+�*V�f���d��������̱f�@����*���f>�9��J��̱�i'�ԿV��G���� Ӱ��m�Mח�����g�'�O���!�?s��w���A�E��z�U�/��wh��5����|�ܔY_�@{�W�L��}��ɛ~^�D�jNB�g��]_�m٫����<������_�nT`9��ꑛ~^�x��\�W�R��lW_{���^��!�5�kZ�x��~��g�8k$u����l�d�l�OvΡ6��L�!��\�"���UJ����R���G:ީ?=�O��S�.      �2�X�L�׷����
���n��CR����l~���j@��NJ�i�_y�;���u�\����ͶɗF�.�mp�N~��*~�#���J[P�B�|R���7�]�Z����i���f�|v��`�����qAρ�n���a1Ls�����`���w2_�R�-�M\t�i"�ϭ��N4�l�L�?���=�m���̗>�n������l3��|1R���|;��ɢ� i1I���B�'������BGHL|�;Qg�/��g�G2f	!����g���b����!���6�i�vXg�~��φ�:���yBH�A��lmv֗-Ͽ�$�4~����T�S�Κ��?7�Q&Ԛ��Pz��>�>`�©Bj‹Vս�[�m��;���a�!�N�)i)I�˞Ζ�-ʹ�#�_�����eˑ��̾��p��4�aB����d}��'����Ub A�}���������y     xP���>���q˝@;�Z���M95���{��DA,u_��T��Q�����8'D��8^t�H� �3��N~�Rs���_��q
���5�m�b��?��nT=���i���������ү�붡�l��s���NW��$Ӝ�JHv2�iИ��QXL�b����Wďj�k<ި�g��O̔�-�[��i�f2~�1�L)!1q�t��>��f>Bz��xb���z��}���nBH;uBG^�����d�b칧��Z���Ϝ�lo`�G�C3_������i7�Lď��l{�`�K?!��ǜ�6�����Bօ���!�\ě��jk�����v�M��	��'��6�i٣����B�*NW�cɱ������.e�f
���ܮ]m�q!�q($5i����B�b"ic��v�Ϩ:�X ��t�.�T��+�Ϟ     ��kI��u�>�3B\r_��U���$Ot(�`�7����5�VB���z74��7��>1�W::��L$ܘ�L�L�1Ŕ�l��潚I���*��f>3���z3�T��4unڮ��>��G!U���̷���_o��V�B�R���(�4a1f�����c��G�5�4�ɂI��i�9/1�9�f>ۤѶǾ�4��e'��l��̗u%˾��2>��f>BH�Y_�����M�%�4�=�����f����0R��W~�\���B|j:�d�%O���0=�=J\��%~��	*�a1ͻM�!�q̬#;v���TΔ2�f�뙄�ħ�����SO��m�4!���ww���'5�6Ci3�s��4�F*��1�(���O���c��q$�S�x��BI/¯'�Qjz�29�<WEZ�>��}��W�o�     �A�
��S/u�Y!R�*Ѳ����Dgszb�nx�^��" ϯ,5_Ot�[��k}ojPST�{)W�_����V�m�a R�73}�m�M��(��4��f��q��!�UNT*�T�b%-$	�+e>�[��=���Ls�k!�e�E�K��:Ue���2�2m!���*�. $&��f�M7]__��#$&Ιf>���<��̫�8U���߇�t���jN����f>s�(�P`�B������^;�b�B�o��}�|��6�"~��&�|&s��x����h�QU��f}�L=����x2�2!��,�Ж�-:Vv��%Tz��ֻ�pbBH�۳�pN����j��(����Bx�c�wT�\?]�;��3� ����������}�Y҆     �1ݺ��:o��{��P���E�'FK�'g����.�T n.-!E��t��"�_���o�AHS\Y}� \W8](�0�[����`��)U���f��)ְ�m�1����0�Z	�aח�4��:���Y�x��4�K\g���H\LT�$!����t���Sv��I��f��i@��;U���	�a=������(:_����Sv���
\?�<SAPL�$�������v�9����⥪I/�'G��k�     �ޮ�էO��B\qO�V�s^�DP�QlCb
S�v��)���e*N����[-��               `����Ѷ��-�R V�E�-�d�;���ԅ��     �Ճګ'�!n�#(�a�ݹ�W�-�^���6�'��꽲x�Y��_���9               X��i��U��/ �לU�'6�[�=�y�Ϟ     ��$*�/�C��#:!ą��<�MZ�g�뽶x�~��J`�6��걎_�o}^g�]               ��k˪�G[߮�tX���<=�����/h��     xH���e�W/�gtM���|DyZ�W���J��w׼Zo.{� �GUF�>��n}t�/t��)               X�;�:�`�O*1�  뗙����v��8�����}     �^%�q���۠�y�����A{���E� �6$g�ю��ǆ�J{/�	               ���Uڣ_�}��� �OR0Ql�)�&g�'�M      ��zH������k��١��o���d��4�U��
@d�&$����w|I�~��                ��{����W�R "�0=P��&e��g     xF@����1��b��ן�����h�G���Y����6}r�+��Ԡ                ���*_f7 �gB��b     ���*���z���%�������3��s+K.�����-o���Z���@�~�����ϓ{               �@ �j^�7m�M �ǄŤ'��ƾ���     �zݡJ}ع���/E?(fF�p^o�Ke&��m��%�B �+���Tz0E3�C               ���ؾ��n��x� D�]�=6,汃�OK�e     x�������EӾE7(惺C��k�2!1���N�g�
@l�i�}�M[�ۉ]               �U�y���&�Y�) ���g���~�ֺ     �\���>�-zD3��D/(�C�Ғ>��J������^Bb 0a1�T�:-,/���               ⍩��պ��\�,���ġ�V(DX     p�:-���/	����E����%�����Ԟ���K���{�ߠ����׳�               ēwU�R�/� �xU�]]��?�{     x�/�a}Y�ҷ߈NP��ڮ�;S�	�͖��3�F �%���7kni^?<?"                �l՝zK���>o,����9}��U     ��
鏴S��6'�B�bv*Y3�3�V�\ƄP|��ԓ�( �t=������T߅��w%%%(3=:�d�0���W����JVB0 ��8}�9�E$��$*=�u��?�ڵ%��-
�����v��ny9��y!��R����}��좮-,	���ٻ��������Y4�mɖ,۲%y���ر�A�
Jp����H�r�5���+p�
d����@[�VRL�=�eK^d���K�e�w�Q&�JB4�<#�z͜$h�F����|���S~n���7�9��1�ɖ���P�_�u��sv�gS]0���)b1��?��D5:��2�r���e�����HDQ�߲)/
(+��kO�Ȭ3��2��r������3��!g߀�
��1f*�/g��eTH���t�.�0q�)�Re|96>��Y��g��|V��)|�)fg���8��d��
)-h���1�'f`&U��m�����$�_&[^n�l��`Ɨã��5$U��/'����4מ���p˟�8S�c�`�w�<O�s3�A��     �\���)g�)aQH��ڣ�+�y�,�s�n��3��d� ���b�j�;�W���#�-BjZ�$[�R��I�c�jn�ؤ�dg���వ�͒���^��I�̟I��U�*�KS�⹖�Ój���̤;��5�v�o4�ɦ>�����I�u�
��2��<Nݽ�j�V��S�E�L��{�j����o銝���Zz5<&$���kr|B᰽�s�0�p�d��ڶq�fg�e�A���VS۠F'�$�{F�����e��}CCK��&��$�(���di��~{C�#Sja|����Q_��҂v�̐����9��$�XU�#�
[|���Sg'�K7���"~��o�J߹����44*$���+559��Ǘ�]#��6�!����u�ie�LMă�6���U�3���]k���������MLJ���N��e9Z�2W���F�"jn�8s���=k��?h���\ih�u�>�|�f2UU,QV��9N��^0�'��9�?Iv�Yk��7h�M�f��e�3�f|��.[�K��D ����hbnZ?�|R      V��ݤ�z^Hy�]��q�w�o��>��B�n�6H�@H�6�[7�K��}Bjڽ�BO<�`��(�����w{Y,
��li���h�nBU<��'��މ��Og��#��+�f�ߟ����XU�D��4uv�*�l��B$&�w��bb~�{wU��ǎ)la,��o�9w`e�[6o\�õ�233USk��~��a�Qz(����g땑n߂���!�=1��ې�H��O[�'�mTlξ�S��w8g��ܐ�VYi���6[�1:�#���=g�գO�+-h�ߟ����c�;���+;+]�-=
�:���Ęq/�K7��>���Z�y��3���`��kllL1�!]Q]Y���>��Y���/�s��n�ڳ�R�=y��XLG��"�ξAp�i�����+c1&���'?�W���5�kt����XLSۀb1���,V{w�ӣO�[�1����Aq��eKrT�����+�6�H����p��1��ǜ�eȾ������X�fi<��3`],&U�&�/S���j]E$H)׬�Tӣz��V      ʧ��
���ćL).����Ƿ�G�,sq���l� ���`��zӕ���]�RS<��I)f�-'&g��=��}���⥹2���׷Y3�*�i�%�2�߯��\�G?�P��14<��As�a�E��ķ6�b��)s�-"1�2v��c_,�DbF���o��fb15�Q���[���܉���W�`Ls�:�&+3�3v��.c��9==);W��a_,f22������r֞a�WT��MW�pm�U��ZM�7����r��u��bFF#�5Q{ޞ���e��M��<��p�&��o8wo�u��ށq����SHw�X�Q�q`��XL�N�-��˨=��E/==��<���7�s����TdBp�|,�Y�){��SSsj�싏/�\�vM^^��o�/��6���q���b��M��H�Kw-/ɋom���#1�Db�_��C�w�v�3&342�����X�9g��7hM,Ɯ7�l�V0S��eʪ�)�_T_!��?j ����[�/�-5��m     ��N�*]�l�,���bnҕ���΂J]��M��J���w듇����R�����'����[&���O$�#��r��2kb1�-}���H��XL�5���b"�Gl���/��q�����m���q���̖�e��m�"�ĘǜCz"�y��z+��#1Db<2�iPln���HL�K��X�捫���4��H�7l�ŘHLO���bS,&���Db��z�,�;kO�~��2Bޏ/M$fd�H�W�W���q;b1�����">���b�<�ʚX���LN���i�VY�1����^�=y��b�lZ��#�V�/���xj~|yB>''�%�b1�HL�����9�b�Ɨި^W����GbZz`|���cÁ� ���?M���n�p��     ��b��>���U������F���oe�ՙ�t��+���4sǄ[��Ч뾯h���8���ٵ��X��Č:���x͖XL��İ��S�X�Ï�P������I���X<����ϳX��>U��">��X�Y�_X�����?F$�6�b^��;琞2���-�Ŵu)2=I$�c�vTx�!c[b1&���S�-�����z�Y��5��9��s7e�b1&s����ǂ΁��3���c�=���N�������i�\����^_���K&���J=��	�=����=�����X̳�5�n�?5=���>�=y�� ˊXLs� ���]�/�+���=61���A�=y��b�9\cs����fLA$��X�o����X���$���1���fs��=���@X�6�[�lH]�i����?�M����      ,����9۫����PL�nu�W�"E����+����]�����tW�/���e,&��!c��XL���hW(��	U&Ý���O�}��c��}+��'c���K�[/b1�HLS��,L��y�1���1"1���b��il��X�܋��� �9m��~�'����a"1���4*6���)���H�=�c1�:\���b��V"1��:���2��DyiA|�E,&�����E|�0����x�����(�Kl�Z����$c�/�c|i��p�v��],��H�Uvl�.1���~"1��:��6��hD�����9��
z0��Db:{��
�+��[/b1f|�����&s������KKx�17�;��痩.��mxg��� R�ʌ%�?ߥ[[3Q�     K��!}\w�zVHI��E������@(�Y��' ���{�95��v>%��x,����[�?19�&RY�xYn|�v,���_Db�b&^�����X��Ȕ����ƋX̋�?��x������l��~,�H�����=�Ŵu�H����ڱFO>۠؜{��im'c����x,�H]���˦��bDbl�R,�Ғ����F�#�/
,�b,���9�s��">;�X��{���cǔ�b,�pB�Db�����܋Ř;��$c�b1�=#�$c�c1�S�M}���Us<þ�&/�bL�Խ�xs�����p��;k�����Ϗ���ɋXL||��+�K���y��H����Db��c�"^�b⑘&�琩��ʷh{~� ,�sW��uo���H      ��+��s�gk~9R��O����S�,a��Y%��\]q��'zT3�$��=�+]��LEf��5�">K��i�GbX�g��b1G]�x;2Qo������f,f>�K$�Rn�bz�ǉ�X��XL<����\�������^�g6(��ݝ;�G4==I$�R�vT�����Sk'�[�X̦+]�ŘHL�E|V���T��1���^"1���b�1���$=cF���H����9{���c�v!3�!c����b�#1�,�T<s�:=�L�2\��v��jbr�kO�r3�Ĵ�)�b�/�|,f�j����Us����_�ʌ/qƗA>G���Qg7sleb1�XLM-]��b[��sƗ6��b�V�7f|��q�H���g���?��X�U64��(�ې��Z�G�/�& ��뜿���N�s�c     ��O{�q]�/�B�Y�i&�p�Q�U�|�^��d� ,N�_Y�v]w�N�GF��eb1�>Y��N�7�e22���~&RY��b����Ov(-��I4�}��`�x,fO�~��q�Cɛ@c"1=}�Db,gb1f�eW<�����K�&Y���b��]�7�H�b�ށq����P�r&s�H�Ɠ��5���^��X-''����ك�I�Ř;�Oq�w�X��4H���bL$����7pi5�b1�Db����<�x��^H�1}t,��>"1�+_Y�&3��4����Ŝ�B,�Db�F�����b�E522��XL<��C$�r!�ޙ�X�|$f�kO�s#c"1Mm�Db,WX��J,��cXss�ng�Ǘǝ�D��&����ە��#ٱ��an��ⱘ�܆��b�Ĥ�����Z�����8����H�"�1�\�_}� ,^X}�N�upCT     `�/j�~�<X(�bv�IT_�d��P����}�_/ �[A([�Z�}�з4c�}*ۻk]�b1����*��ŷɊ�4��HLj��PU��;��$�bF�"��'�*֮Y�&#c&R�$�2�BA缡2i����q���I[7�&-c"1�&�"������B,�))�;L$f�k��b��
=�L�bI��D"DbR���l\�R�G��i"�2L,�3�%-36Qw� מR�����ͩ���ǗfyNc3��T��X�Y�g"1�/S���:\מ�X����7�@��RA"��3�ξa���}cDbR�|,�I�ӑ�33���p�)%$;��9���)!5�1s��WZ�DbR�K����HM$���!�I�܆��)"1)��b�)9������Y
���}��,qC��ܩ�in�
     ��R#�J&���p���t��K�X����f.�X�6�ԇ�\�;~.�6s���'Z���u�0�*ŘXL��؂�+�)��_,��1���ێ����-���9ŘX�Y��Г���'YėbL,f�����nx����XǾ!��X��#-
�vR���/wzO-&�bE��#�����S��];+t��y��oGO����([EK�KB�enn��)��b�o]������&D�4��Y�T��S��baǗ�3�~��e*1����R.���o�e|�bL,���vu��I1&���X�c��O0�L9;��VMm�s�_�}������bb1˖�k.	�˩�)�)Č/w�f��:�{�t�^H1&38<�'vn�ܜ9$�J�܆�ե��X��}���HL�1��������?0����e�3q�Omx�
C9���o�������D9�     ��V}Rw�sR�B�b|�קe�40^Y�K��SǛW�V�x��~^               �M���D�rW	��c}�J}d����ɟ
     �BK�u��o���0����6�y�,quť��)�S�ukߨ��5�w               ��닷����S��ۯmՃ=     `��>��Н������C1W( ���{�6�Ғ�pjJ������wj::#               �K�Å���p�~�tt�M��     �L�f�1g�OH	�>S�w9�e���\}��28��g.Շ�\��N�L               �W>�n�~�2�p�
B���+t���4�     �Ub����m��z뽺P�
8��[�9_��|�r���7���g����1               ^����j}N� �2{��]~�����      ,���nr��
�{u���z��Nx[�^mϯ >�O7V�EW=w�g�               �iS�*���l@�;W���:8�(      �\�[�}VÂ�^](Ƨe������U� ~[^Z�n�z�>U�]�b1               n�
��ɪ���� 	>��ξ���n���      ,��Y}��~A�ڟ��Q�:ϻ䱐/�H� �kG�:]�|�~��                7\��*� ~גP�>��2���     �27h���<�k���>.�o�Z��L ��|`�zz�:&               $��K6�K�
 ���0����     �"e�۝�����B1�T���y�*�To^�K ��	��t㺷蓇�Q,               �Y���Zs� ���f���P��f'     `�>�<�y�0�RZ(fVw~�~y(���c�.���� El�[���F��~N               @2|��b��
 ����l}h�E�҉     �E��f����W��^y(�z-�OW�co/;[k�� ^.���3C�ꏌ               XH[���ol /��g����C'     `��;B1�z塘4��y�C�E���
 ^��@XW��Ds�               Jȟ�ֽY>�O �r�}���]����MSs�     �BL�Z��+�z�����R=�s�n�|�B�W����K6iO�=�_'               `!\Y�Z��( �R%��{�y���~     X§���l��`�WV[�Y�)���%�wjs�*���ڊ7���M�E               �k�J���=�?�ه��=���]     ���a�?��f���PLT�O��f��� ^���\�s�9���               ��U�*�� �Tfrͺ7��Cw+�	     �˕�K��	Vy���[U�i�U���󔛖) x�./ݣ���S�T�               �?��K6iK�j���)�\gm��}G     `�>$B1�y���]�<�呕K���g B����\����G               �T��W_$ X(^s��8�HtF      �D��\�U�`������Ї+.�� `��-ڨ���깡�               ^�����8�/ X(K�����=�~�o     `��f�g�ׂ5^^(�fmUL����tzA� `�}d�%���횋E               ��l]Qz� `��s�9�U��F�     �9��%B1Vyy����!�|~}pՅ�dX��L����;����?�����y������RC,��䴢��ߘBi!M�L�c`h")��¼l
�cffN��Yg�����/�@ �����!yF���o��������:��#���1��}3�a����L)�cMO/��!;+C�SB��O�q"?7[ݑ	gl!�3����8�z�?�����ch(Iמ�s��N��:fg�455������
�4;7#����7��1�?�LLN;��3�iaǗ��i����e��e*�t�I_fgjrr\HC�S����������1I0S�9V�sɅ���tdJH���I�ې��~��dn.��g�נR,SZ0M3��/S���d�ƗY�ؕ�e*�L�*b�=-��5ם���3�dn�->��Be� -ݟ�����ϟ�g     X`�n�V}^�+��P�t�<ri��� $��,�~�sP�sD#���?�ёq-_��������;�Ť 3����v/�J��/��С#M�fBUJhm�?6��}�������c1_*0����:T�,9����t�kQtnV�߉�=��('k��%K�u�h��GG��HLsK���$���d�t����|)�p]����D̅����(Sj[59I,&��k�$i�ˌp��Z;�!J�m~|��N�¼��5kf��J���k��]�$m|y�ɯΞ^�~ѹ�j�v����!��7�8��9Ɨ)���O!���%g|Yw¯�!Bũ`*2����X���eXG�[_���c]��	ɗZ��]�4Kk�4>>&�oxxB]]�Z^������[:D,&5�i���|�%�:Xע��I�~]�#�D��6�L���-��\{:��K�&��S~�3��m&�"�Z�
Ē�o�_����`?sC��':U�,9琹�!9�B,�k�Jt~�6@���l����q��     ��bz��L(�<s�v:ϕ�@��;V�- H���,]�|�~�����Q8��6�^���|RK��������� /���0��V���E3�,�Yk��f"�
�I{���e�����Y"�����0�d�kce��7k�	UV3��P0������ח��Q��\"�������
3U��:N,�z&�����D �����:X۪	��n��"1��@�^��$W1竹��X���B��#���2y�fQ�vg|y��E���`/���PZZ�ƗkW/�-b1V3���um�O��2;3�-��Us��X��L$Ƨ9���_n�,Q퉨����L$���[�9�_����u��S�s&ɵ'��HLfدd}��w��e�bR���tv*3#-i�aƗ���L,�v���e~�f��mC�iRd���L$flt\�P�=U�*t�1�w���'wnCf8M[̵��&��2�������f$s|�\u'D,�r&s�DG�F5ɒ��ƪr���ܕ�ΗO�C�<fnԕ�Ӿ��	     ��t����W���~Uo\q���r �vE���Y�������?��HLª����Zkg�X�g���&��̤�-��������������6z��XivvNuGە�¾�,�P��X�Œ�IH�bj�I##�bl�F$&aI���J?٪h�X���Mn$&�L�޶q�ԶhrrB���Ф����N�"��������������d� L,f��U:X۬ib1V��N~$&��b朝BOo�`7"1	�Y��X��c-,�TCs��I��$������;���0��l�F$&!��,��m�b,��HLB"s�H��&���ȍHL���gdM�H�5�I�{!��dƗ-�D��`����Gb֔ŷ�b��F$&���nXM,�bɎ�$��qƗC��}�p��I�!Sw�_z�*�T�
� ɶ��Z�s�tt�M      ���u���g���4>��6y �ҳ n�����������L$�`ؕHLByY�b>���X�M�'R%�N���XL�۴u��I�Z��9����@�����ֹ�I0̈́�#�}�:��Db��l�.U�Qid�X�M&&���ܣ�l��L,f.Z��ƶ�y�q�ΝHL���}���s�&�&{O��gЕHLB��<g�Us[�k�'�qnFb���F,�J&3>6�PZ��%T�Yjވ��#Fj���ms�ړ��l�Z�/�Y�g�x$&��HLB|1_�r՞0a;b16�GbN��I(*�T��2�'c��㝮DbL,f�ƕ:Xצ��1��#��EbJK��[b1�1A����!��e��rb1r3�`b1ј���I|nÑvW"1	��W�o�3;����Gbf�3�a>S��'b�g|i�9zܝHL��Ŭ_�RG�[��x�=���! ����u��#�     ���<�X�_Es�v9ϫ�7/ߥ�P� �-o-ۣ�|R��,�s����U��HL{'�x�I����m����=���L)to�eB����>�o�X����$�p��Zb1�0���@���V�X�zb161����nW#1	�K�䋕�DSv,�v$&��b�m*ס�V�=9!x�Db��ݍ�$�;�Ks�hn�`B��#1�FbL,f�Fg�Pע�ib16�"�PU�,>���'c/"1	9١����E��ؠ��O>g���?��XY��Gc��b$&۽HL����X�U⑘t����&X�mC�s٦1b1V0����ee�?�4�����/��d�#1	�X̆r�kU$�����Gb<_�]U��[Gw��#1\{��4��rgL��[��I0���+���OC������$�ehC%sܶ)�\;��	 ܲ�`���V�p�      <�v�q��`b�����4>�I�������ى������\djrnz"���b�O�f���~�?�y�gu��遴��@zFV0������/"���a]^�W�6�JH>/#1	��
�F���ݷ��e$&a>�J�ꚸ���^��ܟd��~]���4����x�,�=��I$&!�X�5���$���idtT������eKMԶ�X���&�����~�U�S�b�d"1].���w��ȗ��ss{'���q�w��αu�ty�I�^�,~.��G,�K�Q!����S�s��i=��H���D ���ҧ��W��!FꥩȬ�뻔��ݾ��b|&�Ъh4*x���.O"1	&c�=�uƗ�H=�e$&aEIn|&U���n�$B�
�u}��5kfzZ�Noߨ�UzȻk���ķ�b��e$&��b6U�T�_�1��RKۀ3���V�s꺡�Du'D,�c^Fb�܆��V�h}�K��g�����h$6<3931;��NOL�͌�Ţ��ٹ�I_@�����>(H����23��������?��{]Y�Z}��     xl�n�V}QO��O�/��l���f
����:'&��G�Gf�k�g�L�f�O�<�����{5���_�`{8<=ݟ��y��(HϮ(N�/*
�R�9Žy�n�K�������HL�"�b>utw�!�`�nݰ�X���:�<��$T�-����o�X�L$�p������f�%�/�7�*�y��޼���R�m��ww����{<��$�XL�W��Fb1^1���L��f��M�b�44<�y$&��� �%�x$�_�[0�|1s�I����&3�q$&��bY||��O,��HLm��K�ټ�\5�Z�q/מ�����i$&!>�\_��GE,�#��s����4�PT��j�$�!��H�y~pƗ�7��`m�&&����cS���/��ZiIn|K,�;&��a�4!�_n߰�X��z��448�]x��bb򩳛�x��HLBvV��8��������hm��̴g���D,��DT�CÂ�l��$�gh��r�ou��mH��yښ�F8�E�s����tod�{02~lln���\�@dr��o�?N���}�W/\�!ߙ���ف�k
ҳ�������>o�=����}Ё�     x�o������-w���e�����L��3<3m����yzxv���YS?��}����Z����gs�w��{?������,
�_���aUVqN��꧔�>hř���WBr�#1�vDb*V�狩��	Un�_��aE$&�,.ݲ~u��[��L�t�|$fҊHL���Dc�� �7��Ix��[��b\6����l�sl�XF,�&��ح�l�g$/ɖ/V��Mmο�`�M�G;��a�x"�ٸR��h�9��{�#1�VDbL,&�3w���cS$&!�ٸ�9o �6�"1	�k�ŷ�b�eS$&�D�T��Y�G,�U&��z�IH�bj�I##�b�d"1�OtX�I0��*��q��#㦣'����$�}�_�q��Ĵ��[�I0�������!���a��=�!��C�-��D��#1��������UE�B�:{z���I0��MU�t�x3���H�L$�`Ў9��Tvc�
՞����I��b*˜�N��$zW��©'27�����������O�L��7ox0)w'����7:������W�qᲜhڕy��K���m]�Y�$�g�w�}ЁB1     �s&��SxU�_��|\vQ�e3������y�g�y������w��M}o����~r}���u6���|�u��|Y+�(|ce���L;>�ER�a���A�C��#��l��$�)/�!����~��D*��%�I���[&#���m탚�O��g����ֺb՝�jl|PH��٨jN�� 7,��ehCe��~0�&T���HLB"SSצ�a���HL²�ي�LG�}�q�x��2��ٵk�O�f��^g�,�s�|$f��HLª����剦.�5G:���$��Amް�9o`|�x$ft\��]�K��b��q�OH���>R�a�"��YoƗǛ���M-vEb�9��R���GY���HL��,�7,)�t��C����ĄdM$&!�9P�C*v��XĺHLBYI^||y��]p�m����x�t�֚sHƗn�������s֮^ߞl�F8n0�K�"1	�s��U�:���'7��h&2mM$&!��;���s�`"1�'����$d�z]���d|���+�5o�pj�͜����xd�{o�?����ݫ�7'�_x�w������%iyo��.�Rηo`�g�AU9�:>ʵ     �3u���Y1��C��l_��㪀ϯ���-,n&�8����ɑ���c�?&��}��Y67��{�9/�5������[�WV�Ȱk� LN0C��w<!,�����M��]�%~[Z0��4'���`M�rsB����rs���/&$��ЄN6�*��������|f�������g�8�{�a�,�L���a�ͤ5{w�q"G�N3!���������
��58l���p���霰SBCs���œ����媵üW�x�L�ȬԴ8�K�>�B!�fag���͇ FF�=N��嫥ݜ�F����X}�,���p8]��Y<b��u�x깦x\��kO����Y;���oD�4�94[+7;K~�����2�}Ҍ/}�xߐ���<��3�ZچT�4��KO�9�3�l7�W1�L��9=�7����o�^8=�y���X�
��V�/���%�_&��Ĵ׵[�miii�mp�3����f��27O�`|�l�jl��&�-+;��.y����/�G����a>���{�ŭozd��X����_���������>�sw�Ͼ�Ї�zѻJ��W��\ʵ�x����=����     �4�����G�g~�E�+dn��z��%U.�ɹH��H�Ѷ��O����t����O���M��(ܷ6{�{�rJm��^���أ�v>��x��Є�x�IJ�w��[���3 Ƴ�:M���0;;����.H�w�d�����϶	0�e�u�����|M� ��}$� ������������.���^P{�W�108�Ǚۀ<�%�h��? ��/OMKB��y�X|���N�v���vgo�/��w_J��q�/�����y��V/��pYF�u��Vo�ӄ�圢M�v�W�bn     �O�P��~(�\g:υr�	3`q���n��eb������Es{�*�7����KW�|~[ޚ!?�Ţ8��=E�p�              �����=
���1:3=8��h���5w���Z$���?�_���������7.�(�}{~�ٹ�L��(�}~]�b����     x��\�<���>���_���U��)�Ɖ����/��}�\p�"�͏=�sg�ss1}E�;v�=;3�	)��ҽ�b               NQY��..�!,��#�����eb��t��瞏>X�lλ��gf~�5k�X�宨���ŧ�{-����      <R��k���Z���B_Lg��s�m�{���>�7up����7u��Q�B^��~����e�ܻ�ȯ��`Lj[�S�Xi               N-���Tf0]Hm�3��GN��k��]�޸H���8���7}0ky�K��}���<�1),#��KKN�?�=,      ��d!�b<�_/��s�ۨ�p�X.Ю�j!u�O��>=x����n�ʾ�D���T���e�������p}E���_������-+�$              p�1�/[��z,���t��ct����T���o��Ʉ���{�t�-˳��㮢���tn���.[�K?lT��)uo_     `�X<s������V�9�����k��(27�'��G�������{��G�ͦ�v�۶��FUvi��rvU� ����1              �԰#�����'������Ǉ;����/z!�s�{�t��ʼ�tZ~E���Z�T�$���*���1     x�,�3�5��n� �_�FH=�c���|��>������k������Go{��^��c9i~!e}�~�v����               pj��d��zz"C3O���ۯ���?腀N�շ_z��U_^�^�.���Kv�     ^Z��\_V�����og���*�VQ(GH�sS�G�j��׵����wgTxY�r�On���77���ּ5+��a.�������               ���e��*!uDcQ=6p�ѮK�q����q������?�e���̢�{̍���(�����     �'��<�Pp����u���x��:ǻF�8�>��o�^�{>�`��)��mo���6ߐ��	�+iK�jn               ��OS�RC����#�u7�q�Ͼ*�b/�u�^u�%�?3Ý���4�z&�sA�k�	     �#{D(��9�q�r���z��y�Q�N��\,������Co�o��«�kr���"��3�O�d��ֻ�d�              �E�����ӄ���PCS�T�Y߹�?څW�Ϋ�;"��.�5���]T�C?h}X1�     �{O��P�O��y}���������LF�_s��W��s������gzYg����,ٸ[���%�s2C���              ��-o�����o�:p����}�
�;Wǃ;kn���}���[�<��Z.ж�5:0�       l�>�Ǭ����i�[/�s�.,��n�����'�����k|ZXp��o���9󆯿���-����?M�S���mӏ;�               ���wv������5w^��I����˕c�E9w���B���b��      �֐*�m�����i�b���r-K��U3���\�a�����'$՗?�㫦�~�­w凲��n�s�l&              �H��Ӵ��Z�W�d���CG^��kŤ�$3!��;��ڕ����̥���,\�p ���i     �ί�"����i�[/|��͂��8v�׭�;���?+��Ϋ񭙯�՟U���႐`�9+�,=_=�!              `q�]T.�N�F��5m���_�
����_=��rl�x�����K���Uz��      \������^
�ܬ,�T�Ƌ����E��b1��?���~����}��MU��TZ�U�-X�����%����G              ���%��V��[���߳��	�U߼���+�]Q6����5���9�+s��̈́b     �7b�*��PLT[�ߍݚ�ZE��.&�`ϡ��U?�\��w���1x�6F;�6�$W��9�b               ��@H�T
�y~��阚6ܻo�������7�}Wl���fG��*�*�V)3���و      \F(�/�b�ڢ�;/zv�&�.&��|�y��{���u�U�b���W�	֨�.UI�@]S�              �Ⱛ�Z!�`�g����e��}�gO�X̦}�6<;^���j�`��/�]��u�!     ��\7(__֐���B1Qm�/�/���u�B1�y���?���w���g���?�k�W�V��|:g�f�S��              ��p��-�]�l$c�}��E���+�j��ѝ���k��d3�     �����l\��^��n�[���,�����g?|��u����C���&�4t�,sIX��9K	�               ,��t�(�ya�������Db�s���˺�-��i'��^!X��òa��M	     �U1U�P��^
���	��)� ����}����Q�ַ?�'}_
�y���O�r����e-ײ�<�D�              �Զ3�R!�tmqr�s��`��{o�O��R��o����:�Tf�(<��jg�:����      \�j�U�}5{�/h.����-ݵ�3g
ֻ�����%%;�%+�	�ۑ�N��~V               Hm�0��=�����N����C���v�X�ߥ��	f.	�ϙ�:�b     �����ܨB�97�/V.Ҋ�B�{��=OO�o�o��i!%|�_�8����Pr���}~�[�V�              Hq>�O;
�	������?rѽ7�TH	�~�����K�w>������YXߧ�b1     ��G(�m��;��wRZ��������K���>!��v�����od�{��-
�zM~����fcs              @j��*Qa(G�V����{��|��_�ZH)w_�����C������pCTo�e��i'�:     �"B1.��u'SH(�k����j�����������.9jjޚ��L�LF ]rW�f�I               HM�s3T+<�w���]���R�m���y�Ⱥ蜥�_+xjg~%�     ඕڧ��\1��i�|�}��?M��V�z���on���������}�m�Y�Qذ$�<c>$              ��v����Ѷ���MJ�	�뱎���ۺ�s�
Ϝ^X��q_a     ઠ�T�l�W$"��~��y��x�y�g��}�R!��s����ۃ׿��;�>����ේ               ROf0]�s���LFk�.�{�7�BJۿo���;��_�Y�lN03ɷ2��!g���a��N	     �5i�fI����P�OE�~���LE#�g����}L�����΢o�����g	�X�Y��P���G              ��򚼵
��w�?�������¢`~��wf|�ŧ�"x"��k{~��     �k��,�K�/l�$������H_�������@�-K�3�f���|ڔ�J�               R���Ղw�l���?�UXT�z�O�����wlϯX-xbs�*B1     �mIo��%��b�Vg�h�}�s�Jaѹ�}��B__]�Qt���ܷ)��P              @
ڐ�R����D��H��E�v����쒺�`&��=�1�\      ���qS"S��Y�]� O�Dg�l��w�߷VX��qݿ{�7o�]�~��:.�              ��t�*�Ko<�[{�=}�VX��s݃ǋ���͋���a�uk���o�<57-      �	���ٻ8��:���S����s�ؓ�a$��we�^W���껫��k���꾬CXT\��ADǰ
�����9����sj�0��z����OS�a�j��~�<O=�wfC1�*��0!�B����_�w��	J����%��3=��J�L[j�
�Ob,�              �5��1���L��v������{݊��}`yh^��Q���WW-��&�     �!�xd�x��*�O���PL!L$#����傒��u?�o�;�����Wub}��8q\               P�U�ǽL�k�D�Mw���
J����/���!��Y��[	�      �R/p�G��?�U7{AoM�B��?���^��^AYx~`��5U×/6VuJ�bB1               Ed]�PL!<?q���7=�5AY���ǿ���[��,_.pԺ�E  ��ʷJj<5bx�>��HjDF
 ��4㱾C*�`i�YB��Y�����A��Ӷ'����?,6�?G��^,�-               (��P�r1Tǥ�i9�BPV�c��1��k��#pκ���2\�5�  ��㱎��W�>Yg�#kHee�TUUI1x~�yB1 P����>�dů�	ְ�^/L��������?z뺇Z?�,�8����4               z[l�JO��Y�O{遛v?-(+�����߼ok����=��X�   ��U�U�����1D8� �Cm���#.��@��P��Y=ё��S���}���.�|^���; M�j�O               ��4�"pV"��c�W�RWr�������\�s�Yc�  �Ҳ5�U.�\,�  �b�q�G�����N�7�y���=iAY�u�_�����.�T
�4�L(              �,��b�N{i��ޯ~�ɗe����B�[�Y�j��1K�?   J�ߚ�S  ��y�����0�5�"��ƒәh������]l�E����yj�               @oK���L�3:���2����+wb��4��<   �"`����� ����1�X���ٚ��R�	���T�c��=�������O����
��(              @QXʾOG�����'����n��Ě��n����:  ��qA�� @[�����
������d6%}�ɛe�ᶇ���|wScͥGP[              П}!�_X��㑁�%��xl��խ�$pD��Z�<2��	   ��z�z @s�b��x�T��KC����o����>��] KWb���l�R��J�Tԋ��H�L               �d�q7C����d�i���D`��⟇���
�$�,{';   ��g��Ϲ�  ���o{�UQ�����ݪ|I�Y�����?�[���WN{pY��%ʹ�,
5ʱ�~              ������Qf�~��mg�<�gV��?kj��@���B1   ��c}B� �=C�r߄b�Q���F�3��{n|t� ���oC���
�ZA(              @g���������*���Ϙb^�����     �ң4��8�h��i�@r���Ls�o+���;�9P+               ��=�s,20��-O�(��<x�Ϝ�Ъ��y�����     Pj��b�ޠT��gD'n����H����#[jV�(���               Z#��������	����C�.(G     ��(�Lp�`b"y��������׶�ȭ�|p              �+�0�����KN�� �`l������Z�1��L�      �e�J��9>=�O��0����$o�}����               tU�	������y�cO�O��ǟ|�܇�F[CMA�R>k̳Ǿ�Ԍ      �4(Ŵ&8e$5�-^��?�éӿ�`xmxq�@�&���d̬               @/��qwLOl�Y^Gw|���Pӹ�챏P     @�P�i���KdRID��u�����/�\���i��e0>!               �{ܝ3���� �c49��uC(�-�ye�[      Pԅb��;�#28��-{�R�u��f�n��q@���P              ��Z���x6i���ud��_M4�����      J��PL��Z��prr� o`�g�D�"f�<�@�FX               ��y:�+2<��U{���{��n������jJq~     @iQ���ꍧ"��~���9�];�6��Q�T�7$               ��<�1��+�ILL�_Y��\�Ra��     ()JB1�aH��B��i��F�M��0��ڻV�<�R,�              ���w'L$�?�$L&�OZ7�bc�;     @iQ�	���1��FS���o�I� 'a:���Q.��               Z����%\��pf��Ǭ��(U�%     `�ַ���Y(v�\�K.�d*��$SEm����NR,��m�����|�              ��0���Q����� 'ၛv?}ٷO7C�!P��     ����W�t��=�����x %���1���$-9��y	3�򳈮P�[!               �O�<��OL0���y�e8�     ��l62���������h:v@����֖����/6�	�BaoH               ��
�O|����x��Td@�9�^3����<����$     ���Q��i�z�b�	�8"�I�`�R�q�P�Ba�               ��b�Έ�����L:�cݬ(e��C(     �;�4C�a���ń\�z�L�Y�`*�n�����              �M��=�N�e���h*��9O�c      ��a�|z�C1^���ū��W8�� sM';��-e��� 욘               @^�W�^�L�`���'P��f     0��� �C1n�Z3�x����������(eGb�⒴d               z`��3R��1� �J�����      ��B=�a��bX@Rn&O0Gi3K(�����               ]����h�� s�N�f�      ��f��Q����)	�x��+����Q*��(�5<��               @"	�eͬtF��WƜDf���b�!;A�,x9�     @ØW���f�v�$�u)yX�J2��B�9��@9bY               za�z�l��Ӷ'-�<��p�C�^-�O�c      (w�����LӬ,��\.�C1�֕�f�,�c�2����              ����PUKg�� oBZ2�k�(�     �]6�]n�[�r�\�z,%+=B1�e�$�9˘��r��               z��ߩZ��������	Ũ��b�      ��ܑ;v�����)�43̑�4#�.j�               :q�K�VV��b�d�Lֺ�T!��    �rgƊ>}G>L�JOVX�UΠ���s�@���               �=�`�;���v�d�V1  �`^�<�w뽂�c�f�\:�R�l�e (Iy� �;�cǎ�I�w��p:��`JB1)3-P�-�1w�[B�RY�@               ���$(�7��)��kG��� @9�z��o��-   �����iI$o%�v����|0%��4Hʹ\�b0w.�T
�K�A"              �V�㮞��"��7��kG9bY  �'��#�P�@  (	>�O����b���\|���=ǺY+��f��M{>SIl$�M��n� s�1�j�r|�              �����sy�}�M�<�vc�;  ����JUU�   �����\ozz�����|�;�n�l}��z�z1M���3����}�;�N�nS�T��)�PH�U�|̑+�Y,P�1              @/)"	�y]��]ۛ�v��!N�w���c��st0Ĳ  (/.�K*++  �T�Q�`0(�h�O��=����x<�J$����4�і�2zQ�:6�^y�?�ꪫ���JB13+P+��{�#�˽H���               zI�q�')+�B18i��{�@9.�
 @y�O�6C   JY �x<.v���^i��H$.�d2[��%�h�%��|�ֱY^K4JB1Dԫ�T��Ɯ�ܞ�r\q              @/D��s��Y7��$.��r�q �|؁��'   ����K$���b��oё��}<ߏ�&��r^�G���+���#�$�˻H�T�̊)yz              �-J���>�g� s�s�qc   ���Qr�0  ��t?��#~.������*��$��]�����*O�P�b�L\               ��H�=�N���0!O`�@9�@  ʇ��  �r���O ��꫻���JB1S��@=�ۻɺyH���V���N�               za��3��R� ��/(� @�0MS   ʅ��>>��V�K(��Uxk��:oe�@��4�              �nf�qɚYqz_a��U�+�0Uފ�R��5��  (�tZ   ʅ��>�@`�ꫯ�G�c�	�JpD�7�F����/m_Z�r��$�              ��\(!��7(P��W� �4�k�JM�c�P  (�l6w´ǣ��a   �$�Iё��2}>��T=��P�G4�����U���	�c�              ��d:J(F��@���9����?9(���{.�W��f��� @���bRUU%   �,�J�y:
����k~���,�ٵa�4�0�:��5;�v�m{�U;��Jw���XD              ��T�}��֗���aݽO�7P�q�睨�w  ʏ}Ҵ����  �R��f%��n쵮����_s�5��|%���i��f�R�� R%��#��ԟYw�!����6���D               -KpF�Sq���I�t��c� �<١�4%
  @)I��233������񘕕���ꪫ����R��S���zB�B18	*Z�M�              ��g4��[8	��3�M�c  �S<�d2)�@@�^��\.1C   ����d2�H$r�7���������\q�?q����b�R�2��N�VC |� o���_���
�O�               �3����0X�@���(P?O��x�� �rf�T��  P����̟?�=]tQĩ�U�����p�@�E�����JO�JJ����               �3���W�{��u�Y����x����Y�r����     @�؁�P(t�����|�?w����b�,�;��W����;�q�#���@��#�               @O�q�y:%쪺޺!��T�����q     ���cVTT�X]]�\~��{
��P���q��Ni�U�w�P^��P�
�r���2I              �~���y��x�����L0�     �Y^�����]��WZ[[?��w�k�п'e��j�Y�;W�װs����������wd              �k81)Y3+.�%PkE�y;�v�m{$*������W�k(gZ_C�I     �s����xb����������Vcc�#�\rIB4�,Aq�9�+��]���k���W���ڛ� �              �������4��jU����9�	����:��S��(7��ʍ}      ��0�t(z޺�{����v'��;b�f��r�X�������D^���R�9e�{1)cf�Mm]9�ϸ�*�����e���� ���淄e���T��}_�d�r�}D���.zo��*.I�˥�g|�S��5-i>Sj�z���J �]��9�1*���m;g��٤=1]u�IgOLLS���u-�����#	9r|L�f�u|>�l��"n��?t�+��cD���
����-�;#^��s���H��H�j��qd��>��1C����PR��=�4���[��e�дtt�H"�q�JK�Is�_뵧d*-��cȑ1旪��V3-��"��c����R�u��$\钀���h,%G�Ge|�cH�����������@��O](~���ˉɸ���ǐ*���~u�����!ۿ�#�G�o��'��9c�5�����C#3r�{Z�q��ί�-A��i{o�56�0�T��g�{����̞�	9�ɭIB�5+����e���/c��u�0*cz�{JAQ�/���e/���3'���z{;�����	a�y      ��0��Ν;�JQ��#1v,�9P#Poq�����]�߻���/p�`bB�����q�j���i��ʎ���,;g���A��c266�e,Ǝ�$�Q�z�G���R���-c1v$��XL��r������>I&bZ�b�HL6���N�d��fٻ�S�X��LBF���'�{�*�ϧk����cH��.9��&$�M�r�X��'�ّ���)�u��B9�=�\e�/k����Ǻ���268a��ZI��284�e,Ǝ�Dcɚ��y���s�Z�O�r�Ɏ�t�Z����v�|���h$�e,Ǝ�d2���M����R�ɖM����ů��|v$�w`�z������N_&O?�n��yB��k6�������.���G{��_ڑ���	֥`/C�����_�2c���uq��-5�r��?0�e,fp$"3�1���VK��ކ_��4�_ڑ���!��Zp��-�?8.3�-c1����L�~��kB%��-gnY.�<w���_ڑ����9㴥�܋bf��_�w��z��t2��tb�:�p��n�8����pJ�ߺ�m5�*,8��       ��<�&���@EY(��!��y���u�������V����鋎
^����23�q{��v�`;fͪ9xؔ�I�b1}�Db�V���3V����*3����[*[Nm��^��.�I$�qu�!�pJ�v�;38<n��c,&����c2B
�9�sKrG�����ĸ���p�1\.-c1v$�h�u�)�NZ��)w�[,f6chxQ��YǍ:�bf#1�)	�S6��H^�߭],��w<��s��*d����k����0�t��y�����b�HP8������B�b1����qY�:�b�����a�}"k;�lIc�V�X���L.���9�ކ�k��#1ǻ���i�-��z�����"1Q"1
}rƖ��bf#1�/��uˉ���:��n�'�7�~O��������u�o�����o��kC��<     P��<�ȳ�"��{ll̓�dr�UVVf���S'q�b�;�L4�4�>3([jV�s.ir�}κ{� �+�8%���cڣ��7�[,Ǝ��7Ry�4SkW͓��E��'ť�����)�'��BE�/�y�٣��P��KDb
K�X����)�b1��W�+eI�X̫#1p޼����%cGb&����n��WGb�<�b1��3Db
D�X̫#1p��y��N����_��MJ&C.��U�b1Db
K�X��.�$N�+�b1Db
G�X��"1�=�n�;35C$�t���.S�q���b��g���`Gb����t���)��[�j�ig~9'��tֲ����P^eYռ+�i�     @��?-���2����Dno��{ �����I}}�=f�hLi(�#�"���U/ڶ�m�gO�>遄�U�����#`��&�e2�]b1l�҃.�;��)$;s�酏��у.�"1��K,�H�t������N"1�f�b�Y����޳7����"1��/]b1Db��K,fpdFf���WH��bR�,�l�تE,Ǝ�$�1A����DS�7H$��r��g�����X�D$F�`M��%31��s��wʖ.��\$�c�z�`~YH��bG��%�����6���˧�4��=���韐D2F$��t���у.�;c2���	�Z^�x�����ͻ%({���U����!�     ��������v@&�L���b�4�>�"���՞�͡O��UP���Z�8���9+t,��H��F*m:�78%��:�H����H�&
����,�-:3!��B�bf#1�A$F���n��#1c������X��~uX��ؑ�c���/5Q�XL.�$>:cGb�{X{�E�c1�}�J��W�XL.3D$Fg�����"1�(t,&�%����b�������W$�E$F����ч����b~�kk~p�@�H�^
�!��B�b���б��n"1o�PbR"�����z��� T�9���e�����.���DӉܘ     P����������������QNY\�q!S�v����5����oN�b1٬�F**C$F?���ؑ��^����B�b���P��H4)��l��L!b1�HLǈ."1:)T,�H�~�X�;���ĸ9��J�b1���2�06h�P�"1z*T,�H�~
��ƒҗ{oh�P�"1�)T,�H�~N�bV:�!��B�b�F#Db4c�b�~�*�c1Db�T�XLO�$���b1�-�g�?�h,�H��
���6�&��7�4M��)�V�3N�Yv·������w	����ְ�f��Ǵ�sc     @9z�u�b_3Q�Ie����P����뮽�����ǿ!([K-�gS���#��7��X��9�9�F*M9��'�-�c1Db��t,��w�H������D���I|�r2���t�єӱ;3:a�
4�t,&kf�X��M9�!�/�c1v$��{X<�9�����Lq��fc1Ͽ�n7��HL� R]ٱ�_=}�:�wf�G$F_N�b&��22F$FGN�b�����X��xD�g��_j��XL�H���X̾}25=��ކށ)旚
����b����D,渘g�|\ �k'�Jw��lT}ɺ�A�Z`��S�	rP���     �$��[{t�P�Ö[�޺!S��j��-k��8�#��
�b1'��N$Fw�X�!��	��;#�5�b1�TZ�zFģ��o�S�;��$�r*C$�88���H�A$Fgv,&wտ���"1�s*���t؛�9�OgN�b���ϩX�l$�M$FkN�b��'%ɕ޵f�bN۴Ty,&�HI��'�i+�Ŵ�ўS�;3<6A$FcN�b���b1�c��&�3;�6{]��#P8�$S֯�/���XL���$��mЙS�"1�a�e��b���tކ���]�����W���ζ�M5K�#pTG�=�      �H}(&2(�7���zɒ��_t��ѣ���<������NʘY��ձ���A��^$֮V����h<�&�"0�y��c�l�#1��#�&ST�b:{�%�%ST�b��������Î]Uo����[U�"1��b1�yX�����).�c1C#3Db���X���:s"%ST�b�HLw�('�	ձ;c�)
�c1�3q�c��T�bNDb���	ձ"1����X�˕�b1���6ձ;�8EAu,&�$SLT�b:���M��5j���5wXw�����]��jv�9�xd@      Pz�/���8�e�dyx�.�n���\�낳6W/?E�(���T6-x��X�9g����u�������HUd�X��/�%���|�4%#SL�X̺5��;��3z�F��;��s�bJ~ǆH4A$��ر��E-242����� Sd�X�S����xot4B$��ر���D"��8?<6%6`;��sV�s/��c��M�)2v,fz&&�T�7�O�̈�ㆢa�b6m\"G���s�ޞ1"1EƎ�<�B�d�O���&F$��ر��K��0���ށaN�+2v,�ik~i�{~9%Sd�X��d�LLM�����'����K���|��^.֞�����IJ"��cONN�*"v,f˩K��ូ?vW�8{���yd��=��f�Db���Y�r������{���\,���b��<az���@$&_�E$mf��3:���u���>���{fecgێ��e���Q�EP�      �&�ž2ݓ[`��%p���%�w~�ݗ���������_�8��i����c�b���_��3�������d�l�$S�<^5c����ɽ_�S*E�����M���Wܮ�n�wO�j(F�IA���旼��Ϛ_zU�x=���%~ǎ�\��A6����Q26�&��(������i>+/Fn����؟3�Q{���ؐ��8��uY�
����Q����P�|^���>f&C����n�!�_��y���DH�)�I��YU�@��z_س�]{�u�hH	��h�W���aǣ��p�4     �R�|��^Xj����y��׆�%�Xw	Ŕ������͵�V	��S               P<Lw�)�3�V�;���7����k�8�ukݪ��w     ���H�y�t��XY9��cw���ۯ�ӂ��!��n������S              {��{�-pV�7�Zh�w���(��*o��`�d�      �49�90�%U��kW~��۶�Ӄ������~�m+*��7���}              �x�CEa�Y��o�p��?��nAɺ��^rz��͂����     @ir,��h��xV�<j�=WP���s���jWTP��               ��hbJ��~k��<�[N�]���m�ַ��e%��{u���?d�]�y��6��      �&GB1C�I�����]��k�|����oJ��ݵ�*V��P              @q���65�)���j��=��u�
Aəny顳*7�

�=�      �͑P�m�t�l�o8�m������v|�޶G���qÝ�~bK��5��90�":              @1�c
�j�((�s������_z��'�����ؾ�܆����`�      �6�B1/N�m�b
�5��^8�ۺ�6AI���Z�mX���a
c2��3              �����1A������'"muM�=��mm�<����0h��

�q�6     �R�X(�ٱ#b���(�s�ם{�]�ܲ���n�U��?��U9�3�?���Q1�/               ��ب���d^�NP+*�W����u�RA�;{~�VU.��@|\z�     ���Xdb$9%�!Yj�a}�[w��f�H<�՛�<,(Z����=��z�bAA=;~D               P��?"UP8okXw�G��껯��Ek��\{nú���8��      �:�B16;�@(���}U�ӫW<k�ky��ᤠ�\��K��ָ�C��2��&�	               �׳c�b
�c��u�5~[��oy�EAѹ���ok<�n�����C     (u��b�����&(�U�j�N�̺{���\���k�Ѵ�_�.Gt�'�TD               P�^�l�������B��U��4,��<����U{₢q���z����WE%��Rٴ�<�!      (m��f��H&.!w@PX�֭=�{�{�m�}�:AQ��m5g4�x��f]v�
               �-�Mɾ�N9�f���VVί���h�]#(���YY��FPp{�:%�I
      J��������&������2C�oܴ3qg�Ȯ��@kmmm.M��C-a��%              P�}��b�pz���}��?���_&����w�cg֮� �{�     ʃ����c��h�c������Kޑ>r�M?��@[��C��\�v�@����               ?{��Υ��a[��Kw'��_>������]v�;��_,��o�      J�㡘�=(]�#)A�<ƅM��C���q��O<&�Χ���'ή_{�@��/Y3+               (~��Q9�e�A���M�o���N��_�ܸ�O_ؼ����`�a=�     @�s<3��ɋ���ڕ=T{��w�l�~���/���_
��{��[�lZ�@+?�'               (?�G(F#��i/j��?�wH�Λ~�wm�p祟�������?��g��q     (Y���	���v��r�O�;�w��O

�w��7�k�x�@+��?�%               (?�+��|1C�;��e�K2w������.����S?�#��_��     (Y����A���BAZ/����¦�v�w~���+(�����Ƕ�o�X�;t�5�              ������~YY9_���+�l�{�.W�n����Mw^ֶ���������^鋍	      �CAV�f�qy~�l�[-�K�7�:��w�������Q�ڶy�-���Y�k������              ��c_P�P�~<�[.j��)�=��ۮ��u��r�{�9�q�N�����({�     �I�R��":�=U{��w���U�.��;n��g�����7����Z�l�@K#�)90�%P+�HI4�����^I&E&�LK&���C�1\.1�YA�'�JƆ��_b񔠸$�3���̚.럆�m
�GR��೎ҩ��x��I���B~�=���`24���Z���^�d�7Uǐ�O�񨠸$)I���zp�ݒ����j%��旑(�O��~=�{��^�2��H��Ȣ�L�Y�������x�fV���/����5.���G2�T��d�/��/�I*��^)�������׋Q�z=$����!k��q�N<�n�ɾ��=��f����n��PL������+�$���w������/֞����^���B���%�7��W�j_�����x�tȧ�~��׸�}�\��~_���     @�(خ��FI�L��`㋎n�\�r������~n翿O���r�Ƴ��ri��J������Ǖ��R��9,-���Qhn���G\261.(�_���
%��-�W�vI�XLQ�����䌒����R^>�+3�iAqػ�GZ�J��vI{W��)�SbfRJƆ������SIb1���d���Z���cۯ/��-���b�DG稄*������
�����d���Lf���~%��c�r�%#cc���ʑA����a���v����.b1Ebz&!#���֞���#S��/������\R��~�K�t�p�N���T"�dlh�Y��.�ŉ�{~��^%�K�^_^�[:{�9ɬHt��Y�!!cCM�B^>�e�[X{*v$�C}2�I����1��^4*(G�Im�W��/�����W�$�%Pf�	S6���������8�;�'Muj�6�=9t���Ebd,"�XL���XW)/�h,"�߉�������'��%���=)4���C3���j�@?���;ֿ�yϱ�W޶��o�3!P��3�YU���i5˗�e�Y�q~   �B�d�=�G���C��1���:����}��+*Ԭ# �W�*-�L\~5zP�5l�ɾ"�y���[�@�c_��̯]�{H�w�����/����&i�ɡ�ؑ�c�����:���z��9xD��;ST7,��TȚ����n1���tfGbF%X�U��.kpظn��t�G"����HLu���	ۂ�p�X���H��tD|>��Ƿ� �Ni�Ɔ.I$�j��Nl�������?k��Z1�Y�"�9;cf��v�9�2�ʆ���� ��ّ��G�$\�W�kV4ˡc����btgGb*|���p@֭ZL,�ؑ���a	խ=�_�@^>�#3�/�gGb��Ԭ5ؚr����b������_�Z���t�by9w2_T���HLm��c�����F,Fv$&�L�ǣf��s6��Ɔ��d~���HLuX�ذzyS�Xrh�X���H��c*�Õ~9e�bb1E IHWװT��/�, S$�HL8�noC}]PV�"b1E��Č���K5ǐ�g��-"Sf#1��*�6T�a}�w����Џ�^$�9;\���������v�\�wW�y�[���di�YAY����   �0����������~/3��o����G  ����)��PL�T���>Z��C�s�M���E[[�+:�7��p��=����?�gz�Xd@���H̬�X́#Y�����+}RY��%�Y�P^9�C,FS'"1c�"1��X̦u��hNu$f����/�w�ѕ�H̬\,f�bb1s"3k��z���詣Km$f�}\b�b^>�!�4'��Ȏ�:��$�Y��5K&+26N,FW�H��P���Y�r��r�;we�Gu$f��e�Ƶ�ek~9e~�+Ց�Yv,�4��vb1��(��̲c1���wK,N,FG���~g�v,ƚ^JW�]�􍟈ĸծ=�b1�X��bt�D$f֪eM�@��(�]���̲c1��,����$�a�IGv$�Sa$f���:3ˎŬ�Er�X��TGbf��b^<�%1b�Zr"3k~K8����X�2?zY�]�]n��x�+j��?��~���'A�ܸ�ҿ�ְ�﫼.��ٔ��+    �w����7�yR{����������햚��\8f���A���	 �+h(楩v鍏ʂ@�@o����;������M�\���k��zV��AQ�a��5r����rf�bo�Z�r�<l���@/�K��#N폯�����Qb1��]$ƙ���X����e&�շt���^��rnak~s8������U�q*3�w��nI$b}8�����.wK,F?�HLF}$f��ٸv	�9���b�+������M0�ԍ�	8��U[]!kV�ёS��Y�X�:b1��kCV���_67T�a.�#�btcGbF�&�Gbfٱ���|��$��R+��f.vn~ٺ�6wK,F?v$&��+���
<�~m��=�%�tR��t:#_�מV/o���яS��YU�~ٰ�X������"�7�"1���?��cݒ5���dԡH�,���S�-&�!'#1��b1�t�b1�<�d���ra�f����e-g�c��5<{��?�C�ނ�m;�*{{�)�4���b���}�1   ��&&&����v^��{GGGs�JEE��c^����  �SAC1�ƻ</W/�P�?��+�7o|_������=x�Gsv���Ϸ7���xC֋D,��=#��O8���;�o�<9`�b�̧�W�K0��禹U�b�29���	�"1��XL���{$�d>]��Ĩ���Z�R��%���!g#1�r�����@,F���̲c1�aJ���@NGbfٱ�k���W�$��|Z�Eb�8����_��'��%�}8��e�b֮\l����h��H̬\,攅��@�L3�Ԇӑ�YM��bʉXg����H�,����)�]�k>{4��c1��R:{�����H̬��r�bb1�#1:��e�b�a�X�6���̲c1�����N�d�_� KJGװT����@,F?�_q63��ې�.���=��JPx�1������g��O!"1��T���/����R���%S$���ֺ՛��*�������	��;��8�f���8����    �{��G%�H8�\�X,�����G���zsјW�c����v�3p �s
��=1�\�z�x�l����%���5�S��/\��Nʇ��}�P�׬X�r��g�{%�q栽�ؑ��G���̲׭l�}��2���w'�q�g���*�lm�e��歽t�$!�sg��d2� 	�;���\Ba0!��Y +�,$���ֱ,��h�w��U�JK-���9B-�ݒU�9U��>o�Jǖ���S�=�}��2��MCb\i���肪���UѤ!1S����h�b�����D�Bb,��q�L�-���)Z!1����+�v�loQ�M�YND���r��P��C��4a1�v?$f[����Ú��a1U����NHLvdCb,�� K�����NH�%/'݄�t����E��Č��IVFt�=i鹆
��9!�k+��VH���8+�_�b� Z!1�����t���a1�d����F�RUU�K AJ�qh��h��Xv�b����m��͐˙S%~��/�+Z!1���4�?s��А���i�VXL[��2k�NCb�3��䲴(St~IXL�-��eff1�!1������0���h��X*���<wd�0�P�Z���9�Y"p���bW���e�Ͽ>�q��_�'P�s���|"��S�^^�C��I��    �������;��ޖ��i3��r�v�ctX�2��Œ��-  ����ŭUi^�'
Α��Jx]ɥ7���m�c��o����
���w�3q���_�����s�3�S��#��4I����o:[&��	�^q����d�G/$�RX�!g����(�vH��t~�+�;]c��N��h�vH���X��LXL��ĤD7\4-5I.֟��]#��D�?��D���r�D�$H@&�g�����4�UJ[����y���ݐ����c�����%At���Ԅ�/��S)]}c��D����ep_<�PNXL��uD7$Ƣa1-�#,&j��c1a1���D���'���g�b�'�!1����.�b��!1���J�1an���h��nH�E�b�TIa�Q��lG5$Ƣ�⹳��D[�Cb,�(7a�ܿ�����^H�E�b.4����D�Bb,U:��a��M
a1������5?(pm^�=E���X��y_����}�O/���C�ו���/wF�b�K�Z9'   ���ݻ�9�x<fLNN>�mw����������: �\��\�^��IP�C��T�f�?s�Ew�7f����"�w��?����$w��_�u�h=�^���qA��%$�b�b�4,& �TE����D�˼Q�b�H��qv	��h����J��9&a1�v�cL���@�b��0a1g��KZZ2a1Qb�">K͉��!A��g�e��KVF����������Ґ�����Xt^SW{\��daiQYv	���纤�T�t0��4��~H��
���9.kk���2!16���iX��\F&�Ϙ_F�	���~H�E�b��Wʝ����D�����&��qh�0���X2ҿ�9"��mA��)$�Rw�T��	���II
�f~���n�b:	��8��AH�e',�[d��g��K��/*����H�KH�%Y�6v
��T���221|f�s�X����'_/�	�y���������I퇏�������_���;��篽z6���sO�$P��Hހ/x��#    "ohhHb��Bd���$''g'D&//o'D���HRS�s] �-�Z�\�Iς��
Σ����pv�b�诲?5���3O�җ�zE�[��?P�y��.䜬�⹳}~� t�cїiS]��w'8nAd�-$�RT��o��h��-#���UH�E��/6T���QY][D��Bb,��r�g�Ad�-$�b����g��c��ԉB���Ԭ 2F����6��$+3̈́Ŵ�豁 �H�[H�E�7��Ǥ�Odj�b�H����T��/�3��t�t�뱁�e$�-$Ƣa1*�Ŭ�"�n!1�������(��H�[H�E�O����旑�����"�|��'����%[��X�Ŝ�����3��"���tO�*$Ƣa1="���_F��Bb,y��bD#��
��ל����Y���!R�c)-ʒ�@��� +R4$��6Xa1w;�dy��a�_޳UH��*8�$�=5旡�����g������Ԑ]Uz:�칲�.�1�1��?��_�8��?{�jWɇ��~<5�^�i8��϶�{��~    ���%��|>Y\\4cpp���YYY;!2V���X� ��w0��OO>/�x�Ε����ڒ?>����U��G�����o.�Z����^��S�eu1���{������WgnBû퓶�	�t���=� VW�{E�:�qn�sR��&k{-��������b��`'�<�208m���zl8u�T�n]\�!����&L̮�Bn�K

dd|F^K��woIRS�dk۞��k���삆��s����ֈdf���PZ�++k[2A�N��̮JR��$��2p!!QNT��Y��������i�cCUy�,�n��nã�R\��=痩��R~�4�>1!z%᳹�ޞ)I��SU%����uAxu����4������HƧ�qh�յM�3��U�^{:&�}GB�zi�����,Y]͗��9Ax-,��+5A���~�=_{'+��̼�/������r뎽����Ž��Aqݫ'"�&��0C��9�LNN���R�7��2�4���k\2l|]ڬmXfmC$��kD�m����49V\,SB������HZ�}�'�J��K�6D­;㶞_��k�/C�S����J.
�#�+51Y�Ya��K��.z~la�?|�W��8�~��OU�<y%���i����i>5�m   y[[[��rwuuՌ����%''Kvv�NxL^^�N�Lqq���\
 �`�����[������f'���қ����]��K�9�8��X���s��w2��o�ϭ�I" &f|~�l��y3׉��Ve�q���x�ƈ jxt�@=��� ��g�@��p�m"mȢ{C��-�����1������w�P=��f �k�@�n�dum��%v4�0.��7�b��y���o`x�@1��?�k���Ҁ\�?-p6Hyea�y[�����k�3��~����e�a?�ǯ{eEF��_̯y<#)����Ǥ�5�  �h���<��,..�18��kiě���"c�X���� p0�	���o���OV�J�R3����U�}�?P�1�1���~��?&1��������,��S��r1Eb4(               ��S�&(&��'�������y��T�d�����_ṱ���w>-�_��W'7�d�JuF��r��i�{>=�    �YZZ2ch���.��E�1yyy;�2�X�f  ��&(F��T��h���`�?�H�ׯ�i�*g>z�����[������o~��)��w�3�^�-O/�ņܪ�L��c��ӷŽ�&               �_�܃2�vOj2�	bGbB��˭.����������|{z������,��?�K��Ն��W��P���֦���    ��J����199�����$���1�1��1V�LQQ����
 �[] \�Z�g����,�M'2J2�����s�çF=3_����ч����bSo�����3�XZ�O�f�^zE�+�1-���$I�               �N�]z�y���-�M�����W�����W��g=�kSߚ�v����+������gAr�/�d��*W�K�>5�msL   �D�����E3��r�v�cth���X���kl��"�J��4��LvyAp�)��M��T����읅��/������ۿ2�?������yNZֿ=����S���3���!�������               ��L��T��0-G�*]E��x}���_��󾡵��٭�/��?��_x�V4�lo���]�J�xsqj���,�-L͡j��\6�"    ��<����lKNN���l��1cʔ���� �4�;r�������gu��Q�Q��>��o=�T�ƽͅ�����+��oz�/|��	��}�;_�\S����I�o�Jr]-J�n��()�Nq%
��'ƾ)               ��|�����N�� ~hKpha�����O\�ύ/m�u�z=�^���ғ��Wo��g�彯���������ߓ���X�^TY��k��D���X    8��+���f>���r���a�ʤ�� ؑ-/���3򊂳��@�����4���������ѻ����_�z�6�����z�|	�Y����߿��$JRVR�d$$$&$&%O$�$&��&��RRJ��\�rS�r�Rs�Rm�2@��X��1               ,�{�E~��	)L�ħ�Ԝ��>��C���ɫ���Ս孵�U�gzÿ=���No������>�V�7��N�%���yRrbqb �8-1�XJbrizb��dWiNJF~aZvzfR:��1��b�A    �+8����c�����v������32�c�	 �b˄���{�N�ޢF,y�����%�|zB��g               �m˿-������	`�@�LW�K\E��Ӳ�$@�}<x��c   ��"$�<,D&))IrrrLh���hp�(STT$��� �bˠ�����Da�$&$
 D�w��wuB               ���x�U~��	)M� ���M�|y��     ����������lw�\;�1:4HFe��8
��Lx�幹v���� ��#��
               �o�'������ ����>'�~�     ����199�����d���6�1��1V�LII�� c��GF��W5IRB� @8}c�C��	               �R�2}K~��{�xz� @8Mo,�Wgn    {HII �^�,..�188��m������cdtX2V�Lzz� ���b&=���myC�c ���婱g               xo�'{N�s� 'm���    ����l�b�����/KKKf��Q.�k'<F���X�2�8!!A �>[Ũ�F������DR� �������
               �r�6sG~��{�:�T  ��g�ٻ   �^���eaaA�h�x<fLNN>�MÌv���Bdt�v �����M���ķ单� 5�oS>4�5               ���_~I�}�- ����/�/x�   `/�������^���Κ���������� }���  ���A1�cߔח\���\�P����eakE               ������,t�?+� �����R�    ��'Nȝ;wp"��c�����RSSMh��Ck�����D`����o˓�_�_9�c �2��(���.               �a���/ɕ�Ӓ��e� �����"    쩡�A���/��֖ �D��{����l)..�	��&���. "�1W���k�:~UsN ��ޜ��{ũ6S6%m;M�����)Y*`õ!�[ɒ�s�)�%Aĝ���|IHHķ���Y͑� ɽ�Ο��ՌU�Y�`)gI
�o�O�;_�O�S�%}���r��h�H O���-S|)�8<UX�^��bV]�������~�3ݒ��/�r���/�KB��e��%�d3mS2<赧�E�s�I�A�l3�����/�����5�$� ��������sq*mZ�����c� ��L|G&6�   �=i ���祵�U�x���b�����222vd������=�T���/ʟ^�y�� �m��|g�[���|�\m�*�-� ~��蕩�)Y�^����k-}MZ�Z$5�*�گI��1�y1]Hu��]Y�]�ӣ��b�B����Ι;���)��.K��b�x�O�Kk}�Yx{�����k�hҜG�~p���Y�7�+7�n�V�\�*��LA�(��ccR�Yn�#96�/�iil����^{J�T�4���d����ɩ�SR9S)�_Z��B����n�(�_Bz��-Y�\���z)],įقY�^���+{.�4����E6�7�J��Z�į��2X6(��R7T��2�m�l�kO���%m��e�
zN��T�TOUK�d� ~�\�f�MI��ʵ�6�3�������]?\/%s%
�1���K'{j������ 5[ �(�����c�    ���׾V:::��� ���u3���ؖ��$999;�1&c�Ijj� 8<G�e�_���g���K.
 <*_�/9�%q:���r�E��_��M:�ŝ���.�.�6O�K���ڱZ[ơ5ך�4���[����S��v/�R�U��k�ŧ��9i?�nk�ԍ�r��$���7���f�MYO[7�k�A
݅��������M�Z�]��go˅�& �E�9774�7�k���䕮+��N1_<�;�'E��D�	��/>����F�ѷ�������r��e��B�*ė죘/NY!�j#mÄI��a1�&��[u�dŵb�w�tI`( ����!�ׂo��tKk]�\�,���fw��}A���V��E�=��R5]0m��0ܠg�R1W����ҵI#�x��=o�ɛ1χ��7�K#�8e��*=w�s�ħ�!�������,�-ğ{E�������)�oS><������R �(>8�UY�m    {s�\��?����O~Rn����dqqь���m�5G���&@�
���d�sF���Kq���}Y���Jn
�<��L|G�צ%h��.���yE�<�ŋ�ݜw�,�4;�ŗ��,���b���w!��b��dus�M��4,�b������nm�����Ǝ��nλ���r�����	�ij6獻�ַʥ�K���+���9�F1_|ZM_�ֆ�}M���M�N�f� >�!�P��v��Z6R7̹�^{J��y���z�����}�[��~)���/�����@�������f�j/w]�D?a1�bo�E�i����w� ~�qA�[�6S0c4�����cw�E�6�s�Ϋ��a�W�0kNw�\��6X�pΌ�ď��%�]{�E_�J�N<�Bj��5sϊ�
A��*������x���1� ���^��L�    ����(KKK���O<"}�,//�1<<�����������͕�D֨ ~9.(fy{]�z�+�k�� �aMo,�Sc�J��"�˝�%ۓ-�q	"�\He�)�jľ�Bb,�ŗ�ZHe�b>-�;9qR�vwsދb��b�97�S7���?�vs��t~��n�w��b���h����y�[gnQ�'L7�]2�?��v����rFp~Y����
*��qU\t~�u/Bj��/����JGMǾ�t�a��ۘ_��;�l�)���n��5מʧ��M�!un�s������k׺�I���e��J�2�{CH-wO�5�Bw� ��T?BjY�]��3����DPq�/�t�����uE��i������CH-4/���Zh�_^*���_�/��T߫�6}�?6.�K���}���=�6IMp�} Q����>k�%    ��'�0a����essS �����ݻg�^III������� +P&55U�X�ȫ�_��%�.>'���Z	�p�����ےX�])�m/��y/����|޼��j{诡�/>��B*�ȱ�%���(�бl�x�tZ{��O������� ^���^�3_�_*f������ךkMn��4����b�Fچ)�|���)��;'����*��YCH���봘����r��"�|1�a!�����Y�v]��u:�Ǫ�!�P�Bj���VPq�67�c�^O���V����U��vҶTOVb��C���c�;��t�?I�^.���v�M��d�D8o�E&���CH-���r�lp~���2�d~���֥�K���+�M���v�mqg������
Į���Zh�^.�Ԣ��g�F8��a!�N7������5 ��ѯ����    p���&�����^:;;eaaA ����3�7��^o���|Qx��XGvv6��x��
԰�����Jb�)��ѐ��K�˴������rݜ��b��ڶ�a1,��9s�s�^�.A1_l;�B*�x�l'lK��|���9��|��]��/F�n�7^6$��_�o�ҙ/6=���^��{���I1_,�ߖ��� �|�b���rݜ�҂��b��w��9���ȕ�+��F��Xs�R����a�A{Bjѹ�����x�㒶E��X���D���1||�NNR���*�d�d�@�VCD��5˵��c�ACb,]'�L�o�\)��s�R�;�-�u�r����XtА˭3�X����!�8���_j�����z`A�9H��F8�MCH[�Zd#y�@�~�lD|)4Ez��t}C,���7�E�R�Q" pc25�-   �\�׽Ό��UY\\���%q��|��:�: G���f����Mw�������yyyf;`w��K�7��#���Ϟ|� ��Y�^������ij��bAl8h7�r�����b�Xr��t��>�/�v!�e�h��ә/v���^Z�g[�_��m��b�au,t�A�ӿΓ�/��y/����<o�"�~�^6�8y����)�~��S�+�XoBb�c1�|��r��b�Xr��ݴ�S���V�����6ܔ�����Xf
fL��	*&�4&���1�8\7g�h ��/]���
����ACH-#�GėL1_��ꑩ⃅�Z�>�t�;Bj��6�3��`BHO痹��_�e��sO3��3���!��'�hH�^����ah#�h�[Bj�Nl:l�E��>Q;Z˵�2P1 ����������?#�	��x8�c�Q�ge��k�    �+++ˌ���}�{<&���"&@F�e��}��������Y3��r�^ ��1V��>fm=���+�>3�yUQ���. x�?�������:NvHCB��s��p��漗;�-/�}A�y�U1@���GE1_�xԅT�̧A3MMt�CC2Zz�n�{iXL��f��vU\[�9�'�c>c�3_�0ݜ�s x&p��:�ǈ�vsޫ��w��f)�s��vs�k�u�����$)�$p.����Z���n��M1_�x�R��նQ�#4�TC$�)�k
�/;�J��b>��L�4ř�:��b>��h1.xh��Å�X�������&,&u;U�l:'hihy���_�/�$�TMU	��QCH-8t��\�&�>�f��QCH-R?X/���g{�R���B�I�N��!���'v<j�E���U�Pa11��Dp~Y�h�K'�Y��߻!���+ ����c���~   p&��Q\\,555l� �����P�X�F�~�crr�m��ɒ��mBc4<F_�:�ynn�$&r����j�/�����Ʌ�()���_F�Y薯ϵI���3Ig�l�L�LG]HeY�\�ֆV:�9�.�?6.�G�^�9�QRY�r��w�����蓉��#}-�k9�"WگH�f������^t�s>S�s��ݜ���-�� �4o����r��v��#���~�oU�T
��Q�9�e�o[L@�����W|�,�?*��w��P�LG!�P����ر�#��uE��)�s�ʹMinx���D�9�P��\G!�hP���\m�/��_:�QCH-�e���R=Q-p&Bz����xi&,�j�K�2!����}��CH-]5]
H�|)�pJ��Z�Z9�Ԣ�p���1�O#u���c�=��h��|�)�f.�s���F8:?in��C鿟�3h�y�yr�i��V��� �gjc1x���    �nB��:����|����&c���ssss��u�5a ^��9Y�����IJJ����������׳>OOO T��2�6-O�|M~�� �Z�^�?���W������|�\�,G�漗�ַ�"�b�G�tˏ���B1�s���^���,�|����n[��鶥� �H�J���P��4�������Gg>�2!1�we1�h!1]��AR�:�I��ߝFC��O?z7�*ė���j��������~�R�����(�s��<Pq�RK��6�������Fu4�!����-!���u�K=�$w5W�,�u�QwCBu�H��t~�4�D1����:̼"t~�|�ل���\gY�^2�p�2|lX�	^9=~Z�,�Āܪ�%+����X6R7��\�	�J��%T!����&l�b�B�,&���!�w���).w�ǉBBj��s���6�	�چ���>�k]��,&����!�N��m��v���ᅟ��� x1_�/�����bS    �04�";;ی���}����	�X]]}Q���ll��f��i��K��(�˵�C�d4@�z�Z\��bԧ'���y5r5�V ������Y�Z�x�W�'ۉ�R=U-p�Pus�K�u���CKh@L(RYL1�P���S������|Σ��9�7�����*��.K�z��B��y/:�9O��9屢����.�گI�&��N����:C�}���}�b>��'��f�MYOMH���5Q��$���RKWu�	$*�-8�	�	�����y/S���9�|����ܔb>g	uH�E�FK1���:�ԢA�Fz���dlf�a>o^�N��������kg���A�MhpC�BH-z?��_�doL,a�y:�?6n� B���_h�� ��ۦ�E�BH-k�5||�38�0�t�P��Zh��<6��tJ�&��bk���/O痹��_:M��||��� �����K��    @8h���
��z�;�1���d��t�s��Z�crr�m���cBc4<F�c�@���"IM��/^,&VY���}V����%'�Ee ����w�e�W 2\6ln���<)��Pws����w��ŖN�]�u�t�t��2})泿p�X����ۖvs�_�-]xK1�3�+$�Bg>�u7�t!�.���A����N�{�C��y/���c��sjhCH-V1��6�b�N�!�ˇe��H�~FoU�96T�����B��y���53���y�b>�3!�'�d&?�!�-�c~�8y��fؾ?�|��ҝ������Ody��6�?'�5�a���%��K�I�PמlN�!o6�>�Բ���T����6�W��4�Iږ��j��m�l�kO�Z۠�K�4�p�O�I�#��B#�Р�����}w�[n��M#W�Si�cy��!�J @i@�     Z���w(jjjؾ;HfuuU���Mx������n����Y��+��g^_:�'��O��V��h����'f*��V��?'�^�� #k3�����d���Ylyz���v�n�{i1�.��3���n�E�[He����vR�������X�c�`��i��3�YHE1������^Z��~�]���XliS������	~hgث�W%ӓ)����Is~����|�>���Ϯ���y/-�k>�L1��U�hI���W��k����d�97�/$Ƣ�%��[$BH-:������R�=�;��B1�������������*�;/K�'[`O���I������i��0� �'m8���"�a�9&�T�!ۯJ�v��~���1n�Ǉ�ϣ�}m�l��l��v���"W:�H���vdBHk�BjѰS�(�+%,Ʀ�Bj�i��u��b�
w��~���O��.�M2�9��Ƿ%����96    �]��y)�g'�B��h�����9��
O�C ^�kN������5���m^�%%%RTT�"���+��\O�E1u���.���M���� ~m���޿�-����Ƌ��"����^���y/:�ٗ�Fu��t�t�~&�|���T�̧�-5�b>{1ݶ4$&+rݶ���q�Q����n�{�g�S�gS��漟����}E����n'z9~l\�"�3��j��.���pws�K�כ����K�����G���Bj.6�'�(�3߫�E�u5�k�k�M$CH-Z4
H�<�|v����3w"��(泯H���v�ᦹ֐��'�=���H�)�o�W�������迋Ah������R�H5,Ƶ�؋�����?$�B#��z���H�m0k)��`~iC�!�tWw��'��O�BH-�N�p�(��[u�	!u�{��/�/��k��t��2�1/    �t.�ˌ���}�[A2������l�dv��v ���zw^[���/ږ��$999&4F�c���v��
%-���NswO�j�Kr.�T��@|z��?��Z��f�x�,����]D:$�Bg>�1�j:L @�i1�$�TOT�!��,�a��|�b�m�B���/��8�!	R<WL1�MD���^����U.wS�g����(泗��c2X6(����u_lhғY�@��9�?O!(泑�[Ou�LD.$�2R6b���)泋H��Z��X�ITL1�=D#���}��|��مs���\��b>�1!�����ȅ�X4��|�y)p�/!����i�m�CP�-�s��ȅ�Z����f��yM263��s"8�,���R�l'lK�k�"�!�=&i#��mW%���;0!��������/i�c?K9Kr��v�.�p�'!�N���m��W+�.>' ��3�w噙ȅw   @4YA2/E�-VVVL���	������y �e�|>�K��(}�Z�1:4HFe��ԓ�W̭���m�;;?*r�?JF27��x��l�|~�Y�p��G�RYv:�]��|�d
uNEg!�e�ذx���@��9�eu��B�_� z4$F:�2֢�g��3Ig�l�L]��漗�Z8f:��	���Hws��|��|c�"��y���9Sp������n�{��u]�����Iu�j�d&o&j���q�/֎�rl��h��Z��(泋h��Z����5�ʙJAt�̚p�h���>�Bj��D�P�/�K疃�!�,�,��3��B�I�=E�vʶ�����"�ϯ?�J���d	�(8�����5�1?;�O���k5}UZ[������r�E�u\�ԭTA�D3��B#��{�#Bj������e4E3��i���sr2�TNd���2晓?��     �KNN�	����y`��hX����������Y3���c������uj���WUUIZkB�-�bԸgN�����ku?AJG�צ��?'8S�w����|�D�vNmih����邪+�W��%f!U�]m��/�/�c�EK��9��zl�b>�b��,���i�n[�����P1M��h�f7罴��F����(Zݜ�c�A��Bw� :�N��D�D������R�M�!ݡ�|��E��7t��0�}�m�x�����=Z���L�u�Y�|F��͍�h�C�e�r@|�>���D�Tє���^��b��C�E����d����Q���R�;�-w���Ş��`_�$��E+�t�ֆV��sIrWs�g����\~��4�h��Zt~�a��گI�f� �L��[���R�p�O��;OuF��a�_���i�Ev!u�oK~��c�'���d&�~��oS~;��_�n
    �`4����Ȍ�hH���	���c��h��G�����3vKJJ�ӧO�k^�9v� :b2(F=?�%��x^~��	�V��[��_��:�B���|�XlivYHeѰ:�E��RY&K&M��|��n�{i�����t���~�����X�+����jAdE���^�EOԻ9��t���[2O1_D����w�pJ�b��v7��P�Z�g�9� �Ԣ�|��jjDV��9��/f~I1_��)��2||���E�X�TD?��B1_�������!����.s�*�-D�4D�.ܙni�o��ݗ%��4����7�o��2`�����R�.DP�H�){��ZL#��N��um��C�6]��	$��Y{��Zh�=z��:�!��D��BH�7ZQ�  ��IDATdbc^~����u?�=V yO�gdt}V     ����(yyyf���������������IOO����ʫ_�j����>�uFA�Ũ�����*��y,4b�^@�þ�ȤgApx�l���N1_�إ��~���r�e��d�ORݪ�%+.���X(�<�ts��t�k�.�:)��;��pC�R�j�l�NN�����9�E1_�٩��^]'�L�@��"C��w>�?#vC1_�٭Pg7��"+��۵��u��)�1���)��ts�k'����dlf�ώ!������A��9��BH-�E�	�	���Bj��5�ފ�
Ad��"���Z�\k&�L�Y%�_F����Ե�*$Ƣ� �/#G�wk�BjY�Y0k.�\�6�Yc�|޼��j�����G�yU2=���c��F8�7Y4)�'z�nv�_��m�D�CH���|�|b�����' b��ǿ!ߚ��}    ����f����]�b������b��?�N����g�5����DVL��~��ݟ�?���R��' b�Gǿ.��w	�N1_�-�ͮ�v��[��.v�םRY(��us�K�W:�E�v�47�{!�Hو�R|rz�@�p������X(�;vs���%��b�b�p�_��9�>ݜ���/r�c��/2��kBH3�{Cr!wA�ϴKS_A�af�n�{��t^�,O� |4�Ou�Bj��/2�r�|XF���]Q�9v!��W����jA�]U]2]4-v���v��t�UI�'	�g%sEn��;��e�P�/���/��2��]���r���p"`.N�k���ZZ�JWp~���2�LHL�=CH-4�;?6.��]�`�4]��;���4A��9��I>4�59�u\���
��t{iP�v�Y    �Szz�����n�z�;�1V��5� ��'@�{����@^��W
"'��bԲw]~���������&���.wZ��##\@S��pS�|L�,�',��P�^NXHe�b��ڶ�a1,�9;wsދ�|᧡Z��u@����q�OԎ�R�&=U=2Ul�n�{Q�~v��W�w���UBO�g7�L1_�=M�(��ŜE�S{G��b��rB�e>{�t~��/|���y?��&T,ۓ-=�W�{��3�N��T�P� <4�t�dT�b��sBH�e�l�́NN���	!=�a�[ٝ�-�-r��$�Y�N!��~[�(�/����H�!u�7$Ʋ����$�p�ԁ�ݓ����/赆�U�ȅ�BH-4�	���c2X怵�9O�fᄑ��v�����Q�5��$���;��    �L���RXXh�K�x<����3VWWM��>������M��3�<#���/��Ћ��4�+��=��w��87�2�6#������2����bK��B�I�,�.�jij���q�������	ݜ�Cg���H�0�q���j�x����b�漗�Yݝ)�-'ts�K��	������,���X6�(�'��Z(�B�pS���c�b�ξ ��<��2����y?��R�zN
!�hX�v�6�|a��R�|�c���;#��2R6"���=-3�<�_�:h~�E��nȵ�k��e~JK9Kr���8I��n�'��l�L:N
!��F8�7M eb�Aop��z�$z/�F8��R�p�C�=i�m��4�	��s��!1!�Q��o����d%s=���M�����k    �\.�ee���\[[���%Y^^��md��>֡A3@,������O���FAd��*�o̵K�H�������-l���c�^�-8�|��n�{i1_CB��S�ڽJ靴��B1_�9���~t���K���+8�ʹM�.��b>]�0� d����9�a1󅖓�9�E1_h����9gؿ��^�V ���iǅ�Z(�-�_�6�:*�ԢAh��r�����n����/�6S7���ّ�K��B,�W�S�#S�	��P�z:��Bz'/7�D�h-AR!`Bbj��b�sBb,z_����r��y	*���9i?�RKoe�ٟ˧�G��R��i��pBé!�m���Bw���Bj�N�T�x�8�pBˉ!�N1�>+���1yW�%%�{j��y>�����s�D    �'33ӌ����oz�^YYY12���j�>�Bet1�}}}2;;+��ł�����������& ���ے_����l��a�i�o�/E�h�����Y�)g�H�,�|G��T��B�iݜ�s��-��B`ݵ.7�n8z!�L��)T�����:Nu�\��Bb,����Y�u]�����sb7�(���YwS�2�ĩ(��{���焳�9�E1_h��g��Z�����U�t^�D��O��̉ݜ���|�C�R������R=�;���)�;s[.�\N�96<*=6t�t�Lތ8�|���R�d���|R7T���L��[�:�SiPq˹s�2m���Q���JGM�8Y_E�l'nK�T����񵥩ő!�ᄎ�-u��dm�ۤ~�^J�Kh�sN!��'t���T���6�'4t.���>m�ayO�g�W���c��i���}Nn-9{�0     r���%??ߌ����k����	�q��f�c�n��|��ݻw嵯}� ����_~I��
�r]�'���{=���Ug߀v-6�[�x	�yN��WoU�YT1]!8���M�z�E�NG1�9���~Lg��sR�Lg�GaBbnH,���Z�w���|���ݜ|k�`4}���P��(4,���3�9�E1�јn��7e=�yݜ�����u\�ԭT���J���%mK�d��𶓷M���CH-��χ�v���Q9���^';�>�^J�(�{�Bjqg��N�:�?"=o�8����L1_�%�]���Q,e/��5�`�`���������UwKV\�������|�\k�&����Bo���Z�ˆ͵Փ�'�gBH��Bj����J���d�96�Ε2�|�Bj��_>�';e&��!��M,��:�s�mR�Q,o�|� p��ƞ�����59    �=h�LAA�/��������������|aaA66��8�344$�����|��u}B�s��R�yL 8��=}g�[[I[�|��b�C���T���~� ��|�c&6ވ��T��M�tsޫ��M��d�b��X�X��ck!�;�-��ަ��b���~t�-�|�����:%�P��h�I~��pӜw�
�K\?w�b�Gݜ�>>l���Vʖ���BH�E��ֵ�do�ݮ8�X��WWu�	J+�-\,��X��;�|���w��H�.:g����b)��2S0cB���#���ބ�.�B����p�G��p	NC}�9D,9>"�d���Y�al�l� �X�_����R����ۜ7T���0bq~i�υ�t]a~y&��d����F��F8�&�BH��#��Jij����� p����LP     ��r��(+������,--�����l=֡A3@�LMM��瓤���;��"��\y��m�ot>%��R��# ���ǿ%�0�,�,S��x�,�H�J<��$�������H;�颠ʩJ���y���5�RY��O[>���$�b�=��S���Y�Y�X�8ڙ�x�X�򖳖�N��EZ�����|�yI���/�L7�3�d͵&�H��.�^��5���o���y/��´��:��@tn�ߌ�n�{Y�|W:���M���*�Bj�b�@R@NL��<����X
!���NV5�����s}�E�p9x������V3W͜"i1��i)�|/O�m��̼<Y�|y�y���Ŝ��r��L�4Fz&���M�H���`:�l�o�+=W�9�����!������S�$���r�R��y���5V#����MX�A��藩��
!��W��cC�a��!17�nJ,�����V��}��� �~�]sc+�Ԣ�pt>AX���~�^[!�N����9)Jϑ��5�n/��|�y)    ��222�x� ��++++���(���j�>֯i�s^��Ĭ��IN��k�����o.����M�����\x��d	 {���-����
�C���`P�ǆ� 6�7������Ov�~ +�+���@�9��H8���9�֥o	`�b�_�ђQ3 ��ι��z+{� 4,���_�>-��|��|��7А���V�D��i��t] 5P9`�������<�)��y>�����w��,M9�v׽2.���1��    �����%??ߌ��Ë5�cyy�Ƹ��>��_X���	�����Q������)�I� ����yo�gM�                Vm��MX̻ϽEj���=�M˯u��x|�    @�JJJ�	�y)�G�X]]���������!�1� 6�A1jxmڄ��Ϧ����t`/��w�{�>CH               �oC�{Ǉ�νU�2���Lx��u|HV�     ޹\.3���=�z�;�1���d��t��@�:r�0�>(F�Nɯw~D���fIOJ ���Ҁ�n�ߋ/�                ^,o�˯�P~��OK��H ��̦[����,n�
     xy��ɒ��oFMM��wɬ�����	��P������Zs`7�b��syT~��c�o���Z�h���o_��~�                �F�(���!y���JIZ� ����e����1a1      4v���������N�����:���dkkK�xB"�.����������� ,����!��Ώʆ�7e               į�M����'��M?%%i� :4�mOʽ�E     ����$���f�����k<�	�Y]]���e$c��,,,��Ɔ ��4�=n,��o���V�ŕ�& "�e�O~�����                �Mz�����Hyz� �,�yG��2EH     ��r��x)^�WVVVv�c4HF�[_��@@ � (fm�a�ն'�w��,��.�z�]]����W                �7��_������ ՙ� 2F�g����e     Δ��,���f����|��_�����KFF��5>�O�~�lnn��ښ	�� ��m��A1/�wuB�k����7KnJ� �gg���~Z|�$              ���V���F~������
^�kS���?$���     b�ì�������B���0�2��鲽�-�G���eiiɄ�蘛����-"����X�2���nz�������T������@�               ��V��o���jz�4fW	���X�_�xJ�|     ���5cIMM���"3TBB�$%%Ibb�x����h���������"@��2�<s�_�5u��r<�@ ��'ƿ)O�<MH               p \�?�?,���'�r�iZ-�}�;ݟ���    ��c�И��,3��ʤ��фɨ��M����۽&��5�Ff��"(� &=���_��?)M9'��g�>࣪����{$��&M�M������Dľ�UWwuWײ�������
� "�TtA��&@$��>ɼ��?�H�B&	�7��r�̝�D'w�������ޅ�"a�                �/�0_�m���Z����@�����zy��r�
     PLL����W�V�J\����Wa!�G�=�bܔ���#����vWiH��p�����>GkRv
               @ř7����I��/����Ԙ/l}p`�f�-      P�����"���s��$��C���3��-3�;+A                N��������ڏ���� T������kI�F      ���
2�hS�N�K�=mG���G ܳ?��:SG���               P9�'mQb^���t�����{2�9zr�ڜ+  �������
]&�-   �P�)����r�g��\�P�@(�j��c�\��	               @�ڞq@l|KOt�^͂��lqىzb���q  ��5Mk����+t���p   �bN�O)�t�7�X�k�*�� ���r��C+���o�:�               ��8���{��G��R�:@�V%o׿v�SVa�      ���P�i2�����G�������d;����y�!y�                �y9�y���9�"��nmu�|���E�"������)*      P����.��߮O�-��js�|�|���d�߶�RBn�                T�����d%��sƩ����]zA����֥�      PS��D�(6;Q�0N��������Q/�Z���               ��Mi�u��7����!����ծ�x=�m���
     ��	WJJ� w��d[�cu��7�P�1��F��$�0_�ٻH���                �K�O����-�/Ѩ�}���%�l�r�4?a��ٿXEN     TG����b�6B1g�#?C�n��+�Ӕ�����Ì�o��c��ڟ}T                ��|�S���R������c�&��K-��;?՚��     �΂������b���?j]����5j�@@md^�^�7�~-��P                ���S��u���vW�_�s�VkSv����R�)     ��.  @��Ŝa�YGu���hJ�5�a_yyy	�-̇��o秊I�%                �_ZA�����.j�Mw��\�>�j�|�S��[�	��NQ     �چPL04��g�~N٣߷�Bu�C�t˓��ݟ)Ù#                5˷G�kWf�n�ڄ4P���J�s;�*.;Q      @mE(�
�v�Э?���[^�z���K@M�R����|iC1                j�ج��w�ը�nj1L�>�j����9�B�,��U(      �6#S�2��zi�gZ��Q����AQj�˥�{ݾ�w�2�9               P���4?�G�cT��{���j��鱚�k��$	      8��Mi�u׺�uC�!�d�|��TW	����3�O�+                ���f��-�5�~W���R�����N|����Ykw�
      �-�xP~Q��ٿX˓����T������P\�Yq�+��               ���7�=�^�R��wm.���T7˒6������)      �lC(�ؕ��׽�a�ꖖ�(�/D���Kݣ7�-Rl�Q               8{$�g�m��-���h5B-C�9I��w�~J�%      �lE(��p�������t��j�_~�<=�z�r������&e�   J��u
���|k��$�           @M�>u�~��u]Ҡ�&��:�����qK�y�j��      ��(�T3��\����>��njy�FuP2�9�sp���ANW�   ��>�=��M�           ��L�c��-KڢqM/И&����G��f�k���:�����      �PL�u(7Y�l�H��ӭ�.U��hg���|����D�N><               p2�cJ�S��7趖��gݶΔ5);��ޯt 'I       ��PL5�S�.Ť��Q�tS���$(R@ep�Y��U��.V|�C                P�ج�����\7��P��PY�d�i���1m�       ��PL`�˓�ب�	�Ln1\���	8Ł���� uu                �`kz����=uo��ZӹuZ
8U��4#�Z��W       JG(�)����]C꟫�U�����r��&e�f�~�=Y�                �kKz���G����}h�ڞqP�|�U�      P>B15��U�o��ײ��uq���|5�'�$��"-Kڬ���^1                ΀u�{�~�^��w��i2@��[(�ƴ}���J���)       �#S�廜�"a��L�I}�����
;`��뛣?듃?�h^�                �Lr�\Z��ݎ�!�tU��5$�\�xyp�Y�ةY�i{�      �8B1����t�c��B�����0�,�R�i�A��W)ә#  ����v���M�-L^���            ��;+A����ޏ���j�_���@��cv��$q�>9�R�r�      ����eve���?8�DW4�a�]�$�~�2苄5�>q���B  xRN�:�=�\E           @����=53v�F6�{�a`]����qhё-:�Lg�       �>B1���@�|��־oԯ�9ٰ���i-///��0�/Kڬ/�hO�a               @u����G�i�����Z�女Q����'�EN�r����1Z��W.�K       *��Z�|Ⱥ<i�M#uI���AE��5׮�x[U����                jױ�u�{�x}�B��э��eH��:����G���#?+� K       �B1g�C��zg�b͈���E�����w�v�k��9IZ��Y�&�W|�C                P�e:s��p�Y��a�ua��� �������/%?S+����n�8        g�����U�I[�0���50��.�� �1��ѼT��خe�[�%=V                P۸\.mN���=_�cX3���Q�*�/D�>2�9Z�ة�I����~?      @�!s��/*�*�;^���GuР�.��F�^>B�;����ɛ�}�f�ʌ                �-�\Ev'�f���k�m��ƽ_d��
U��a~Hަe���>m�
�=G       <�P��*�շG����N���=���GvT��(��0�o�<���;�.u�vg%�">                �͜�B�I�i��no�	i���α�mH#yyy	gF\v�V9�k]�^mJ�o�       �G(%�+*��3�ٿX��{D��z��m���K�t�M������Mݭlg�                 %+riWf�3㖨�_�Ϋ�R��uP�z��$��tg�6��۸�v�Pr~�       T?�>����%���c#��O�Ú�Kxu
k�����(��u�'6;Q[�b�%#N[��l(                pj�
��<i��^�j�@��6�����؈Jw4/U���5�l���YG��      �zN�S��Š��
�)m��ױ����T��:�5WǰfjXW^^^:��iwf�0̶c���\  �j����I�&j�\M�4Uh@�|���c�]�S����tJ;���x�Oٯ¢B�f0���Md5�h� � ��ٹ��ed�@��IڣC��r��
           @mW�*��;$������������)�������Gg#��P����(�֌8�I�K      ����l�"��f�����ڱ0�'{�� �Ip�څ6V�h�����MT�?T��#?C�2��=v��r��HI  �
������jH�!�Ӭ��5�&�/���Ӷ��s F��.Ӓ�Kt0�����v�V]w=���;󕖛fGjN�����7y�bSbu&<4�!E�D�8��w�#q��B���{�Xl=PZPx�{{{2�ӊ}+�����O�'y�            pv8����&��ў���V���۷�mݏ6��U;I5۸o�n�s�:jG���R     TW�E(g�)���kQ���C���u� 0�À_�����1��H^����pn��Ä<���ˋ
  ��g6��v��<�N��0BA~A�|]��ָ����E.�K?�Y�n�T3bf�@�J�ݣ:����ʖ��nc(���Fo�X�3W�����v��lS�Yߙ����������R�f�O�:���e/��#��Uq����W5{�l
            g�BW��mܗk����|��2��ݦݎ s�ǎG���K�+"St�~$�g�Hn��m�S�?6b��(ә+      �,����E(U*)?ݎ����xL���+�7�~�^��a��_N�������K7���/�z~�/a�g����������,9�3����r�  @�1���z��'չa�3r�&BӳiO;�z���_����Y��*<0\�w�܎����n��g�{F�6��1��Ğ��%O�E��z��[��㉋�У��Q            ���6�����[�^>vǨ�#��p������m�Ͷ����c���������ۭu��������3
����:v��m�������Yv'��yi�r      �=�����P��wq���������z���"���"�\.eRD  �:6��Ƽ�!m�T�:}�}tY���X�o���a����3s��wo�:/-�Q�y�	L�qo�v�����j�9����O�PBz�            ��2A�C��vT�����}�� o_��R������e��       N	��
��Lg�=^|  ��cr��z������pA����z��7t׼�T��z�������k��������lX�a�h�G����u��<Z������c�*v�            ��R�*��6�      ��A(   @�e��3�����{*t���tmHؠ����K�SF^��yv.�/PQ!QjZ��ZG�V��]����zyyix��I����n�N�_���UG7��Qo�{��m�q4�V�[��;��S��5�yl^��:��Z^����r��qxc-�s�ƿ?^�,                    ��    Ւ������&�����1b4w�\}��sm?����~>~�ٴ�.l{��>�juo�]����/�m/O��"�"t^��4�� �b(�6:W3����߹\.�K��=o�;�ޱ�wYLfF����m��)�~��O�f}4���
�,u� � ͹q���~�[�                    �@(   @��ҕ/��1a�g�}F��V��z

�*v�����P���p�&���ЀPU���jڪi����\��b=<�a�)�Ȏ#uc�5=f�����]dc@�EbL ��E��P�!��ۄd�k�-���y�?5�ۄR���񷱘��֚�5j3��֢nPrd;t0�}/,�yo1���<߆�2�2���:��4O�7�WZn�P�� ����j`��j�F�"��9���M���u�h��/W7���7T�_�]&>=^�E�                 �g�   P��?�~�u�]e.c�!S�L��;���uo?�]wz���1=2��s�=6�P����f����/(�7����6�o��n����i�#[k�����.�KM�⦏n�'?9�uť��ڙ���m_j����T�r�y�d�'�=��gP��	���/�[W�w��5�vyOؔ�I�w.�g[>ӏ�?�e��z{��'E�L8�YD3��<Z��\���}���Em9�E�3�~˼���6���z7�}Ҽy���/}ZZ�'���k
�Օ]�ԥ.�sM�4=�2�}���yk�[�j�W              ��쐼*v�z��   �   P�to�]���e.�|�r]=�j�<z�nGJN���a���U�>�u��0Bՙ���y<�L�c�%1_�{�X��$o/o͸v�"�#K]&13Q#���1��ޙkg*��ϧ|n�%1�Ѵk�i�;���zM�!�z�%�q���_=����O�I��v+:4��'�L��־��>����7W�)�c?��H�Z�Sӈ�v����g>\��?���S�(���������n�`�`���ϱO���_-߻\��֔>SU����ꕫ^ѝ��T��V���Z��1c鞥�q֍:�z@              �b���"5  ��|||�t:���,�á���FQߵ���    �6L��D�|�J]f��%��(e�gU�m�M��ȷFjr��z�ʗT���8W�^�o=0��R��u��C1w���P�|vA�}�+3S�82�𖅥��Fu�	�&h���jt�n�:��`/&���v�p�a���\���Qm+���Sj=Ȏ�4k�+�\i��#[u�����o��	��#>��<h<�V?��}���˜��;Wh�!m�h�����~s���g�Y�ھ�                �V���6cFaa���󕓓���,����0̑#G�q��%�2�   Pm���vuiإ��]I�4f��*���ڻ?�k�����ϩ:{�����~�*, ��y����QaQ�<�nP]=}��e.s����c}��@�>��^���R�y~��y�r���+�yv䳺���
�PMЩA'-�}�>�����ߕ������լN3�)(,�χ~��Û=�>�)���߲��G4��s
r��=,�y���15��DՉ	M�bj��v둅�ؐ                 5I@@�BBB���`(;;[������PZZ������A�"   �Z՟����yg�S�̸F�9��G����Ru����y��iR�I%Λ�L��m����"�"J���~�f��y�o��+_��.����K�71.zqy�1����ײ�-�9��&2�3Jc��^]���.������Чy��ϼ'y{y�6i�V������I=��                �:���1���@��������UVV��<xP111�`P��   P-L�=Y��:o��7��

T�}��RC1���'B1&t���:����?{�Jn��`����j����W�2}؆*L��j��W�^jQ�������3�2l8eJ�)56㎨�(���jr�ɚ��D-ۻL��������0��.�[�4����U'����srV��d���۵��z��                �ʖ��c�/fdff*##CyyyJHH���q��    �Z���m�Ι0�߿����M	�ʜoR��<a\�q
/u��/و@U1a��b�ӭ}o-q�qxc��0B�o�\@Uh�\S�N�=nP����/����kҬI��~�j� � ͙8G�w�\g���u���=���oi��5"�                �~�1#55��`�HJJR~>;6E�A(   ���m�W]v)u�|iܑ�ܓ��T�|��<��7�:�_��WV�����e��-}n���W��7���Pθ��=w�s���������u�\.{X�k�$��Z{p������������Y�f�������uq��=��]I��cڢn�
]μf*�z��@�@]r�%vH=��?�_�l�D                ��[aa���ӕ��i�C0��OKKSQQ����    7�Ө2����=�}&�P??U���hh9���/�~���xU�mG�i����zP��&X����g�9����[�T��6U�^���|���Y��m�q^�����]�e����+q����0��u�|���%s�f\;C���Z�e�j*�xͺa�G"1?��A�/}^���>az�˛X��{�ײ��l���Q�+�?DU�YD3ͽq�^^�~���*r�=                �VN�S6�b�/&cFq�Da�w��P   �j�N��:���VmL�(��^p�2�==1Q��o�X�2gÜRC1&c�����<���ܹD��yd���{9�6�aDE��WhR�I6Sҿٛ�ܬ�������_=�W�zE�v���u,ݳT���:�ѹ�}{Md壉�����̣����������_���c���j�=��̵�s̹ctU��*m��[�s��w_�2��v�w�~g�3�-m��[Iv&�Ԍ�34k�,�M�k��~�L^`���=�c#5��                j���~111��1Üg�� �#   ����U�F]K��v׷B�4
+;:a�UmX�a���_�Sn[(��m��텄bpZ�F�U�f}�>����y�Y�{��J��ħ�ku�juj�Im"�ظJY���){��⧕����1��hQ��n�}�u��˯M�b��o��=�{4���m��}ſ�0��I�߳iO5y�������|�N����8�o=<�aM�h�b����cnn������L��q����͸vF��&��ܒ��̷��P���������s9����������N��H$�P�!m?�]u��G��,w�����+�?؞����mG�i������                �sL�8�R�)>m�0���Py�    �nM���˫�����
3�Հ2��PU�ޤ{�s6�@���s�����jZ�i��=�V^� go/oM�5I~@]v���6o����;}����Թag���|�k�Ͼ7����˘X����Z�e���bSb��7O��_������N`;g���a�1f����;��?�%�\r�u�(���O|�B͛4��8���%�f�a����?���A/�xI�bn���h`���u=G3��~h��L ��yw���o�ߟ�Z:i�3}��Zw��Z���C��H����\��v'�>�:�E4����I�I�Q�c��?�Yi�i6~4󺙪l&4T��d�'z�gl8                P�
m�%--M���6�b��6�f����Q-�R5F(   �G�1�ǯ*fD�e�o>�YU���_�t*u�����i?���PL���TDdp�>��������	h<��Q
1�Օ�ڹ���5��H��8RC�����=��ן�)�����?e/����m�&!#A����\rv�.{�2�y��GN���ﳱU���kj/���k��u���m{{��)�os��|Q}��є9S���SU2���RC8�Z�w��.��y7�;i��t��~�V�_iO{�1��_�f�7�n�u�9��5qkԢn��w���O
����Σ~����rۗZ�m�VŭRaщ�_��R}t�G��u}�k������ݯ�x]                 �9�N�1���L���� ���8�)**����`�^^^պ~D(   �G��l[�\V~�bSb��o�_�Z*u~o�^�J�굲���l=�U����]���B�l�����[A~AZ|��r#X�S�c_��|y{y��dh@h�����?i���Z�}�	��L�i���S����6^�u���E�b�?��ɚ3݆_�EΓ�1�?/��6&l��	���M	�l��X|z���>T����������;�^%f%�˞;!6S&�0���L���tUs_>��q��Ky>��&̜Pb�k�c���1�3���~zOw��=��m0��b�-�O���^o��F��3���;4w�\}��m;���e�7֬�g���/�WZN���O��z
���2���Ƽf�ӴU�                �Enn���������Ogee	�>>>
	9��T�b    ��"��:g"1�K�pO�o��^1��e�����Zӈ�e��s쓧�J�U漹�b���^��J�Ę���ݬU��t4��I�u��MT�k�O}��U���6��-Y1�߆b~-)+I��|�w-ݳ��e>Z���d�G?�mso;)H����U�]uR,�8���留�i����n����]<��3��y���8׆ON�y�n���	�?��]R$��c_=f�2�����[�\��HHOp��6�����ֲ�1��8�<��2���q��0A.*���u�Ѥ��y�?էy���|�F�Jz�                �6���QJJ�233���n�/�v U�Q�F6SK�T��   �QM�4)u�|��1��wƿS��g��PU+�96RsR�i���~�5��T�7(�	^�s�=�r]���������֒�N)9)�9c�++_��5o��;]n�&������)&(���66�R��X̷w|�-��~�z��7lx�ّϞ�m0�/�|�K�]��l�	��Xs&�9�H�	��8�F�1�R�ϙ�ʅo\Xj��D������q��Ӂ���̳��,��ۍ	ݺ���m"ۨw�ާ};L0��A����	             Ps���m�  ��\.��������94!�_a�N���E�B�    ��L�4���(_ۨ��q��oѿ������\��V7�n��i�i򴣙G˜�\�} 1��,{NTv~��w��p�<���j�A~A�)ȑ'��)fb1WO�Z1�����ݟ�=a�������CC:��0��@�;�]M�9��ǰ":5褹��*�7മg����q�/�?~ފ}+�:n�z6�q�;!�SOFb�%��He�gU���M�������*嶌�4�P             ��ٙ����U��G�z{����Bw p�),,Tvv�����& �p8�y�xAA����[�nB�    ��}K��-ȭ�u��J˺-+�b�(5'U�b�	Z�=o��s���ۧ��
t����	e=�FuŔ����`����J�����n�~�`�.��H��g֕�]�<g��:i��_�Q������2�q'�2��8�;�Άg*���͟<_aan-o"0�>�'����v�z{�I�A��u���%���&8�H��Σm謼�aѲ^K��d�e              ��6^��H7|x��)]urc����7�m� ��e"/&����f�9^<�i��읢�вeKEGGU�P    �
�*u.�0�R�uK�[�ǡ�����`-ۻL�ebω�j@���z��@�M������苇���fyBYϱ���N��D���/s��@���ˌ#*=/���˴��`�`5�h��T��)u�|�}�Ƿ�y���z�	s�.�p�FtQ�:��6�oТ�N����ɬ�g�]T;��7��fߤŷ/>����D]��eJ�I)�r��ɚ�i�j+�8^����<����������a��P��]X�o�P             ��жC�����q���j�W��9�XGӮ�fwg����  ��N��������p� �9n�3Ü&���l�?|�p���   �j�udk;΄�A/.Q��R�hU$xTg&�Rٙ�Sp_�3Oc����A��?��_��o�۾��V˼o/o}x���5���$�9����%O�@�;Lf����vd����������^���{u�2Q$��(���}L��"1             p���h-��P/�|Y��vgv�лYo;a��v �ʔ��ic/iiiv��ŧ�a^^��$�����&M�U�P    ��)�QDPD�s>©s9���G����=z;rr˜7{H�I�'��9o^�@yv'�.s>�/X�'L��W��p_rv����xϏ�
�ҡ�Cڑ���]��Zu�*��jW�u��5o�{K�q�)��6�?��[˚�͕�]i#1��{��=o��4k�~��Q���/}Z]v)u�H���             p2���{/�W�w�u\g�ǫ�u?w�s���  �f�����8)����N'��eiݺ��.T-B1    <*�YzD��xJ�&n��w��\��R�sl�P������9O(�X�e���k�O��_�Z�/�bL����ҷ����g?ߑ�Ш�G�XLi�bC�ѭ}oմU�*�~�Gi����qk���ަ��p���sl(�ϋ�l���L������̊}+             (۠փ�����i�M�rۗg|}f'qfg{#;�  U���P�����̴�)))6 �p8�qs�Y���ر�ƌ#ooo�j�   �Q)9)ju�$�!т�

��������CS6��s\����Z�����`��ɺC�ԽI�2�{|��6tr ��P1&2��qZ���(ώ�v�&_L�B�^e�h�D�p�BL;X�u?2�ui�ŭe_��͈�q�y��̹Eo�y[�8�yu̫�>�Dx             �=&���͟��/��R~a�Y��6�����qxc P���󕖖f�/���)>4������6����СCu�y����K�z�b    xԡ�C�ѤG�s�V��ĭѴU��^~\�q��Pu���.G�C�oV���t�'��]eϫn��c�\W�V�k��� {e�+z{\�!�ЀP�0�]3���>��Y��/ھH�Z�/�q�˼��S�2�]��n��C�ztأn-�:n����O'�_�*"sn�w�z6�Y�2�)�o�/             �{�{��^�i�GfNPlJl�]��A�c=��\�{�,��\ �[999ǣ/��3�����UݺuU�^��͛7W��x�    u �@�s-교����r}e��i���zP��b^Z�^\�b�˥d�(57�F���Yi]��<�}t�2�˻@1�p��s��F�ic�F���e�_4��@����2�����=~��en]�#�����˥��?��'�7�n(P���$9��             ��>�>��qY_��ע��=�N7ts�찫qxc}p��fH��nJؤ�3� p�1����;233���q����Pn.!1�L

���q<c�����    ��I�K��V�z��'y�j;�ٛ�W����R�3�~ѿ$�v��unعԹ��G��v(�����u���Z�|P�А�4q�D��H��^�MnRh@h�˚�����o�m�׆e�q��{�߱_�\�zMR��F�.׵qWM�3Eo�~S             �_�Z7K����y�L5kP�ru���ӛ>մU���pf��S1��0���a�]����뎹w(� [ ����!3RSSmƌ��$�����gb0��Ѫ_����GaL&00P�y�    ��\�|�&�ϊPLmVPX��G���$&��i���.un}�z�:�ѹn/?��x�yџ�'Tj��W��+���\��}l ��=��kԿ�*`��K�\;S�\�^�zp��n/�̈g4g���	             ��ow}�^S{��>��V�\��~��W�^���2w
�[f�{��/zl�cvۯ�d�e����ۈ �f*,,Tzz�233�aq��p��iii***�3���Waaa��/����8��G��3
   ���Z/��U�������
5ۺC�J�ti�E���ɑ�'��j���K���`�1#��h�����ӄ��ܒ����uM�k4��2��ۥӂ-���0��?�&Jb�h��gbb�ۻ�|th�&����V�$             ��L;����c=Vn̥G�����ݎ�4�h�Y7�*w�=��h�� @�s:���Ȱ�1s��<s���T������3L�Da�����\��b    x��r����gӞ%�_|��B��ݮ�ts��K�3d�q�f��)O����eΛ���w��jY�e�/wE�+ŜE�"�n����k���S�r�v��#��/K�h�Cn���o��@G��yt�/3��8B1             P�¢B=���~�����(�Q�ˆ����?�;]3;S�.�.q9�-�;�߱;�,ϴU�t��{��� ��rrr���i�/�!�1�8�����(<<܆_L ��_��0QQQ���P�P    �3_�/-�.���[{p�Ps}��k���҂㺎�X(�J�������(O�&�N�r�Z�S��:�q�Rn�����7VlJ��v�7���o��w����(1ӭq7m;���l;�M��|E��B���3�*�Bf���ޤ�����             (ْ�K��n�q�]r�%e.;��D�=����k�������s�?�{�c��*�ٹ�ߪ�7|, @�0!���Kq��trr���vU���Waaa�_�����m�DaL�N�:����B1    <�-���Ꮧ:?��dB15\rv�V�[��m�8o�4�<���R��vum�U�[�/u~��E� n	�,w��1������h5kh��q8��TV(���@)9)����6���Ou0��V�}���w��AuK]�¶�(����'�o2������~�
��1�z^�g�v'�����̣vc�^������D���ƞ7*4 ����D$             �a����=<�a=3�Rwitj�Ik�[����gw�ֲ^K;a��6�[�z�ĭф��ϱO ��QXX�����/���r8����4���@�

������@e    ��L�|A�|Q�$��L�S����@���O������}�Ӄ�?X���Ae� �Y� w�8Ky�{��_<|�oKzn�f���F�l��U�V�p݇��i�2�2u6I�Jҿ��[O]�T���s�=�2g����C���Ly��Y��w|�����ˠփl��D��������J_OV~���>��Gu��ο���9r             ����K���q����؝ߕ��Xl�5�4��(i3��`�,E�"=��9��7g�S  �9������L������L���H ��������m��`L�8%g�    ��~��^�z�s�~��������N���n���WLUDPD��w�K/�xI�)�Ur{�kt���q}��q�q�f�7ܱ|��r�11��~xM��U�t�'w�C�zv�z��W���Om��N�w�/-�F�J{�1��z�����v�V�>�8���u6i�Z�{O�Ğ����G>�[T�m0��?.�G�ˬطB              ���
��������xg�5�C�b@Bpw���-P �-Z(�B��o[�@q� ���S,��	�A������/���$�����z�Րyff�;�3�y淜��yj�m+�}E����h��-6��""���A0�"!0���ɿ���D�����C��#�0Q?K�D	�A1DDDDDd��ÐC4S軖銀#8zd�$�a���*�GG;G�o4��42�k�Ib��M&���V���;~ǻ��@d�������c(���fY��-@�ɕ�g���Σ���(��F��]w����`���j��2��ɫ'*�jh���m�W߂��2_��]�v��W�Hv\�k'��zy��p��5q���<L%D/�������m���
Q�<x� ug�E��=1��(����j>:�ja+�zzDD��˗/U��������S�"��d<%��0OOO5D��H ���#���b������,��|�������Su��`����Q|\qu�,��=cѳBO�pJ�s|��ѹTg�84ä���*ߣB�
����a֡Y �		Z�z��6��:����G|�wm�M,����0��X����cꁩ������2 I�j�i[��
�)��
�+�<G�k��5-:�����3���!��`ܞq���H��� |W�;�m�=���i""""""""""""""""""����Wuy �zv;kʬO+4�����6��5Q�s��%�;waaa*�����>����I���?������D��A1DDDDDd6$��K�.(�����Sd��kQkF-U�N�G>��c���6O��Uo� A���Eo�>���ͻ7 ���V �z�g,��]���q��m���Na�ٵ�\�3~���K�WÑGT`L�@�x��DƖ�\�VE[i����<�=������?�������$I�UsTE�2]Up�����[L�7	öKР���*���5�3d�D��Şt>Wir%��w
n�nѶ���|���n%&
�j�*�����⟳��'0��8"kŠ"""""2R��6�-Bz� �]R�mJg.��]����&{�<�NC�"-Uѿ.�ٯj�
f7��+{����yj#�?�6ک�+O�TQLI�햴S�0G;G�m���B8F��� ��)��`�����O�^�;�e(��f`t�ј~p���擛��L�#�����0���<4Ӫz;���M�6�[�/r{����������8}�4R�\5���J8�;�m���*,8� DDDDDDDDDDDDDDDDDD7yR����K
�)�R��w�v��5Q�q�����ꤓȜ��������0���eppp QbĠ"""""2+R��wM_Lj2I����{߬�K�/1��Ib�B�����_�	l�ý���Sg�����f����e&I�Da�m0V��*�C]WtQl��sF����Go;Y'���һ�W���
	��@$�i\�q�������W�^z!�X ���S�O����_@.�\�m�)�
�+�w>��sx�A�d�Эl7�(���S��凗�om?������cf���rQ�s�6�[Q�H�c��LFr��O#�E�,�岔C���94""k���c�����\\\T�K�ԩ����!���666 �O1(�����������U!��h������UQ���~Ŗ[T�x\I��_?�2 �Se�Fhx(�/h�-]���F�����#f}5�7T�\�ղ�G�?���yj�m�2�%�i����(.Jf*ip[�)�5eV�-����ϑP��=��>���>�4��9�`뀶�ۢM�6���&��5;.�%����|�9�h�����ȍ#���:,Y�T�T�Q��?��/�����=c���k$$yh�?ah���gCڗ�X7��Ŝ���7�Υ:�z�C�>G�����bY#�]Y�|9Cb�$�zG�H LTLԿ���@D1à"""""2K߭������]�
Y+`S�M�p�V�Z��g���ͣ*��Pn�n���*�篏�y�"�sj�����������l� �"������}y7޼{�w�pQ9{et,�M��h��D�@�y�j�!���.(��l���p��_oG��5���S$��g�b�?�UP׏�T�a�RV�Ad�s��\�����Ҭ9�FoP�A�8��J�T�U�_o�O��r�j����an?���&�ܴ��b��A�\5U�L������Act�9m	��"���b��軦/^�}""kr��qܸqD�?vvv�_�`>���'"��EDDDDDf���w踴#�x��ڣ��3U���w�8w�B�C����<{�L����'C�T��͌��\|]w�S��m1W��h���G��-����s;��s������=s�t��H�ܠ��f�a��� ��9�:S%3���f����Hh�4j�(	���E��`��F�+����y;��p��6��.����R=�������3��X{f-,�����~>w0� z���`��>�ĪG��������������������(f�o�)�S����Hǌ�@�@�k1����۾[�n����4��;�ADd��ƽ{��(1rrr�$�����C ���Z
"���ْ/���돣7�b��T�.o	�T{�I������髧 㐛E����2�qIm{�Ψ����J���m�c7���� �/6���z�(����`�+�`ߵ}�Q����;������fbjө��S%�+�e W��[�cىe#�Q������%���퓰E�Q1���G�0p�@��i6�\��B�4�h爰�a��������?��H'�ӚNC�"-�m{��5�X�B=�%�̪���{bT�Q��m-���!�W0z���f����]�z�=�5�����>��DQ�vtt���ٓ ��0����['A^Æs0h� �
�$_����d��h��a�,S֫��z��� 2������}A��WFޑy���+X��P|\q����|�}�cH^��X�?T�öC�� ����Gcs��q���N�a5��q��:��G໵����{0G�N�R��Ib��=_�z��mK�?""""""""""""""""""�^��E�3YQ����J���㗏?�N��w<�T�fI�Esz'{'Lo6�U@������sY���D����...`���?�xzz���Dd�CDDDDD���+�;�.|r�`��p��T��ˌ|��'�c��q�֭���hN#l�k�_U �)H�������F[��p��{����l#7C�S�?軦/,��G��e'��Юz��}2^�IV�]�c7���?a�ٵ0WGo���Gn�9���O5~B�B�T���.ܿ�n+�aǥ�Q!1�
4�W����vߵ} """"""""""""""""""��o���SU��>�!�<s+�0Z�3��K`n���������.�%3�D��8q���,Qhh(�̝��Ӈ�$FBa�~��y'Y��E���f5��\��tC�����)���/���׃x,K�/��gw@�+�tV�Y�&�MЭl7T�^Yg�AL�{��/m��}�����9�ʂ��[�����]�7�\كU�W��\{t�gׇoA_�o8���2�H�"X�a�
�賺_?ss���XO+A+����#j�@�`kc����o_�������-��X3���m^�y��SA ��!�W>���.Z&��DDZ�!��u��m����:y�b��:�-=�4Na��H���O:�=x� �w�Y.WGWLo:�7���?��18�E�#ȳ�=����z#�`��6�gn�y0� ""s���%4[[[���}���@D֍A1DDDDDd��T���=*e���D$a�D�pwr7x>�_>���'�M	m�}e7�?�o��<+xv]ޥsܑG`n~����!�˩ۧL��������Ր�5h��v�g-�E0��On`�3]}z5C(�L=0�+�G�d)5�Hqj� jN���W��Ҭ8���oCЯR�/�I�e)�C=�m����7����/&ȴ� ���e�c��p�9��l#Ƕ�+����s�D�ΞX�q=<�{�m7y�d<{�D�8��ȉU�����Q���!w�ݵ��G;G� ÓWOT��O��UЯr?����=��b��%��GJx*�b����+��K�x��)������������X��#{��Ѷ8��+���6%�8J��t4��	��ʦ�V�c�k8N=�ii'���%x��޾}��`gg�!0���j�KH��M�:d&"�Ơ"""""�h��"���65DI��RdB&�Lp�w�KR������wx��)"�D���Oo���{��Z�_ܮK���b��[Oo�  ����M���7*A
�^E�R��^f` %	��}��W}�F���QaR��s�F
L�G	���|.����x	�iV���}�Α��L
Mڣ�Gꆴ���Lk.�l�ֱ�)��/�a�5}0/d��{-��7uބ\����{���8'u���}��!amrL%""2TTI\��G�C3r^+Z�2�wZou~(C����%��߾��%���c���`�!߱X:	�Hf�̠�����^�'s}D�L�Ó ���Z�@����Z���X�O��E3E�tEP$}�N�[^�9]��"߃�v =�9��K;���~�y�DDDDDDDDDdy�o�em����Ao;y��ە�b��9�^V��W���B����m����B�-�tDD����� 2y�G�`$F�_�a������%3�"J�CDDDDDVG^��ĭ �#��ʃ�2���{�·�/Je*����l�5�װȰ!7g��+��>�ѯR?���~2>�Cr5�S�N�q0]���%R�����O�_%�8	M
��6�
Y+h��t~:/�B�,�����E����7+�Qa1�B��Ս2/)J��=9��ܽs8|�0v_ލ;��(J���0����K�;#ǡ�On�ԝS�������?ypS�3�嬆J�+��%	T5��z$�P��=��W��b�e'�a⾉8}�4,�Q��j�Am�$�o�p��5ė?���e��V>�TCS��sy�evaLr\��9.��}B}y��Q��T)�y�x�D����J"U2�}���T�Z�H����
$�Y�n��F���t�T����WCkU��KT����'ADDDDDDDDD��@�ц��3�_|��w��yy�w��M�m�o1��hա��<r߷�����1~�xY[[[���~
�����b���������L�H��#�W��ފEZ״��mjͨ�#7���~��DЩ �m1yR���MF��h�n�v[�-���b#�w�"��#�D��ma��Fg)`�n�w�<+A�x�J���]63��\U�D�'�{�:/�H1��u�P�!,:�H�����u""�x"��;z��F�<������^��������ͻ7H��|��wcU�ml��u��ѥt�B�u�q��X3镩U�V�uۯ�<y�y�� "�u\J�^�k��S����ٌ��b˅-}n\���`ݨ@2�gBb&A/5s�D��T/���.�s�=��������GWADDDDDDDDD�/�H�z��؝�IG���Ò�K��#�f;���k�_CDD����C��#�0Q?�3*DD�Ơ""""""""���Z���NTq�>����vԝYW��TQtlQ��5}*��hR*S)�3v�X�<�������c?m\��ǟ��T�8k�~q;:.���PX�t������/ڶ����	��fU�̥�0�g8���ڞk�>�9������\sȦ!�A��V�_.k9���|L��M���v��賦��k�_�?ނb�=����	�mT��$W��hF�C��Zn�!F��Bu	rPe Zk��L%�|AB��[�
M""""""""""�$��=W���C3M��.���b��;Eu�@DDd�>�I�:5<<<T ���q:n "�	����*�(�ހ�(n�n��y�Ϯ�]�w�Rɍc�M8�T洘��;;����޾躢+�^�o����+�ӦvN���5eVus�'��f����u�cʁ)_(��=�
L��s��V�^�Wo_�N
������+ꇦ��⃋ ""2�L�0��<�,�����0�!��$a��TNW�}�w���I���~��˒�}"�>E��ή;1n�8u}���[�iJW��L})�gn�:0ޖ��>���h��*��Z������������ٻg�<�9N�9m�e={�L�ߕg*'7�l�2���b���...*F�_���?��xzz���DD�A1DDDDDDDD&"���9�3�wZ���b��m�d���C�1�1��t-�Ug�l��aK�-8��k����&]e2�I�icB�tzU��>���?v~�p��X��)2cG�j�0T�T�A�`ڂ8��|���K�5�����:�T�V�]����;�:�ӲNL�ſ����a$`�^�z "�$I����<s�M��RbӹTg��yX�����g��.Ȉx]��������%�N�""������!�E	��P�����/��`P����E��p�9��&������G����_�n�rYz�~q;f4���sti]�5j穭�b��)U�^9N�� S~.���W�2�l#��k~��#"�E�T�Qo޽��wҋ�lCQ���ث�y����]6������������I�\�	ep��]T8���T��\k�9��ȗ*��%�Һ��wodI���yv(�A�"8v�XX��[�5�����&[F�B͐�.)�Ⱥ��[�Z�C�-���/޼���'�yý���w3r�J�,�
�-��$�m�ѯ�.?���������������̗�?�z��<�`����s(�W)�^�w�,�DDD�bkkWWW�"0�
�*U*$M�g7��z0(���������D^EF߃��6��v]�����VYH���r���b��(����6�=0��|4/��v4I���V�^)���k,����:c��6��P�6H��E�v��Q�5�{x�$F���P�s�Θ�h��4�=fd��iH��>��R �GN��\�\��	�Y�z�
�1e�5Y������Ѷ��O��T�K����%�A�Ϛ2+�Z��j�����揝������aI޽��M�^݋�W����c5�}�s[߂�h_���9���S�?Xwv.>�k��95|r�`���&[��cQ�	���f����I��ʾ2�W>JW����W��R���N���k���vb��]j�^{���v ���|o������[��տADDDDDDDDD�G�'6hn�����^�z���'7��� ""2���\\\>	�I�:5<==���%�!"""""""2��U8�j���߼}��K�Ú{�����O,����!5��0
]���SߝRa1kϮ5�khX��*�v%ڡ���0�,)� �e�*��G
y$T���[�VR��2Jv�_��B�$I4۞�sd�'��ĺP�`ڂ�Q��*p����)����펿��DDDb�х���f��+���U�f����Vo۪9��cɎ� �9���a�$tGMV�^���ǿ�x������&�p�\�4�;�9��Z?�傖�To޽Q�%�<s}1ο��ɂb��ʆrY��w��iHS DdZ�^�sp��h�+�Ku��*~���_���(�=�����QF���/�+�`V�,���$�w婕j���f���U��|�7�w

�)dp���6f��~��$�H �Â�����ȁ�&[x6��H��H�DD����I�D#�0Q?�{���(�`P��09�{K��#�� �g���hV���6m��Q���uV=�Z+�ۆm��a1��<� OgO�n���O���W��ĕ��W�_��ӾD{���UXkm��ń����E�M������E�M�R�1��T�0�(���ŏ��O��Ӥ}����b��̭����1��4�{����,ˑGT(Ʉ,���R�wK����Z#�C��޾���[�ޗ�w�F����q � vtݡBM�4-�}]����۰T�.��>?����������}��E�u>����s�à"�p0������V���W�m�d)ѹtg��5?�?���`d������O�X�9�	�m�o�~q{��SZzb��mx{����Q��ךx7���ADDDDDDDDD��ĭ0W�����*�_j�����<_x�hW[WY:[[[�����	���P888����cPUR��������k����ňv%ک����Uo��l��M(�g�h�B�ȭ�R~[�[T�^E�JPE\H��Zˊ	)���O��#N�I�B�����G
���o�=W� 1Zc(��m���ۧr=���:����@���K�]Z״h\��*:'""���������8�� 2�Ȭ����-��Ĝ�s`�$��TB�CQ}Zu��wJ� �bgc_o_L�7�j��^s��N�N�o3���_�_��W�Z��7 "�"�W�Z{�ك�95�IH�bL�U�+캼�C0��]����������6���⃋�3����o�9�i��T��b���������(F$��ڸwGDdjvv,�7���Ӈ ��`�g�h�&""�xD""""""""2!	E����+G۶n޺��u�Ϯ�{�����zz��Tƴ��жx[�v���ǡ^�0h� ��{<����/+�sjLh4�ҽlwU����XM_){%�o9��3�m'�g�4TE��N��'5��.���~������(��G���
��؛A1DDd<w��A㹍���~8�9j��+�g�A1�v��U��:���]�M՜U-:(F��}���|��_��@c�?V�$p$ %2� Y9.uY�;���lS0mAbv��]�q=�*S������uδ���X}�f��wN��u߫���T�Y�N�x��1����������������#lll���{���`�wwwxyy���C�#""�aP��uZ�	�{F
�Ѷ-��$Bz�������_k���k�[�'o��Ⱥ#akc����m85rՀ�"��7x�X�f<�=���a����Q�R������I���C1��Ϳ5���{���X;	�Y�UrV�5;x66�� J8�_���Y*4IK�UADDdL�n���ѳ|O�6��U���+��z
����f�ڿ� ?]
�) K'-��b$�3�[�xr�h�j]�����|r;/�dP��P���vj^��w �2��+ū�/����;��z#�W^���{/9֮;�DDDDDDDDDDDD�D���������ogg��)S~�����-�0��� "����""""""""����bmǵHf�,���3bO�=賦��k���?q��i,n�Xo�N��u�+X��,�G���~���"�-�kZl�էU7�wp)Xh���m'�=�2#��0Y���l��X�z)һ�7���K;���o@	oҾIz�b<�{ K�,�������e��Q���b"��3W�;#b�����ЙSd��[vb�j���%����W�#w�4�r$��y��:�-:��޿Y��g��=͖2����]�_k��٦P�B�!"""""""""""��%K?~�����CLT ��a0�CDD�A1DDDDDDDD�@�U�̬�mW U�TѶ����M&�M	�x��l˅-(5��tX�<��h���z@�%���r�v.I]���"��W�R M��ug�ŕ�W4����.H��%��~�6�mt:�Nz��_�?~��Ytb͙5h��^�}Jxg���Uh���9M#7�X=�W>dI�E2�;��5�+""#�.w��������p����	M^��7E����\]�kvst��W��������w-��������9>L[P�3���N�Nx��9n>��sw��`�A�7�+9FNW���G:�tpN��K/޼@hx(��9�������0'�Z��z#{��*`K�o���e�Ku,���?8v�Z�̙l�r���ΞH�o߽Ž��p��URq���/W���B�4���%-�9$S���վ�ԝS�/Y/��8���Jj�)��0�b�H�.��bd�#�s�G�D��pU��[���q���6ZPL�<�5��Y s��3�:�ʚ*+R;�V��$����S=x�@c��;���ΛM�eT0�O$�P�%���r"��ze���X��U�Aʬ�;j[{����|��K���<��i�B����"Y
Y������aPY�ܹs[TP���-���>�HLT� ""�à"""""""�x���nW�zR�w�hQ�*e����:�kv��E��X�;�G�L�4�IA���K���?��U/��BA��+��_�
	����mUO�k��Z��t}$B��Cq���m1e2�1x����ۊn,�43�!븖n��<)X.��,�樊��+���J�l�]܆U�Waىe*X#������E�����-�}��޾��N�������ͱ�H�~���'A/���s\����u�Q+O-N����켴�LÚ�k��O'�$6hV��o�*9���k}��|�����:~'	�}��7>�}T@�!��ץ]Xxt!V�Za�0	=�_���qR�?~�x�㤈�[�nhT��:�3x�`���/~߽lwdJ�I�4c����gw����;�o��
}�
Y+�(;}�4�G{������`��:۝�u��-��eK�]Jw�?b�p��쾲[oPL&�L�G������s�l��l����m)�����~=�]�3(F�%$L����?�%�3��1���HHr\���:����f���r�2h����c�ŭ*�F�>b]�s��{�PP	��GΡv]ޅ�!�x,P��\��H�{��~��6�K���s���7�ux�?[x���$�N{ÂQ�\ȵ�.r}!��&�4�9N��~ݦ:B�G�X�� W""""""""""""k�'O�sagg�O�`��ԩS#U�T���Y�ţk�����қ����Pv}l:�	�LS�O��mW��9-R�;��@U����/��h�U`p��������)�tX��#跶�*��7��P�T�'��>�_����{�N�C�~�7F뿐B]@���/���0]��'S���P#W�h�=��p���al���w���B5L%�Cr��Vbj�9;;�PLR-A,R<;x6�N�h^)��Ā*t�;z��A1�i�1�w�
�1��%�D)���{��AB�B��M&"�gn����K�Ed�~q;z�ꉳw�">�qC��~��#
�+��e�����F>�W��j�b~)��Z�d�yP���'F���d]6�փ	�P:si���8�q��� t+�M�=��4���S�WL��9	����w:�IhTb��^�;ސ���V�!��7`I�\˘S�Flm8�Am�~�9�_�5(F�$�D	�H(r��c���y����O��2$ `Ķ*�L�LM��6����<�w�<@9'뵪�΀��$糝Ku��U�GF��1�^��$DN�S�Oa��*��������S�	R�k	]$�)>�bU���=<dY$|�髧����=�5�{�>>>X�xq�.���I��D#�0Q?G��2Y�Q�5��v��� 2Dhx(�>]Q��Ɍ�5
�޾R=*K���nSE������QV}��"F}j婅ýc����]�w�
�E��h�1�Ǡh��h��A�Ӝ�w>�}�8���'7���,(�� 2��פ�p�wT��rVӜ.��G���Wdn)��[�o�V�H���>?�cɎh���]�g�eH���fӑ9Ef��[�X��\�y1��	)$]t�·d{��m'���?�e���J!�c�A���t\�OG���+�Ŭ�Y0�\��0��tT�^�(�K�OD�bm�:��*�O���������#F�%A�Z�r�²6�P!k�X/w����p��_|N�%䘿�������:��"AQ�������.�	��"!��@��_��>ײHKX? NǬf�����y.:�	A�If4�����A�Y-СDt\�W]���(�B�WI�_leM�U|ʱ�ۊn�|��V1[E�w�$�N	�j���V���ў���Ix�>�_>����*��Y7%HƔ�M��`�ܵ4�'d�Ş�P_	�!"""""""""""�Vy��A���b�y�������C���sԿe<Q�����(ƶ]�""��ӷO�p�㳤̂�i�GP��L
7[.h�
ݺ�骷��,?���)\Vs�AmC���ά:*(1�B�Ca�� Zm����9u���$�O�w|ě�8Ϳ|��&	���L����v¼�yF���Oh4�6��T#j����4ʼ$�E�%�����0�����y��F����#f~5S����8���$T`N�9&	�(��$�<��ͱ��ćv%ک@�,b*.�>r^���dK�-N˕���#�U��ζJv0iPL�����9��q�g�e���H�Ǘجs�?���RNs��k�a-d���5�����V�ӎK;p��-�7	�Z�ne���Q%G��A��M���N�Ͽ�����F��L�ӻ�G㹍վ>>�kTu�:���"ck����B�Y�T)ş�r��!}����#�䟓�ү�~��ɖ/A�����'7M�� Ӓk$WGW��#��Y��u���������������C L�������]]]�vo������$"""""""�g�o�1�m���,)������H�$$Gzz������= ��>x��+	�^s8W�����q��q�������ǰ(0��l^��آ8�Ϸ�/&6�h�"��"]�
����ʾ�o���7�ckL�1F����Paf?o�٨����wUo�Io��;�cM�5h0����b�歋��f�:,)	b�>�L�;o�UH��|��qh�fPL��Ց�=���$�F��K�9D
�z��W���*��һ��oM����҃K���eЃ\��v_)� ��	��o��Z�q��%5�2d����&�����ͷw��Yo$��V�Z���բV059�Ȳ�ok��HP��n;Qir%�
'�v>�}4��yﱛ�`N]��}t��J��)�bd�Z�:,�%[2��z�{/?�""""""""""]�\������߿���ŉȢȳ^�k�F�p��!���!22�`>���"""c`PQ<�p~��z7G7���䭃#}�����~q;�~���9�3���k �'uf�I��R<;��T�Q5ڶ��M(A��;un���>�k���zq����s�_>V�4�����]��PT�FG��f~5�S1gZ״j�6$$�ڣk8q��<���+	y�����5�+<�=�7u^U|��!9�K���W��4ǟ�sZ�G�_�����"Y
�Q M�P,ڠ��[�����e8LE�ѳ|O�� 58,X}��7�G���$�D�ȓ:O��Vs��$��䵎�?ڠ���=���P<�x�g��� �Je*��)2�^BV�[������0���F����{~O}&��q0Els�Z��9�����P�ܣ�Gj��3���A�re����~��R����vޮD;���t��T���Y����ET��ϱ�J��?���9���[X}f5���KHh���?׸@cu�}��E���_�_�~L�t:�I�ͫگ2($F�1��V�(�(�wM��)3�dƒ��C����,G���T0f\�����ǋ.����'7�k�c����^:Si�Ǥ�EZ�P�!���r�ihH���#��%45U�T�)�C���Ҹ���ΛQ|\q5=����7�n�9^�s;&-8�@���G��|�t�M�*�dD�%!B�(�j䪡w��GADDDDDDDDD	C�.��<�窮��d�Ȯ�3�}n�G��\xp�Ba�ŭ����b��X���g.�~��`gY��3����(>1(��������(�I��;����'ڶYSfŶ��aىe農�*�Nl���ۊn*,Ư�,�0֞Q[������)�~����<�#��o;~����R�`ڂzۘ��PBJd���^Ut&�[ё��f��u/�W>�vN�N������x��]�^��~P�Z�Pt⾉�{x..ܿ`�<�!�9����
4R�ȶd
2_	������~x�хj{<{����r����w�Z��ސ�!Շ`ۅm�wm�M���7����}��1v�X�xrCsz)����hZ��fy�jz��*�%�qX�^���m8Voy�%dN֝=����-��B�2�ЩT'��@�$,�ȟELR�<��d�$u���R����b�=�_���"?/�N��U�~l�)�Fm'���H���m��p^��"鋨�Z�j_L?���A1�}���e�/�A:c�@�����s*D 1��}$�b�?�|���G��Ŷk���&��	r��ػ�
U�)�b�:t*�_?G|���em�E8'�*r��������l#���12�[�y����6K�1&.׮��Scn�ц��9�#�����yH([�h��ɸ_k����7�TT����6%ｄ�I؍�"�E��e1�� ��[Ws~YRf���3�7MH�6�S�u��󛛫���sp�}}���Lr'��
<q�N�>�<_�Js�뷯�FDDDDDDDDD1#���[��}�3Z��|^��h��!���Ig9�L¬C����+��cPQ�w�*��N�mP�f���p�����bFc$�;�{�-ngg4�� �(4<զVÝgw���\O����c�H��H����W�h� ����eY�0y�dT	1u��}L�?SLQ&��F2�d:�M_����UQ��J��������ƪ;&d�'�22L�{�
��^z�ؼ�xQ��(���a�?���^
O��V;/o�\��\
�紘��
� c����å��;�'o��vz)�m6��x7��su�7G7Lk:�g֎�k��g��B�ےζ_��n3h�Ҿ늮j���Gʞ*;~��z�2�z��+�
���|����S����_�#�t�lb�ly��s;/�D�U=p����@_
�eеܥǗb\�q�3���W�Q�.n����۾�v��	$v��W�;���+���p��F��/-�����_�6r��Bv]�P�Ӡ9���S�Gc:b��`1?d>�	�&� ?��T�7Lj<	m���l+�79�o��bkB�	*�O��&�qiG,9�$�yIP٠�0/dV�]�z�"!:r^k
����L}֝]�Ν�Z1:d(a�{g�U�h#=�R+O-u^j�A%�@�ee�jQX{���]s$۱VP�|O5p��Xgj��}��,���$�R��pɾ�����������ܧ��bry��yR�Q�wU��O�N`HODDDDd�CDDDDDDD� ^F�T��{V=t����[�W��7Ɔs��H!w��0�2�g��i8�!�?���F
1��+�o�ك�.R?��t�����Ǡj���Yyje��s��=4e�<{�,��Xd^{����n;5kV�
�c��K��5TX�.���L�QAq%�-#w�T���W�1}��Ja���\��|�B�)U���~��Y��-�-���'���AB�*O��Y�����y�fh�a˰���X��IM&���]s��c��yigDDF�x��SqRE���2���曲ߨ���0i����d�;�.v_����&@��e˺��Z��C�+ￄ�u/�]�4Jv0jP�j�L�� ��L�y2�g��&�F��Y�� 5-���F�T�4��>��F0R�+(�z��H�V�J�t�ys_y�]�vz�H��=�z�h��vq[�zzK�3ii^��:��qib�L�2hV���x�.�k���h��f�)�p���%&�(�r�s����U��.r�9|�p��:"V!��WqrEl�Y�����`ىej0"YW�d��Q�G��I-��JP]l��⃄��o8^�*���n���h��U�L%5��b��:�_tAXs���o=�w���cJ�'^�j���%��ɳ;DDDDDd�CDDDDDDD�@.?���j`s��H�,���I���;�W=�\?{��Ab���t��`�rx���['�Xdpˀ!5���lb�5��K�mE7�y]4��̪�͂#q��o��Iz':}�4jϬ�=�������=s�\�r����1��@j�e�QBb>&�[.l��H�f�-c�⃋�-��z�*��Ez���	O3������̺1�����Nt^�Y����g��c���7�t:���U�x��Qgf����'N��������s�MH�1��;>�!1�H؁VPLc��H�,�
q2�%:h�[{fm����?�/����i
�,�N����a�y�C����Nױ�cv&�,W^���Єq�}&���[`잱�G���]��k�ΰ�����q���ޱ����T@I���4��\�g��a>�_�\'�4$&����ձQ��brS=+���[�����a\HЛg�{�<�J�]�tŘ�c@��}�9�+�9$�KRu��}�|S?_}dN�9�i�_�=֝]s%�%�ϭG�&:��vm̠}�		���)�,-��D���5���ɜ�"""""""""kӶx[�l6Ө�����Ʃ~�T��<������L�A1DDDDDDDD	�ȍ#�:�*�tXcP��Ǥ����wc����a�8s��]��4{e7w�޾Xqr��\�6ߔ�F3B����۠o㵐�#��6=����n�?�q���8/�!1Q$�D�����E��c��5��8)ƶ4��ga�ٵq�����w��v�H�����qhLa��8y�d��1?d>�k ߂�:Ǘ�XB-컶/F����O���5�5$&���H̎�;`����_�
}��5I�Ȉ�#$$����跶�Q�)Ao�a�:��X�W��M��r$ģi����e�L�zW�*9��m#Eɉ�bu��Ȗ*�����J�e� $s%C�mP������f��G� �NWX�i����2��J�]Q5GU�s 9>���?M~��YCs��3k�/�p������g���:��������?eY�n�����_���9^�����Iϫ-E���`J��jځi0w�#�ﾲ�Q�%4V�4_�Ѹ�R������m���r-CDDDDDDDDDѫ��f}5˨!1Q��@����aؖax��-������|0(��������(�IAx�qű�o�ނ>-�7D����cUL�?�L�V,Uݼu��.)^�}kU*S)l�	�N�1�V��z�L�E���;�7F��>J
鿮?,�;�P�7R����9��x~^�^:���3�+������`�>w,�Q���C�&	����ю��@�|��>\���:ƨ^��d��kU/�x��"a-*��8���^����;�t��i��=�MB�,�b��d=�#d=6FPL�"-��>��q7����[�XI�ר���m7��LP���6ÎK;�XH�����"鋨�CB9%TF�'J�U|iW����6��WO㼜篟c�����|�f�?��پD{��#�E�c�1����{����d=�0<]�5Ϫ�Fn��2zU�쩲1.kʬ���v]�2�7��`���m�
"��oP�()���b��5�� K�/��rj殩
	t��]	$#�!���Z̃���f9w��JDDDDDDDD?��ׅ~M��|/�C�P m4hn�ϽY���/�����V��*��*R����^E������7��A�f9=r�J�*�TRl%E��C��Z
;�>��ܷ���ܜ���e}�
X���M`�)��v�v�*�G��ҙK�N�:����A��Y��n��%��m��,
ϓ:�z����{�/y��:�����&후;��e^RD����1���^�%`*s���1��:B��凗1;x6���s��C]�w5xy�K������&)��k�ΠQ?}��H@���7	R9|��I���b���O�$u�b�M_Go��2:��9n���0����p��*�+:F��տA�#�פ��0��T��{���s��2)�R|1ο��
W�G��P1]�Z-��úr͡E�ӌy="��[��
�ŷ�/���n�C�Ӵ`S���.��{�a��}����bm��0�v��i�����zz˨˓mw잱��Xw`Y�|�c"�%er�v��]X�&��X��e��/�=cŴ*�Js�ʵY9'�����x�����������(~�Q�����{,�1��g�U�����e(�3�^��N�4��ب�Q�1(���������L�MX�����X�j�f;)���
~��޾��bH�!���쯳�T�EGY���6am>�[
U�7��s��M��X�i]N�`ǣ��m�d車bbc��1��o",����uňi
�������I���/a#�bѱEF��l�i0F�>\�iF$�5cy����iR��#� e����˻��������9^�LA4�>���)�~1�\�rjۗ���@t�ɕH�B�l�R�x,]Jw�9�C�8�����TR�8	4����"�C���婃N�:�����{$ae{����7*�hىe�<+Q=�)�	�w���%����?��LK�B�t���4r�/��F�4�����;bJ�%����G���膲Y�b祝��+�W>����'�!���=�6O9�j���zߘ�;�k̿����>W=Wu�iH8�G2�M�W��]|�DB���b|r�������z�r$�ZdD��A����z��X�C]s����ʋ6���m#�bM;0���f�]ґR���u���}}j䪁-]����F"""""JX�]YCDDDDDDDd�v_٭�Ȥx^)�\m������1
2�T�=sï�,]�h]�5��k'���0L칲�!1�@�fa
��"�wM_����9塚��_��.��Y�'z��Kp��9��}ʨ����*���t����Q�7�۠B=�i�~��dtϨs���Ŕ�X)���9N^��[a*��t�H�A�t�p0��Q����*DDF ������j�.cơ�A1~E��om?�z�*V�-��Xr�m��
���6�-R%O��/g/����h#�����Aq#a1峖W��4��5Z�%�s5	-е�˾�R�Jz�N�_�]�w�Ɠ�/UsV�'�.�fl2ϑ�F�)Q�)GU��b*e��9N�*�GL�9��S+5��!�Z��<���P�B��pu�&�����ʏd���؜�5�}+�U�IC6��gwa	�����+Ȗ*���8�U��0iߤXϿ��c�.������������5� �5@ ��`c!Bd!hwwwwwww��=w�����������٧��p������nu�����L��#�\����
�C�9et�і�S�ɻ&�譣      @����G��ͨ�7OKPH�쾰��r^>(���L~^����g~�r�]����2�=�v���   DA1      >�ܭs���V)�����
�)`~x]r����w��gF�,���5pDW���j}e
o=�%QQ���䃊Hろ%F���~�@��E���?0�"��Y�Kڄi�Z֦S���o;l�V��l;��/
�����Z��q��u�M�4�FG�r���P%{˶�G������S��оD{�m��-(f�i{�㮝�w�;��U[�l��vH�tE^i�0�FɄ�^n��X�!*ds���
Y*xt��vN�o�|#�W��ɥoݾ�0Ci5��_��j��u��	m���*���e.�M�g"��kH�8�/�~�tz���T��m�;g�R�sz�Zw�����h(��9��'�y�QP�^G�w��s�\\*X��/�&��Ň�������L0�#z܋HPL�bm,�4`��3c�A��e���$�疮S�
      ��7f\iZ��e�ѫG�ʠ*nfp��Uyk�[淭�M�¬MWTV��Jj�a~'   ��      � -v��NG��IG'�~�)P�QA��w˾+u�ԕ�"c�2�� SpU$��@�o`�+�QGtqOL�~Ϟ?�!��ЍCM0��iQf�TyMA{���$0V��4Ò.Q:�6-�sǊc+,۴@wT�Q�X��%������
k4���u~�e[�$�%~��r��][���p��9�K�ϥeN[ز��������"���xCd�W�}zwDâ�S?_}ss����&���2B�L�b�MN�7�:# �$��X��Of�E%3�4Ǯ��Kg*-���$�U����KT�,4AC����0�K���x��=��{�D&g�#O'���ny�?u~����9+�蟄�����}�݃b^�# Z�$��P��K&�S�b鋙�Ύ��������~�6v�Xˠoʞ<�)(pW��i�Z�j���6V��4qQ�Ef?�r���R��      9j�i��v�ᓇ�ttS�Bb�N�)�k�j���J�TydM�5Rmp��b�	   �     ��Fn)�V�ԭ��LI2Iߺ}�:?ȆS��SwO��/��ґ�	�E���EZʂ��(,�J��5��E�R'Oˢdg�_���b[���Ѣ��|퉵^	�ɐ8��2YZ��+E.����h،;��Ro������<�
53��v����B�>������r��>g����?}�T�]�'�����s�s��:��y���+�œ�ܽbٖ6aZ[֡!�^'O������M�DÍ^V%{ɒ4��7�u,�ѲMC+<y �_7�ߔO�~"m�K�֝\����֩T'�\����@�����R)�gy9~�DeV�	��$27�N�9镶6��8\֬�����;Y�|�#E�v�CQ\]��gگ
}�t�R�l��1^V�x�8n�/+^�xN�]>$�t9��e�]�yv����kJ���>Qzs�~��;���z�4�����-��$�j���¼L�)�������r�{�@�vv���i_w��s�`�����O���eυ=       �T�i}_�w˾��<��V����Z�H�j��������VK�AU���#    r     ��tt�6�ۘScDw�+�qVt����f��{gȌ=3�j���a�ĉG���M˩�d����/��R�a�o$�s�vX$�*��sݟ����Z����jJ�`y����ש�0�Wx_�f�jy���~���o�Z�jan_�,���c��ܭs���BYvd�	��"Voy����|�#˾~�	.K�0��v-`�#(������w�:�F�s-�<��+"����hȁ���۲�{�����^��p��m�(�E�ۗh/_.����i����f%ds�����5l�0黼�\�sQ1z� �_W�*?����X����=���8��	努��&�)�敠�ҙJK���Y4t&2�<V@,�vO���|�i��#�o� ��X�k������\�r^�^��y��Ǖ?6����,d6Y�d{���,�F� �(�7w8����l1R���.Ǯ_6v�X��<ޠ� ��o�sɴ�����<y�D��in�a      D��K;�������umY��?�ga�ua��h>��1��{M�5R}Hu�{q�    �<�      ���6H��-d|��N���B������'s?�_V�"�NQ�u]fF��t�y����Z��u�T0�Ì�^ֺ�����D��o�ЍCÜOtS�O!���lɲ9-vUoK��M"�G56�b��'U�t�-����}}͉5ft�>�����t����%�6�Ҡ�Yvt����*�Eo�d���X�hȊ]��[n�p-�u$�����: ����xKx���o��0��=l�0�A1J�b����s��o�Om=�Uv��%�;=6�9�F��.SvO���o
쥣v��՜�F�e�Oj��{�ߓ�V�&Q�UhB�\�$E`��	�j[���e\�sIZ,�)�s��{W=��ºtۜ�$�*0���{��nײ�O����Ů�<���7�}��5d�����jC������WM�5I~����k}���h�J�ߊ�+�M�G㶏�.��m5֜������s��       �K}ț:��6�=�ڽk��oʮ)r��y��i���4����]�   D2�b      |ش�ӤFh32���]1��<�sݟ��4�bN�9� )��P���ሆ���J�eZ8�ӊ��W�^榃��b"+�h�G�����ݫ�s^O�����H�U�H��On9_�|���7��.S���t{-�����/}i�v��	��!q��~f֟Z/#��47�h!�'iP�'9���<�����'���a{X�!Y�d�bǈm�r"3��uGbH��Seυ=R M�W�2&�(5r֐E���=�v(���=ds�Dڇ+�JC�4 �Lnʍ{7�쭳���>�wi�<~�X�yZ���\=�Z�Y��\?У�b�6q�D��	���5�����0�慛[.�S!zVc:m���s�Ȱ�����o��s��=�'�b��#Y|>��s�ǫޝ���O��i9R%{y#�2��|�U����B	��]�	�	�iS��e����yZ���o:��`iZ����>����F      �4�E��Yqt�G֩�UTUu^dy���Ŭ�Zj�iD   �y�      ����WK�~��*�J�r�%i��.?VG	Yvd���6����;�N�:f��$q���B�_�e�)��uկ���,�#3�͔�R�R3gMɜ4�ˏ�"q���M	����]�W�l"C�qZ,ֹtgYr���:ʶ��~��o0���q�봮���v���O�#*�B�{�����G�?d���������	�qR�'f[�a7VA1a=���'D{>g��oy��A��oئa���v�ֱdG��b�d�b��vL����ؖr��9��k�_� _��������)�E����}��Y�&�-���A1�`6f��la�~y2�+���81���m{�P��)vń�������D��z/�-+ޱ���V��O�(���*(F�>���K�m���*�ʲ��F��Ǻ?J�R����oU?�y��      �;��WP[�z.�E>��,�DR�p8���(x�	��vv�    �,�b      ���GwMȆc����P)k%	���q:r��;e��=>7f\���&'z���=���'�3��3{ȥ;��W�r�L�s�s�ˡ�eƞ2r�H�xj��?ݸCZ�ma�I���b9߀Fd��Ur�����R�J2��@��Z5dér��A9}㴜�y�l�7=}d�+�$��'�;�O�q���;��44�jD'W�����<��H�o.v{��x����q�������za�ÿhA��j�e������L�=Mn=�%�7h �8Z���Z$*�(3p�P2cIə"��kh�#�/���ͯa��<y��>�^oZ�31�o��m�����=��<��Zyl�쾰[
�)�]���$L#n__5g���pr�7�kP����|�򖁲zM6u�T�o�Y��|R����2R>��|       ��l�+�W<��]�wIŁei���.Q:��� x˺.���js�   �a�      ��Ї�2x�`3%��܌Z�?u~��c�{�ߓ������eѡE���9p逜�yZ|A�<u����%iy�i�m��5̈���B���`�7U^)�����UK*d��(�e���̌4�#�����}Fwɞ<�T�Q��<z��x���#"�Ĉ#ÛwZ0�E�Z�=l�0�qn�<y�$\�J'�x�ބ�cF�nQ���.�Z�f.�P*�Y���TZޝ�n���#��œ�N`�fW��������<�ｂ�i�֔]S�]�v��iX@�bm�5X>^?�oxӲ=ds� �r���rf���X�a���4�QFԜ}s����Ge����V�&���s�X���Cz�T�J�X�~��^ga-���$g�w��'��Y~t�eP�~6�e.��!)����vɷ�k�ƕ��ϊW	��M���;�GC;M�$ϟ?       ��(�����Vq�2��	�ɐ8��yt/�:Ցu'�	    � (     �O]�{�(;�yA��g(n�4tF�btTk��޻j�y��e9{�칰����J�*I�j�����?Z���J�ҝ��eߛb-O�jQd���LH���20��R�OaF~�I��]Z$�)���(F��c[ȾO�Y�&T'O�`~��\:X�&�jٮ#5�D��:'� �=��a����8�L������	ܩ���)(���2�Kˣ'�L��]�*���5����C�8	-��zZ��L�&1���6s�:���4(�e����kұ��j�i����A1$�#y9t�DUzL�~x�R�^i��s�ϙP��i�}��q���V��îݻ�u'���i����ϑ΂d�ƈk�J��������<��)��]fAԵ���G�X���TƧ�b��\Y���W�|V�<�c�x=&j����{'D�i���7J�h�,����V�Z�      �=}d٦��u_�����ʛ�p��]jq��Rx}Yvd�    �A1      ~l���ҧz�������yS�5�����К��h�PP� �G���aM\&��d
p]��L�9�֑_����	�	Ͼ�9��x�ޥaR��XF�m9��D����p7�-��e��k����N��ݡ��M�+�3��ґ�*d� ��V2Z��3�^��V��l8����tO�8Y�vמc�'���ǋϲ=���1<s�̲��N���cҁK$O�<��i��m=���c�
���������x��+����N�:J�(5p��v_����c4�I�8�����N۝��#*Q�DNۯ�w�m�Ρ^�76{*L-��W9;�k g��1L�"��ˡ���[�(�K^�2&��J����,��:���urױ�����|K�<u͵���O��9�M��'       "ύ�7,�t�������~�\��
���Rɗ:��y����gK�e��%   �^�      ���W������
�{d�@ѐ-��ѳu��EZJ�xI�˕"�i2D~o�L�3�B�8�B<y��n;��+������s^OAԥE�p��&�hȑ~��^��
�S�vئ�|�Im�Q��y���?�L*M�4� _i[����\6��S���k���ET�q$y�䦐�nZ|�6aZ���w.ڲ��ҋ�貵X�JX�Ao���WC�ɜ4��<OP���i��Z�W�mz�t��I�rDC�a��R�%��I�F�>��&��qJ2%��J[��>f춱�-n_pڞ!q�u~�G���5����Mϑz�iV�A+�
�I�؞�Ù�g,���K�s��IA�VP�?|������KϪ����k㴏��V4�֎�اr��2�������m�z!����{      �7ܸg�20������,z�D��UeI�%�~G4,fN�9�lL3��o�    �A1      ~���^R*c))������"_.����iq_�Ty����Y�L�����ƌ+���6��hX�e������n�G�����?�}S�nW`�����i���+�Q��Ͻ��u��YΣ�%SvMq{�q��5o�<9r���)K�,�k��z���f� 	��V�Z�r��ɲJ����m�i
������hٮ��v���x�ҝKb7}m��|?̑���V�ȳ'��=g���3z�h����44�������:��h����� D����j�4��>�����˥���>u�T񖻏���{�-)4��E0�ݬn�U�뼬�2z��@���h���z��`N;h_F��P���s�Y���/߉��6�2(�J�*&������󫛧��r5l�C�C�Q|���\: ���6��       |���o/�b��V��'�}�W�ŝK�tEΣ��Ln;Y��nj�W   `�b      ������+�L��9kFxyZ����Oe��N��?2%�$��7���'el�0NB���k�EX/
�t�vv�)�<x��)�9s댜�q��Z鿶�l9�E�7�/�3��6=x�@ޛ�	BԧEfP'O��^ҡd�a�[�u�1s�L���[v��u�A�����{�߳�O�l�I홠g�ZX��	�֥��A1Ξ�{5&,;����������'����nBa^�(N"i\�������z���Y�<
_��[΄>
�ׁ�&��7�z��~ߥ}R!K�m��c�!4V]>�R���K�-�b��/��;en�Ӗe�>�c׎Y��sV�Ň��d�9mw����s���v)���+m�L�ߪ~��5)��ah�Ұύ�6
|���w�/	b'��G��j�!WB�       ����cs_���f�g)/#����m�z��	�Y�PJf,�p�y�[S�Ř2c�   q�      D:r��ސ.e�H��}�(��u���Q���6�����($��M ��8���ΊJ�48FB���y��5Ġ�27��4�_�$��3����oƈ����'=�����
^_-��2(F}V�3�y��I�U��d�l;r��)z��7��=0�)���	�r�b֊���D��	�^k=v�Y<��a鑥b7g�aυ=.-c뙭��֑
Y+����_�m�0(F�]���	�i���e1���L��$L��ƽ�:� 0=v����2ަ�#���RKI�h�L��N��2��X�ﾰۥ��k��#�곕�`�r���jS;WmȊ�)m"����S���[�(�s�,��� x��<먾I�%������RcH9w�       �M:@�UP��ܸCj�)�X�n��Ni7E�Oj/�<    CP     @�E�����GH���]�vR%{�Q��xj�vo����l;�M���.�n�2Ӆ;���[�����Η0��p2&�(��d�lɲ��}]�m>2i��'B}��<#��L���!.$ j�rf�,>�Xj��=K�,�`Нъ4��ʥ�Kb'W��+�������j1�a{D��^V/o=sް���p���Z[�ո`c�a��.S���rղlw�98��#�Y�g����V��+�M���*e�d�Ǯ3�ݱdG���:����*l��׏��B`�
��zEZ$ަ�w˾�M�mJg,-Nm�u��L��9�&W�|V��a�K5d�ڽkb�&�����^*-
�pئדY�e���^����DC���g1a����O�d��+"�R�}�����آ���h0ո��ާ���.K%U�T���1V9^�[      ��]�w9����s�� /ݱ��W�y��֒���[��D���Gr_   `�b      ��O����Ǌ/�rT��%�K����u���#Y}|���?O^$/4EJ�z��R�50�v��f*���D�M^':�K��}e������~���A1�󪟛��Ϟ�+��1D;YQ�*gE�bbW�K⸉�{:g��K���${����;����a����
q��s��쭳�>Qz��V������/����)�~��:�� }�1��sT�\�����z>����e��	��>/���;'J����&�}��O���8��O��SZia{PL�����/?�ܥ�9������>�a�z��K��R5{U���sM�_�h�_i����ʟJ�i]Q���V��4P�_\�sф����)�F>�����U�V�y��BG�/u�Բ��ɐ8��<�ܖ��j�O       ߴ��:����W��S׫�;�yxG�����q�T�V��<�[����    ���     �(���{f�u��u�E��O��Q[F��]��H%v� -^ԩ��ޒ1qFi]���tD��A��I�J�*��|h���H@9S䔦���iW\�wݲ-e`Jۊ5��a���O�޽�]���Q�Ju�5(�s�Ζmz���Ë�n����缞�-��s��#W���=O��>N>����ҙJ��O�&�Q[Gɷo|+�b���V�����_��>�Bj�_����! �ﳢ�~w�����&��\�r���6Z|�<h0C��e��˗�����oڲ>���eZ�{q�����ca�l���
���!��{Ktt�:B��K�V�Z��<���oMh���y�;ET�O�2v�Xˠ���D4I9;�r�]z�^�y��H��r����K��e뙭      ���wy����G�2�-����>�:Ց�fJ��5   �g     EiȐ&C�J�*�i8� �[�O\:)�<}����3i����7���]l�k�Xl��{�E_�k���Ϟ
^o�-�NtZ`�ޫZ/��k�KE���P�e)g
��0��&Xş$��ܲ���Gr��]��U?_}�����>�:��ʛ*�t,�Ѳ}��Y�0�n�O�\����y&��j���T�R��]��1d����'��!?�,��Xe[�"�ވ��s�BM_i�p�7r�!틷�|�� �@b����t�y���݄v�/4��*(F�Y���ќ�lY�W��r*4v�{!�vN��)���	 �#�R�U=��(�w�����#����O��i.��ƌ+���/��h?ݎ~ud��w���?0v�+m�[!kZ$]��\�F��4�'a��� x�HS�r}���nb�O       �A���Y*���z�M�mȝ2��|P�I�$S�M�zy�	    �E�     �א�hz��}L�RT�-Zp�wy_9��׶c��ufʔ$�	��P��߅P�#~���/���� xJ��8�C��Zxp�l;�M��/�]��4hC��r��i˶&��/+����V���X|�cW����_�~����ʓgO½�hѢ�c�� �?��)����� mƷ��r�Ĉ#?��Ѳ���n|��~B�o/m�9޶�i
J�F�����2l�0�A1����9if�m�ܒ���
`%i��r��u��G����Mv8��b5e���� ���|/��$r�޽|ws������e�Z���÷�7b���hP�ն��N�C澩��$��X<A�o����|�H�B�L ����MC�F��4�C�u�����A�w���Ү�㐬�E[��X�Z�`~����U�R��C��w�Ή�^���gw�-%2���G�ێok�+       �eѡE�bT�bm�����m��b�Q�eJ�)f�"    �"(      
ɟ:��k=β(-*����.Ǯ_q��)�2�����'3�x��-LPBT�� ���,?.�Q�Z�U�%�߾_��L{k�e{�j�]
�Yyl�|Z�S�m�2�2/���
�vV�ZQ�4"vK?����wZ���^ۗ=@���nپ��z�ש���ӺJx}]�k����e�lm<�Q<EW���"��#\����Q-GI��,��m�\�������ҤPD�Hp�`�y��|6�3�C�^Ȗ,�|V�3S�z��aA�-;�L�_;.Y�e}��*$FM�1�* V�Y㟦���/e�I���*Y�d2��$������4���v��m�~�����a{��X��Vn@9s�	��3Ȝ��8��"WB����;� P������z�ɨ&f����X���p��������N,��w�K�P�u�ǶC��W�X��n*��~B��H��5�Χ���W�,�HC���b�l*���iY�����Zڄi-�VU��½���J�*YΣ��~5y�d      ���gX��_�vɷ廥���oк���4��m'   ،�     �(@�H�-����e�yD�H��o���o�����U��I���H���$s�̒&a۷C�Xޙ��,8�@|��״�J�nj���'Q�������������!0�/헼��:l/�������0?�������E�4���+Ԣz��2��L�+��ME4�DGk�������tz�-����u~0žVf�!�ХLs��f�7�z�X���O�~*��k�_�❋2i�$���{����Y�f���}tW�Z�U�������gAs޶�I�O${��<9X�ݻ&v)���)�o^��	!
o�^�� ���߹�8}=����b�y��=0WB�Fx�z{��[�S��L�3@��p�}?�����L�]�l�;/�z!��<�p���%}�����⿖�K�C�=�t��/_�(#�ߨ��������A2��`��y.<�P�n+m��qخ�ߑ�G��W�SGԴ�>��٫��U?7�gگ���=��S����GXFn)������rs-����%������)=��?W�����Zz��̇�?�
      �1��`����0�W�4�����H�U���� MF7��m&ʛ���cI��لg�zL�x)����   ^o�      ���qʨ���^�ߗu'�Ɏs;d��}����������5Y�e1�1E�1�ڻRLe�M��?��(62�<�R��VD���y�Z�^O�=�37Ϙp��w���+��O��'�'Q�D��2i��毎r�Q��Q:Si���i?������
�.-���񱭬G��@���b4xc��i�#�'��L�t[#oM|��B?���^:��l���Ϊ�1��8�A�f�c�ĝe	r���p-O��YZ���C��r����7�9���׵���)s�{3�3Ǟ��1^�m����t���������n`�����Lh=����^��9��ECδ�<�Ѭ�]��ه��տI�ܵM��-�����X7����8�#yi^�����/�[F�ύ��B�Ƿ��*��j�i&=��͟P���v9x���/�B��d��Qm�����3���O�}*�n��>=�<�c�r��<%2���l7!�s��qi�z^�x��N���|=���+�W$<�\�aj����<��ט]�v���¾q6v��&<�O�>�\���w�K��=�l沒5YV���o���GҴPS�y��&���~�#%3�4�v:�5 ^�-Y6s=��o�o���T,}1��%G��������P`����ԑ�e�Z>vʮ)� Y����J��=nXɖ<����׭����p��=�W�^Ҥ`��yZR'L����z0      �^c����_P�S�q���c���ci6��	ҷ
�]��
5�;bō%    A1      ~,g��2��Lɓ*O���A�0��|YulU����N�e\:`&]��w/�����zp�N�9I�����ga�!��dr�qϟ?��+���C��䍓r��Y���.y��f�s-.���T�V�x��M{k�|��;�rї&<��|j8�a:R.s9�����8���r���_���*XItZ ˎ,37����r����GC�*f�hF"jR��	�y����c�?dr���	ZL�M�o̴��N�xj�	��zv�9&>z���h��#�p[o��������Uxw��q�pr�+!/�S'O֥�[�}�5C�oろ�K�.aTiA��xsM��U��o��~V�3iS���0Hf�!�����M���+j�k���5�pj�����m�#��n*뺯3����q���*~ K�,5��5�ט� =?���/I�%1�C-f�I�'�A�p��	\�0Wh0 qc�5�]����5����&$D��W��I 	c'��)$O�<�O?V|��7j�(�a�����5r֐���ZΓ.Q:��q�l>��]�9F^\j����r:��(�3s�SwO���Fh��|ݨ@#�aj�79��A�u�	��|f��S��u�.G-]�i�F�=߯��M?uC�� j�ߨ�|Q�Yth�ٞ�'�ʹ��^�y[?��,��8ϗ�Tʄ�9�w]��������+=�X�83v�X�4��C��v�Ϣ����sA1i�	s��<���b��T�      <a���r��5����w��y'��5�I��h?���W�]�v    b�     �SZ�7��I'Q��q��=ST7h� �vv�x�����OH��z���~�gZ�W�&H�|��aο��n�5�W�׫EKˏ.7�ٓg�7r�!urב��+�D�d�@�BiI˱-M^d���ehS�����z��!*HҥL��U�Q�L�❋r��u��#�;�	��t�w��+Ǯ��P8ma3I���7-���Q�n-d��_8��W��4s�L[��ׂ^���Ad��-�I_�K���ҝK&t U`*�`��i�y�Q�M�'�O	�-�oy�([�῭���t���cd�����;i6��-=�:�ZKw^f��#�50��<�ݽfn�Ҁ;���a����㶏����`(��6k�,�<����t����h`�3%3�4�zS����ԝs˖3[�㤎Qz>o=��l|o�dI��r>=7�S�3)�~�n���5�Ί^���^Zm-�r��Ay�7d~��a�O�O�#h�}M}������1b
|��1k�-{/��aJB�c�:y���=�V        ����oxV���(�F��8���>
�RK��n��v   �날      ?��lÛ�X�����׎K���e�֑+�Y��	̨���BC�т��@�G���$�Y�� :�����v;z��y�u҂��%�K�2]_	�����A���2������Q[G�5����;l�`�2��ȆS�.��Y�ҙJ��^-��U�,�FFo-E�o	�h��3����a7v����^�f'����<��k�?}l��7��,����c�˂�������;4�'hx���uV�˪8��Lo?]*d���c�y�r�ȱ��b9}�dL���|3���ɛ��a�����S��hJݿ�����.��TX�&�l=�Մc�yxG��Nz-���r��u)S�),D�ab�y~�G�b��{*�YQ�t�cB{�;FlI�0��,=�T�Mhg������ʏuty~���       ���.�F�b�M�&    "��      ?�A��_P?S��.���%����ͨ"���
�PWm:�Ij�%�ܒ�D_��&�e�v,��r>`�P�%��xt{4��տ��k~�j٫I��=�~���,[G~Y�}��R��#���������~���O�>R7����<|�P�j,�;/�|��ٶ}Z��������:�}��g豢�CWI�!�e~��.[���rlK���D-�m2��Ll;Q�Ĉc�2��W���v��4P�꠪�Uͯ䳪�Y��M��4����B6��׵�v:_��|ե;����2e����*��HH�iU��G֡�I���M0���_�/�U6A7��d�e�z��4��L�5Y"�>�"����K�"-#m�ڧF�8v��Y�G&��BR�o/?���ٺB�e            �Y�      ������n?N�4X໥ߙ`�Ȗ9if����.Ͽ��n�9���~p[�"-��,�bI�bm,����&� 2
�t�.��e.'���3A/�+E.Y��r�4����uN��8LzU�e0�F�7�h�����v��9����_ZB��H�B�"�]��u��E��'v}*wN�Z�j����W���ޗ���m;�M�('c[���`�Ž�|LsS$�f�e�Wƴ#ْe�в���v|[�x�x���Y�G&� ���Mj��u�v\Fn)���"��C�o._��B�8l?q���8�B WL�5U�&L+urב�؁]���Z?H~X�C�틿�<y �ǵ�Y{g��0��v�zE>�����>N<���R���2���Z��yF:L� ˎ,�Ȧ��V�Z��^�HS�c��~܈-#L�<G�gYpp���:��;�:?*:{��h�mX���b>�            �,�b      �Ļeߕ~A��~���҄�x�HkQ_���\�_���B��|a���H�Y�e1�,�迿U�-�ed�nۺ��L�2&��o��&�'"4�ay��RyPe�p�� j�������73�#ѢE���{K�Q��\����B&� ��������=Z�<x�`鷪�)~�}�z��=�T�ZA��+U�W��i
����Ϟ���Q[G���S����Y�^=*����e��'U>���3��x�����'�s��������)�ka���ҭ\7I/�[�?t�|��+Y�]�g�Ҋ�/&�Wx_�o(	b'��25lׅ]���b���ĚH	!{�iQ��k�$g��۵�?���~�7�)N�8&D*(_�T�RAr��m��u_\r�9ߎ�6F�<�#��&�l��}G����~��\?Є�j�Ӯ߻.F40A1���/��r�^[jP�n޿)ޤ��B��ڹjK�rݥz��&@4"�����Fs���o�׮��*���F��z̄ jS��wݕ����c]
��m�            ���     �M5����w�0Č�~��}�j~%��Uvi^-R�Q�O�<-��\�2�|�GR�p8��6���*9q�D�n�L�9���o�_ڗh��i���N����#���u�hd#�=�ö�#�e�/��c幸P���̽3ͤǒڹkK�lUL��Q�LC[]>$Om�Ȓ�K������I��88��3��M�<{"+��0��+���PB�d*c���s�#EI/��2t[w��-��m��g������ܭs�-���|��!&��~��R.K9ɕ"�����M߫�7N���M���s<��������W�M�9_,�B~Z��	�	�$�2��,I�����=r�,?�\f�a�z+Pe��m�nB;�#�T�^Մ��X��K�����k�!?w��A�sq��<�R.ݹd�v��������x��X�/�~�[s���� ����$=����O�vO�t��~���a_��s�[uR��`��鋛���y�Y@�#��>���Å=&�`퉵r9��Df0}�t���&���_r�[��VC�t�����T�ZQ��+��'w�j9p���.Y|x��9��+��_���f�7Mp��>�n���'e�٭����cy,�>��˾w��=i?U�Dq��m��eM�DC6��������iߥ}�ߨ�y���u��y>����M��{ߙ8�����üEC�f��|�4���V�jd����������l�����x���{Ao����           @�     ��Jf,)�Z�r+$F�ޚ��L�=M��fΚҫZ/���c��Xx]h��{3ߓ	m&8lO7�Ln;��h�LdӀ��:ȢC�dp����1�
�-$�[�7�&Z${�R ��mܸ���j�N/$����&�����ޣ{r)�����zb;_�c��۬4@&0v��
��q��NC.nݿ�@O�`���IiA����k'F���9�y����m	�����`�t�S'Lm�����	��bF=��(&A�c�$L#�b�}��>�Ź�>hѴ'?7�Df�qDu(���MC��<#Q���Xr�*o��v�z�aj�0NBsl�c�#�8����c�2}���3��7??�_Ґ �^о~���̾��znѐ���o�/�P:���I�'Jo�Y�u�<x��E��Ru>o�j����'J����2}��1�y����aOo���z����4*��uSx��6��S�=���5%           �A1      >L�f��i��\��|uC���Sśt�Ǵ#ѣEwi~��-���;'J�R��Z�jۋg(.��"=f�o�m�tz�Lo?]
�-������hF�"J�:�S�������Ұ���̓�O�?����A��XҦh����!x�J��KIt�'�'9q��D%�O<~�             �#�      ����2��XI�0�ˏ9w��VK�]�'ޤ#���4_R�t�1�^�o�+J�ӷK���Q��u�u'֙�o��*���쎳�B�
�^·?�U�Vɜ�s ���y��"0�ö�w����s               �b      |TϪ=�R�J.���I�2����M�bɴ��I�4�z��mc�u���J�}a�LS�r�-F��[ge퉵�-7�ߔZCkɔvS�n���ZF�h�dx��R�_!9��  ��(�òmĖ���C               �      T<Cq���W.���-�7���Cb4 �fI���z܅��صc򺛳o�Ӡ�81���3�\�rr��!����K���d|��Ҥ`�p-#y��2��(�9��<�\  �
�d*#%2�pئ�a�	               ^�      ����2��`�ݵ�n�<{"��4�}���}[�[i[��ۏ�x�@d�������ϙd���N�L�2r9��x�㧏�����.Q:S�sT�VEZɸ�� ���G��m�-�#W�               ^�      ���e�J���\���Y��co���gҫZ�p=6a�����κ4_�dYeN�9RmH5	}*����i8��lzo�dN�9\��%�����zpK  �gE��f��Y�\?P               �� (     ���L!������'�$�o�Q�����7܏O�(�Ď[>y(�3w�RJf,i�b��UW�=�'�r9���u�ׅ+�'u���u�����!  ��x1��_������w_�-s�                "�     �!W�X�M�ҼW�^��f�'�֡D����ZF�q�t�Ҳ��*y��L�����U�YgIPH�<x�@�e�Ž�cf�bT��N�w�տɩ�  ��w�[��"�X��͒o����               DA1      >"E`
y��.ϯ!1�C/�7�)�F�j��D�=��jU��k�+E.�S=Gu��n�4�X?},�2z�hiQ������+ �|Z�S�6��  ��l�?���1bK��TR&S�����o+;���{�               Q�      ���+},��]�w���2a��&��|�-!1/��{Ao�z������������K˱-�ɳ'�-]�v�=q��طK�-?,�A��:+  �=�j����>{*��v��ϟ               Q�      ��x1�I�2]\�W�?��xSp�`�d�m!1J_��� �S��u�!AM6��l"�[?���[�㧏�N�<-=����ot���cĖn����?  ��~����3[               �A1      >�y��(N"�杰c��zD��G��G�?$Z�h�/�cɎ2q�DYvd��n:��,��&��2�j*qbƑ�����'��n*�Wx_r����c;�� _.�R=}$  ��9��H��               �A1      >�k��.����S�n�w�-�T�D~���ǖ=Zt��v������v\^i��/j|a˲������4<HB�Jd�}��e�˨��~l���~��2u�T ����2B�M�&O�=               �.�      xY�4�dƒ.�;e�9x��x�W5��/k~���$��T�w�/UU��/HT+ �Lh=A�Id�2+g�,s;Εz��y%,f��qҧzɑ<�ۏ.LP �/=�\�].?��YZ$               ���     ���<ﯫ~��=Zt�w�K�r�"m��R�﬐ZCkɩ�$���vhӡR)[%ۗ��\�y�����ܸC"��gO��e�ˈ�#�~l��UMX��{����<�#SvMq�v��	�ش��$F�WV��յ{�dυ=���Z9{�                �BP     ��5�����]9$[�l��;Fl�r�4-�T"���l~�4�D֜X#QM̀�2��HiU����Q&SY�m��1�H/\�}��T�'I�­�i~���d����~n_�fc�	 ����5               �*�b      �(S�LR8ma�����Ȕ0NB��~�T�^U�%e`JY�u�|��[�~������
�%J'�[���Y+z|]�S�u=�I�a����Y?},�wM�n庹���                 ��b      ��^�z.����s�}�D�T	RɂN�H�"�m1b�׵�����K��e㩍��Zn!�����G�:3&�(k���z!�"���c|��bj�%�bɣ��                  �AP     �U�R���6��$Ǯ�Ȑ;en���<ɚ,���b�����eҮI�υ���W��?)�����T�Q�+�O/�,�L��n*�̏�un8�A�_;���?V|)���߇                 ؉�      /*���K�-9�D"���Li7E��M"�(Z�hҢpiZ��L�3M~^��l=�U|Y��e�g՞R/O=���/f<��a��;�]�i������s��s������ǖ�\��                 ��!(     �K2&�(��wi�u'׉�u*�I�9Pb�_=@�jf��v��-#e���r��U���2�\*X
�) �$F�2��Pə"�|6�3y���G׷�Ȳp�h�N�U�                  �AP     ��h�+�>{*Om��vD�]���+�T�D�Q�tE��k�_M����se������~y��y�l���6T�VE�o e2�1��/���ǒ=yvi3���}t�c��tz�<y��Ը���                 �날      /)���K��Wn=��m�(cZ������Ӱ��Y+��z?ɍ�7d���&dg��}�u<~��	މ����K�d�$��R0mA)���	�I'��}�W��J��/�o���:4�f繝R<Cq��:AjI�B��^            ���w�Q\o��oHB������]�\K�ҖiK�O�8(��N^�	\B<�{��
dg}�@��\!{Μ�����<��b��������M�t���`���N����R�'"OgO4*�HM�D�D�v�m�"?�x�ШP�F�":6��������ƑI�K�{fW�%�RYJ�Ч���f8v��M��/h��A1B�#�!"""""""""""""""""""""""��b��������I~��F����՗ݰ@C��0_�$'������USR���K<	����O�m�j�ӥN�~�B�,��z/���̷���`P�A&�'�}���������������������������CDDDDDDD�(�R�!w��F����Ֆ�"E
�5?��)S�%	����?�~y;N�9���N���K�����_��l�ِ'm�)���UՔ�5�U�������C�,�1x�`����Z�~�#_�| """""""""""""""""""""""�1(��������(d��
G{G��Z+(���s��A��-�¢�p5�*��?AdL$��=���<�=Ք�-#�\��;|�0f������γ;F��2A��Դ��6L�7A��P-��D��7]^����*��x��h3��>�5��66L������������������������(9`PQ"H�����)��4�-F.�\H
�?h?v_ٍAp��%�
�ep���U�I�,�а@C��Vv)�𾋍�ŲS�0�<^?h�q_�|��wO�釭?��O�>�T���AD�T�UGE��[�`KI8г�g*�����>!"""�j2
_T�Bg[��}0��ti���?ޭ�m�ɥh;�-�������������������6CDDDDDDD�|\}��'��a�)R೪�adÑHe�
�$���j,:�;/�DTl��c����-��;����ӢI�&����(���G������q��q�/��ͣj�eV�~����JV������7ǘ�cT(�%$�H�"&�c���������$�4�wn�T�d���'<�=�d�>���4�)�>��s�����k�{��J�&P(}!�P�}��5�������q'䎺�y58,DDDDDDDDDDDD���\���쥾�x������b�����������^<2{�\�aN�9hX�!l�䝓�gV�Z���p��-����j���>��9>*�*vK�xPb��oqȊ��hq��a�w,~��z��
M%�B���B�<��eq<}h�:1(�(�8�9 �guR���R�H��KR�,!_AO�&�����}u���I��S��G�����E�oDD����ʧ(������~&$<!�Nb"! �لtsvpFUߪ������)�Y\\��_�Uv�R��2��z���t���[�/h�o����ᛇ���R�u�/u��T��k�,�P:Ki�z�j���?v��`�U%g���CB���<HKDDDDDDDDDD�����;y5�j����
�Whd(��9��w`��E���������:CDDDDDDD�����3�p�A���f&2�e��칲���?l��-A�P\?���F��0��xU(�T�ym�Q����A��Y���OƟ-�D圕�G^O'??	��~��Ӭ1̹:}�4�H3,:Dd<)4����*z.��rx��~"�&A��p��q칺G����?��g��*$�V.>���W��B�헶#*6
DDD�Y7o]����Y�ܡ�=%`"�e�3��e�bmЬP3T�UM�Ř������R���M=0���N�+d�Tc��E�\�M�O�E%(G������o;CDL���;Jf)�:F~���eTX���2(�@��]�7����A1DDDDDDDDDD�X�zd�/~A��m�_��誂�e�����x~#���5N�9"""""��b���������wjo��Eǚ#oc��E�ҝa+r��/����C@P ʎ/���>��h8�;!)�qh��ȘH$'�D�)��e�/�C��
A����lèݣ����n�����_��tX�b���h��]�W��22i^	�ɝ6��Zk�n;s���3s��Ž��@֑/]>5�*�K=��&a��xUXNDDd+rl ���q%��
����_f����3���g�������ː�K��%�!#6��Ā�	�*R�H�����5���K������R�Zmu��,GBKg-�:&O�<F����l�ФP�7]^|/�%�źB"B�E��<�����γ;F�+���$����	�����?�m?%��Y�A1DDDDDDDD��ؠ�����lY�%&���i2��J��o�c��ETl�|I<y�d���R��vR0f�^?8��M�_w����bA�����1䄁�j|�f����Ҟ&]���"T'��D����ʩޗ��t�j�s���k�_�}��U!��=Y�����U쇁�b��� ""��\޹0���*4F��\?��`V�Y�+� ˒���$�z���o���?���\\���R4*�Ȫ�J�`�� �-�ê3��:v�l��~���������������X�b�<��@���%@�g������7`��a8��ޱe�ojc�:�Ō$���O�=�)�G�CDDDDDDD���1&\CBR���E���SwO�ゎ8s����wN����X�X]q$1I�|i���}�'�ǒNKT�9�ˇ=��`R�$u�_D�08Ot�yA1ƾW��'{'�5\��
����..?������i�Sf�"E
x8y���GgvϬ�	2�^�;~��;F�����z2�eĲ��0�>_�y�#"�O���1��5�T��.�]�/S>���u��U�a� ǁ���Bݼum2����gǖs[���Z���Cb������������D���uF� cI�f���~���0���.?��_���Զx[�E�����H��<΃���M��3�'�����CDDDDDDD�R�~��&����n��=T������EpdL$�����bN,�[��EZ&�:�92��y%$"�f5�c0��@�Ɛ����I�&�i8�X�7����#]`%Ge��łT��.�����S˱���_�GpX��1=�=Q9ge��S����#�1���P����ӡ�@�5�� 8�;� ""J�9rR�IputU�pߣ��$�nNn*d�������f,��=7�ꤪFl�jZ�iF���}�~y�
~���2�gB���Q)G%��-�:Y�i)*L���Z�����������(鐿����/t)���1��,9�,�c���Ƿ��Bdr!#[�V�^?���#�r�r�g�i�/n��@DDDDĠ"""""""�D��θ���>������H0@�
}Ք:Uj[��
�齼7�>�7����(����;�WWIH�e��X�/!D���������/
��;.���1t�Pl��Mg���qf�Ϡ����$�I޳��#3z�hl��UoИ.O`ݹuj�b����&>���o������~�C���}��D}h�=���7��WN��p�@��UQ���T�SwOa��� ""����ta�Q}�󡧋'
�P�!c���W\�����<�9�����6�}u���_��ޫ{p- 7��DL\L�~�޾��[�KwF�\��[2sILn9]���.r·���o��R��KN,�������=����qvpƒNKPz\i��$��?��{[x��!�����������^���/�ļ���߫s��!�>�n;���F�Mj6�߀�!�ADDDDD�cPQ"�+�C�����c����t�D圕Q*K)�W�����bN�ڏ���I�]V�����b�,�a�C���R�꼯����
q�d�E�H����[�3p'&�O����_U��U�Ro�TƽW�>tv)�0��4�(�#^���3h� �q�*˒m�����T<Sq�m6��"h	��ۊf*���z�,������Ҟ&�#�?	}kY�%z���Q�H��s�q�����6�ژ4��
g(���~��+|�t������{g���}�����{�?v��
���vΑ9j�P8cH�L���F�l�0���XD�<*���b�C�q���f��������o��a����@�>��`ՙUX�D3�._�|����#!]	����d��%�/�[pl�X������������l�v��Rc��Ɠ���<��Q�r���n��#�>
TA�O��"�\����k�9�r!����K{�������Ǡ"""""""�&Wo�����%�C��"W�1�.?�����Hp��O#�G6�/ﳵ��xߍ�3/����&�-�f�j
Ʈ�]��$�F�����_�U%gN�NX�-
�x��Q/T����Չ7�p��	ԜZKv���U��+��t���7��o���pP|򼜻NM������_���)������F�ar(�+��9u���d�#W�Te�ޫ=�;���?'���˗/���jL�?;.��8J��ʎ/�)MA�2]����a���j����ѯo��K�Wӿ��j���f4����nWǟ��<�K�؂�
�9z�(��:�'�O^���Rއ�"""""""""""[���l����̑�3�:?E.l�Y��4�`��q�;�B��TྜoҽlwuQ"-~�����o>��������
�b���������Ȇ#�~��J�5��|/Cb^���>Z�����]J;�-G�/W	�P��3�d��տ��xѪh+��iV���V�ޫ{A�ɉ=�;-V(��`  ��IDAT�7Iq�l�lU��&)f���|\��NKP&k��mM5��NK�bN��ŀ�������U�󪮫�������C���#YB��>_�9��<���#e���};���|��?DrL����?>y��ƍ��PW�tvpF��m5���\�rT¾k�,Z^.�\�\��f�<��7)$�9����_`R�I:��n	�밠,u��5�y�u0�Lo���6�N"_�|��E�����9u�F��iU(��h�R����}&�L:�뺸+��\�w�ѱ��;�����u^�y�<9��k��s$������8�!"""""""J@r���E[#)�b�Sj �Q �w�o�8�q���6_��?>4J�'m4/�I���@���Ua'Qr"W}��zz���]���|Ns<�x���#żU'U�B����Q�4.�3��D�%��>5��s�U����4�8�;�m��C3ADDd��/R'�Jp�9	W��������'9	����6?�e�,��YK� -�K��8(F>��E�n0�>4{�)��Р����loS�������f/C����������������#a.��9��7Ǻ��T@̻�d,�a5��]�v���7U�YW��ěGƩ7����u�w
�'W�ƞ�غ�.֚A1DDDDD&`PQ�B�QMF��b5)x�M�j�A�ļ2b�Ud��H�\s�α�(.���F��~���_]�>�(��,:����(9\m0�����mkϮE�ymi�X)S�����]���ԩR#:.����Q�Bn5������֘�z�[�&' �����d����ѯb?��ɯ٧n޺�!""�� ��~(���f��!��84��ː�!�`y��}j�e�2��s�Κ�������!�C7��w�l��m�*��6%���Q3wM���7���V:b^9}�4:,��C��a�S�Wf����|�ݖ����\��vz�i�qL��x���q���� """""�CDDDDDDD� rz�T_�V�Q	I���t\��fWVO,a�a�rݗX�u�UǍ����v�*	j;�-�}v���H*f���^9���_�]��K�_޺mg�N�Cb$�Z�jhR���SьE�h��_c.=���k��������:��{�ײ^pwrG�"-_��s���?h?�������p¾	��r�f�r�ˁ��Ț�����"�E�}Je)'{'�'���gV�a�C�sM��=oڼ*�E>w�C�|d~-c��QA/��se��<��YK�l�P�����zMQ�$�]�wNࣹ}��'��5&4�����7&U�g4,q��u��=
?��!^�\|Oέ\uf������0��X�R��g�?Օ6����b��5��>�Z}�-W��%'� �q>d�]Ơ5�0��L$v���Ϩ��.:-�Oo��C%ſ;.T��W�JN�g77x"�v����+�W!eƒ|Jf.��������쟂헷��/A'2���n���o��\]jA�(�GA<C�m��Mo{V��6/�wvpF~��j��I]�K&y=H�ZXT�?������R'~%..(��(
�P'��9�!�S�xI�QL\�E<SW��d�o<���ޒ�
��L_�2�5տ'���d}��?��7'鐆l�P<sq�x�x��(y|�G<ǵ�������cI*�MN�,��0�˫��^.^걗m��n������gq��$�`:��J X>�|ȝ6��ox:{�� �٫��b��������{fG��E�'m�O�^-[B)�=FГ �~\ %]�ϯGtl�[�oJe�
�3V!!d:�v�1T�2]u��Iι�s��9�o��&ۀ�V�Z���#��
�+  ( DDDDDDDDDDD����]�{�~+������ѽlw�������u���Qg�Π�b��1(������H�!"""""""��2sr���]�7��M6aԞQ�Pɗ��o�����ژs��Ar0��,4*�-
�@RRշ*N|qBf콺D�o�|�
�_�Е6�ڨ�_}$HiF��p�R���hY�%<�=t�	�h;�-�~\��Y�	=_��
�_�@� a�H!y�,����z��z���[�sVF�H�"����c�ŭXyz%֞]���+���S�{-��P�׺:�Y�㷏� ��A��1��!��ɺ�"�e'�Ż]�4z��%;�L�2w	��rq��&9�Il�ӯb?�.��22��I��>�Z�T�X��(�2m��A�**�4$���㋰��:>dMsTD��]t��ܩ�	�%ۄz��{����>�S����$`fR�I:���z���~��MB->��1�j�b������������7���+�
�[kR�	l���v�m���G$7r\q���:Ԓ�3����.}Q��m����NGrv��E��޿Z$ܧF����oDxt8�e����|����"�$�%<���.�Ё�LO`&L���������p��M�q�rT��&�!"""""�0(�������������o�j���A�t_�=I���skq%��*p���'ױ��n$}��U���2ڊRl�tTaD)����ۅ����\МG�w��3���Y�k+�]�x��X���m��¬C�I���C͠���f�2�d,�v�۩���is[4���7ڗh��{����]��PS�Ff��K`\�q*(���R�\�rjPy�Z�m��a��1&�U��iZA���fP��'�V苟���?c�8����$�f��*|!1Hp�7��Q�r�k,�_w+�MM���n0�=���������O�>*,�T2O�b��t5��
�����v�,aGZ�!	�z7(�f��|<
g(l�2t�$�Hk��nPLF���d�چ*�f?y�h-Og"(����.?l�ɕ����dH�A�����zn��\��b�?���]��(��<\]5����Ú�~�1h��t�KhՈ-#@DDDDDDDDDDD	G����}a���\�ά��VSu~/("���z��uLgP�|�KDDDDD�aP��IQ��t~����\�Sy褠wΑ9�@�R��/B��8$&$�c��ER�d�������z`*�>CkU'�����>�>2[���j3K1�#�-�/m�ᛇ���#5	w'wU^(C!�!��ԩR���hг\O��S[�.�?��0t]��ߓ�'z۝�,����&K�B^7c��QAt���ǭ:�����7���v)�`m2~ろUp���*$hmy�娕��E�H�Á����1jϨ���뺯S�K�,�R=���z+H��d�(�ɑG�crk���ŜvsнlwtZ�	7��@B������}25,,�����f����˕c����\�깪�p�K/�V*d��#WE�ux��Ga�����r����5,*̬q+���7��k���� ͠�RYJ��epEDDDDDDDDDDD	#m괚��o6{\9�D.�&|x��{��z���;'u���l�w�DDDDD��b���������(�cl�ML%eRԿ��:$�?��A�OL���V$7��OB��P0}A��'E�rR�����#�EωL�h�c��� z��{�cɎ��0�����0}!1�.l��[�7�d gg�Юx;�.���u�fN}q��{�C��n�w���:H��������-?�O~ؚ,c���h?�=V�Ym�1]]���FT�Y�+���ξ;-XyEC~o�;r�͍~+�����IȐ�J(�5H���%j[7f�X���f���Bil��oUt-�T!^�������V�N�:f͟2���X�4��x����\����.��]3^?	��U��\�%lEv�l��7��Dr���.�����������Z2sIͶg��I��&A1���$����# """"""""""��!�'j������������>��~���L��QrƠ""""""""+Ie�
+���($&�qn?�_/_dt�[���u����xz����r��f���Hn����cs���5��l�8��������VSQ=Wu�Ɲ�|�>��S�A�>�^��ڗ����z��sB���U��t�E�D����Xt|�I����֫I��%�r�К�kТp���(�#�� iK�:�����O�>p�w²���lv3l<�Ѣ�$<B�D��	\Z�m��Bb�$�#a1�$ǡzn�ZH�+���n2Z_L�7�j��U��َb����ҹ�S�Dg6�ޫ{m�	h��q��!1"���3G��mձ�<W�X��Suň.������ 2&����6��h�O;0ə����v��C�+���f�����+���f۱��l"v��!��N�!""""""""""J8Z���=,=��:o��zk���Q��v������?�!"""""""�)��~.j�m��R(6`� �;�N�.��-��ĴV�����V�-$7�.m�((&�Z�M�X�[.n���Q>{y���?�����.>���Sk�[�n�t���إ�������#쾲D�%:�������+A�ZL�Y�/�ݵ��Ɓ�,Z9hɉ%F��{��ѡd|��;�|�_V��*tB��s�}U�7=�|��wN�0�k��!$<!!��1WGWu�.		)���e/�,�Y�g���:.B��%p5�����q��U�!��î�]����>����^D�P�9y���S���P�3FьE��c�����g��{
�oP�-�1y��q��Y=��
5������?��1.=����� �ٯf���M��A�� �In>����(,#�i9�jT���F�#���G��ta���+� ;��D��E��������>�{~�/��ދ�<Hx�L��?u��*�܄r�y��a����=}��Ї8{���F�������z��z��>���T�}�cN�9�!1�X�}\-�዇j;%W,,�S E3Uag�.w���굮+Sw���O,����􃋃��6	��|�������'�O@��G�<�4�%T%&.��q%�/�WN�vٗ�����ն_k��7]^�69.)���
2��O���5"�#ن�zzKm�N�=�;������������~N9�RZc�F����J��{DDDDD�b���������`dÑhW����I��Ā��q�*n~���V�ʣ+���*H�	��w,��헷�z?�=��&g#w�TE�搢�����M^��{���"�E�H����X�m5�O(����7%2�x��V����߻|o��ʡ��ߊ~�ĘC�y%�
ry�R���RYJ��ͣ��j殩�]���`-�����?Xyz%֜]����#��5r�@���T��V��~Mo5����'�����N�}���<�O2u[/���WD�BMмps�I��P%g��ױ�����/��M��lѷb_|W�;�j�5�{����I�2�Q6[�x�K������;�9�x��*�pH�!Te�
6�E�	$):��E�H�����!1�oƯ;��sk����]�����Vs�
��En_�e%J�+e� ����O�>�n������S���Ru�^��_����j�ɚ�2��,8�;�k�zi+�����j��)'�6)�$^ Ltl4f��o�|�s>ٟ�"(F��"��u��_�������<m�����]L�!a\��i��s&�%aT���I�*嬄u�ס�o���$TK��$@x���V=$"""""""""��\�A�7�=4��Z�M����%G�!"""""""�P���e�/M��a�Ct[��o��s��	��2����5���7���/��V��67tG
�3)V��C�غ|��U$���KT��&6��>��R�'����I�\���}���!�ѿR�m�Ϭ�ܣs�d}��X�ᵆ��M��bt��}���	u�v`��SƙC�۝�;�� �h=��3��[+O-��_�/l6y9-
��,D��H��U��9$������l�:y�`P�Ax	��r�U:k�x�M
����~fp_(� ̞1X{v�*0��_g?9�OB=J�+m�������_�_B`��e֜Y�B�ҦN���<�㚍C����^W����[W�]��>^�
2�<3��l�W!��@�B
���ߪ�k��'~В\=�_38���n�w0���'*���m7��@����q�!��Yx|�ζ�f`X�a*��]�����K/�Z�9�:f���Q!�ə3��Ϲ��@�� ���k���T�}bH�z�o>�	[����VparW.[9�瑠-	���A��5z�h<
"""""""""""C��P��1���9��b��������,��=涟���M�ϭ�lv3��m������j�Uѐ%��Գ�Fr%E�R�(���H�Œr2���l3Ӥ��XY���!�}W�U����cT����f,����,7/l�(�T�����[/m��[:Ki�N�[g��%��w�#�k��Q��}T��xa�l����y���'�O`-�.lR�^{?ًl�t�Zc�YA14�l��sCb�%�4y�����[�@���|R^�@ԛ^����)�����Y�g������!1o���ƳcG��A}m��UǺ�#�P_��Z�]B�Ϩo�1��:֚Z+��PI�|Q���r�2��Lu\��Wջ�貺����1�x�y�����sT�r=U����*�K�M�Ø�`�/�}���j�URA��Q���6i�}�l�͑>Mz���d+2�� 4�!M��I0�7��Q���6S�[�8������������������>�!"""""""2�}J{,�[oo��[~j9�,ꂰ�0��G�Fa��i������\�:"&�ٙ{g������n�ɥ�|�f��.R�oja�}p��],� v��&z��;����/Jf)���/�^���#�}��4$�����HL�|�o��K�~/��$�mh�W��������ͣ/k�Α���O��������c�v	���Ua��*���ğ��=3�'I�����R��pfC����t��`�9G� 6.�0e���8��:bu��:�%$D
���Ģ�o�~{��y׳�g*��Ҡ���p����>;�^����_a�ꁰ������	 ��&WS?�Eutň����Mߨ���ܝ�Ѷx[����#9���"Zi����A���	#j�w�}��������Ko��[ي���YF�i���Y�f踰#��?�b���������$E�UrV1i�
t��}MΐpK�b��u��YH���;k�|�|={���y�s�ҹtg��Y~�Y�Zvr"�#���r�"p}�����?�<���N���gy��l��c�5���VN��w!�I�F�@L_P�.E�..6�x�|T�#�}rsr���u_ �������ÐC�I�G��-TH�)2�ɠ��c���}��D/��쇘���9u�F���k��]�K�x|�镰�{��a�ơ�����~Z����S�SB]*d���%z.�;k�Q�����W��w�q��C�������$xH�迪�UCbĶK�p%�
ry�ז�5Zia��?�R~j��K�� l���UV��X�eR�H���M'��6��H�%�~�Yl
��&Ǳ$*�nd;�ϓ�P��p��MQ�Ơ""""""""3��ʉojc�<�����U�)�Rؘ�+̱��*^y���
�e�|R ��ktP���q��e�;��u���������F���A�������k���z��)��v�k�H
���P	�8s��+;4���T�u��1�桙�se����×տԹ�����IA12F��iu�=z��	�p��%��5r�Ht)��@�7�~�A1�7ǳ�gVk����]�%ۉN�:a��aF��qŏ5��]ۧ�I��^ڪBm�%�M5�����L	�z�	m��6y=I���S�G�?t��.��*%2����g��������-��z���#�=D���ޏ����f��Ǿ��E�H�Fo���ڊ��e���|&�}��=�Y�38�9��OO�Q�/�}w�ꤪ*̍�����������������/��ab��pvp6�����ʁ����}x6~l�|�������^U����a����f��`����O0y�v��a֡Y�~y;��2o�~���f_��v��;,���kH
���
�x��XCj1�OOܝ�������K���e����d�'x_H���
��V.^[�leMK���Z^�����D��x��VO�����t���>ܜܬ�"$�`���VO�O�N�B����kctP���VE[i��ٴ0GcI𑮠� ��<}�姖#1L
�d���3�O�ҹM�����c0,M���˫m�.ѱ����_Hnd?�y��ѥtا4|j����s�6�~�5\�]��uqW�}vע�H�>1�CA1��|�$q�ŭ������8�<�b�t��m^�Q-W5�.����Ǘy�wY�Sj��%O�!"""""""2Q��-Ш@#��o��=���($F�qX��V)�����C��"~	^�W��J�@�,s⾉(��z��a����FCdL$���ԩR��{hd�޾Z��I%���������d-�&[Yqj�,�YL�T�}\gP���2�g���F�%��Ln���.���w���������$K-<�?��)R����h�*9�`��V[޲�ˬ^����B�cY_o_5]�jp	k�
l����
���=W�� <�xm5rװ�$d21 �u���V��/��'��s�����ݫ|/|��+���]��fۺs�,�H,�z�����~NN�t�T��B
�r����_�vC�Y�gaW�.��$nv��z�q�㬲}6�b(���b�wP̩��0���9�F퇌%�X2�=:�������6��WC+娄��|g�`4""""""""""""""""J�CDDDDDDDd)��l����_A���R�)c�c����{B"B̚���ۓ�M6cJ��!�W�G�L�Q*K)��˗.V�?v�����Ё��0;N�N�m�n�M�����M~~��&L�8T.1<}�����kRP̥��t�H8ҴV��bNX��-9���c�q���GP6[Y���rU�jP�ғKam��$��
�Х�oU��b�o�ٶ��J���$�)�Z ���-�GVU����#�,k���H�/lFl\�M�1��T�A1�k��f�7ff�;��m���L��J����l��2^?����x�_�m���W����nj��i�c��9CcZ��ћGQ~By�q�ⱞ�?U�Y[�y�f�z�Y�K�����؉�������������������y�������ٍ���sZ��Xk�rˬ�$ԃ��2EJ��sHɠ�7�è~������B?����M����_b���x�DIQdl�[���O��W_�*�F�"�I�ڛlY��>���������&Z�X��$t���fdL�f[F��&-sg�NT�U]g[ろ����[�^DRv �mƽ~@3(F�ԬE�B�8k����
Z�އr��i�����?����2+{,^���}�AB-lM^�'���|�sM�EZ`�	�Ö�J�ivH ����A��ڏ�3��m2���v�ݡ�b��}vm�1+�HCAir�h��P߱�xB�l���cV�γ;�3�����^�zi�Ke�
#�P������������������(�aP���0���W�q8N�=e��#EiƆz$�^�<u�Ԡ�\r�^<B��i���fP�������5�4c�|RtܷB_��3DIѻ!F��\����)R�k�r��Hl�hT��$5!!�w��n�rS�z��d�(��
g(����p��9�Ye�4Ų���}��5jj殉�_�U!xs��U�8I-dG�P$L�$\C�<��r��e�E���>h�s$$_�|���-���fq�b�e�mDbH��1e�Lk5Mg[���
���0��Ľ��M�'&ퟄ�������g��}�#O�<�}�ÂQgzRd-��$L�Y�3؂��N�Z�l�$/C�hR��f����b��aV��MDDDDDDDDDDDDDDDDI�b���������ԩT'���aT�=W�`��x�._�9�
�N�NF�#Ş�#���enP�̻:�"4�a��}\���s��o���b���4���1y�d�G��(�		; �[;R$,A�Ӥ�ז�-�
TJl>�>o��X�I��Ll1}*�A���p���Yn6�l�Q��*,��a-�
��%�ߥ'��]�v�}�Rڡq��j����ᛇ���Vl��GnQA-�����6�9y�f��;�;Z%�A�rl9vv��痀#y�Ck��T�����}��r�!�H`BXx|!~o�����F�*�C��U.[9�cCy?�>2��}��aȆ!��d<	@��{�
W�"a-�gԷ�����͔���`PL,�b�-&.~�py��x�֯��7�k�@T""""""""""R<�=0���ƨ�����Ke)e��o��[������2�!"""""""2���9̨�R��ɪO�~�z���������y��:���bTcevˌ�/��eLP�-B�$������o/R�Ha�|R�ݫ\/4C��\{|���ͫ�`p�Π����cW�.$��is������H`��	�pstC&�LFl�P������{u/lEN����O*h���4s�S��ٚ���gYܳ�+�w����]��T���`�����Q/���ܱ��r�E�����F�ǝg�s�90�������X$P�$d"�$Բ%|q�?�пR�xm�Z�Y��
11V��5�֜Y�����ݏ�8�s�����A��ϒ�{m�X�Ƴ��ͣV_���V������؉���������g�?5�4/ܜA1DDDDDDDDDD�H����~��د��'""""���A1DDDDDDDDFh��A��w-��O����_��JSH�4�'�{f��eP�.=�d���&�¾k����4.�ؤ��WU�QR�����5���`���P^�z��T�Q)��U}�b�ΑHLܑ7�A7����C����\�Ө�ƒ�'�嫇Υ:�-*���u�סƔ8v��o-
���63�Ia	͔@�W�=��泛ccύ�q�1i^)d����jfѱ�8t���\��'�A��ڳH��*��t��JP�-���-A+��������#a8I��Bd���q���H��M=0UgP��Z�+���-�b��#�ж��j�O?8�;	 5�u!a"Oß���S�����p������zn@��e4���圖��o�u0t<eN8����o�ݐ��ن�P�x�x�l/����}'}xCDDDDDDDd�ne��O�\~�����C
�Mq��q�2�e2{��`g�Nпn?�m����WS|��;4*�Ȥ�<i�p	�!JjN�;���k��K`L~��8��ξ;.���*���^3OMju;����V�g*�4�i^�~��i$G�%��2��;틷��5�Zܜܰ��R�[Ҫ!+��fc�2EJ�O$���RX�i	*�h�8v��cF7���7��4	[�	i�)Ɨ �Tv�t�[+�Ė��P���+v��}�k��^D�@bH����q�ս*��]ռps,=���8KvT!C�>
Ď�x�I�K�ƅ����vgm��:C�^��~����������S��L�*�P��� ۑ��[/nE��u��~�P�B6	$"""""""""""""""���A1DDDDDDDDH�U����;1`"�>�ٺDǙ�q%�
�?Y=��=o��%@�1&�A1R���v��[Ǥ����ΠJ��X�UP���k�l��!!pwr�v	����g�n0K��5��]�Wr���K,<�Pm�6�ڌ��u����[N��B?�,�m��l�Q�Z���]GWTح��T`MXtb�b��{4��]�t���
��ʓ*�M�6���O*���)�ѴPS4)��έC�U�q��MX[XTlI�O�;(&����M^F�����}��������\�;e��A1�w��F�H?-3�P�7"s9�;be���o��2ݗt���+m�.����۞�3�͖�u�"��ٖi�_o_�%��O��ʕ+���������	�۳������{""""""""�J�����`�ȘH��o�u1%xC
��G>��p��f�[2sI��>�k��-�bĄ}L�i]�5����P%%���+��&��+��Y�f��j��k��������8u�C������A1�����l����Mg��%;�b�y�̳hY�6��4�!1Q�QXrb�
b��������n�a+� ���2T�U]JwA����$�B	����":-��6Ú\R����/��,��v������]��!����G�4��I`Z�(Ps�r�ʡX�b:�d7���K������__����,�c�~�A����[�jH6��k��@�e( 8�{Q�x���lق�g��l�s�ҤI�:8F�W������ ""2�b���������Z��Q���Z
mɔ���!�Ao+������P������!�e�M�a������2�e2zWGWd��aJj����A������+�_o_\������cЧB�N����%�ay��(3�B"B�����lֲ�ƞ�{@�9w��,�U]Wi��l,֟[�'�O�^��~��"��Z���߃�R;���I8����j�Oi�RYJ��j�����4�iL3m�X�m-�j�m��Ym]��`+N�NHe�J�=":�*��
2���C���%�I����4�)�4�2��,�5<^��(ի\/�0Ds���{k��:�J�W��a���;�G�B�4�HH�'�>��C3d�n��BL\���/��rl)�L-�3(��m��3.%���`̝;W��h�]����x����*4���G����x$#��w�0""J�CDDDDDDD�G�(���Q}�:�lM
��u?Զ�5���_0�C
��窎M6���y7����� E��T�Ĥ��l Jr�=%�c�+�W����W��W���_��~��������̓��h>�9Z�^��4��~`�o}1���2�Β��gVc��hW���voo����/�_�3��~��R��gy��)��t�DB��ʡ��4r�HU�_4cQT�YU|����Ӥ7j,;,��F��'׭�~�����]o���VY�-���P��� �i2h�kQ�5��t�1D���յLW|��[��y-�-�Vs�i���)S��춳ѦX����)�� ��1����q�.9�r�d��7}'^|xd[���$H��������������VTT�͛�7$�111x���egg��b$4F�c^ȼ�)!3DD�|q/@DDDDDDD�Gݼu��'E����ak�oD�D��S.[9�Ǩ��>�b�?c�b\S����+N�09(�V�Z�Oio�} JH8�*(F�(����w������ݿ�n��*��]�2��O㇭?`���3z=�@Z�'T#A���68������{H�OW�������Cg{���1i�$=2y�VE[��M�ˏ.�e[+$Fx�x!1�������j��o�z���ZM5E�R���#���ݝ��}���mI7�����Jf7���C��߳�r��g��d�����0��ӛ�m�~��'�O@�	i�xa�
�{��[�n����ձdG��F�^��+�Ad*ه�l3S�?��07��$�c��iŔ�RR.�~њ}���/ٖ���+1 """""""""��c��-H18��(qm߾O�>�-���"88XM��I��uh̛22�Nm�=Q�cP��Ŭ9���Y��:�!W����W��1�o�O��v)��I������^<}�t�錞GB��1 ( DI���	=��WN�N���o輨�����i5��~����.�	㚍��Zñ��B켼S���=~�_�)��+'�e,��yj�"!�[Fն3p�Q��c�������m�����# �$`�]�adÑ:�����/踠��c��]C���}�d_/_$%�s��!5��2�7W�\޹4�@��7}�;��X���>��h�h���b��i�I�JTl�U�S4SQ؊lg�H`�!�_�۞�'^?z�L=0UgP��]��Π�]���Ux�)�xhj���VFp��/F��� Ǌm����&���f,j���J9+i�����;�-	��'42DDDDDDDDDDDDD�p^�x�cǎ%�j����j�~=�97���*H�U�������������2eJ���A1DDDDDDDD�j�R0o��V !��Ǡ�7��_��1���3f1���t�4�'���b$(c��Q��I���W�A1�$��������J�a�����Kg��`ԜZ뺯C��et����AU�IH�����$<I�-�%��U��[����g�~�'`@���Ig{����Ǯ?p��	�ƕ"q-+O��59�9�L�2H�d!�h��o���kQ+O-��䘯N�:�{t��˔Ǥ�O��7c���ػ����?2!H @(A� �	((ME�HQDDEŵ��E]�u˪k��� XTT�4�]�PB-��>����>a�̄��0I���dfν�N�{�^r���vn����4���?y:T��+�&?�W�ےf�W�󓠘����� Z�WW5��=�>���k�ԻD�"\��ce�	�?d����<�{a�zy��:_�����\�����b�\�`4��q��y�L8(          �g�����ʒ/3�/..Ζ������*W�l�cr�d�|  ��#(     �3�=,��a�i�Z�k��CA�b��>G�Z-U�J=��u{���ďO���Z��9�)��Z+��(xP�E�5v�X�f鞥��q�nlw�}n.9�K��O{���Ѥ���~�>�u���v���Pw�$e�f&��,�r��adƦZ�Dț	�0�@��������!_)P��6p�zZV����(����z������սQw��K\��2��t���m�'�g�s.��ۀ��2צ�vt[��P����VkP�A.��7�o�P�d����+?�+�_�Ug>M�S��:��ݝ�v��w[�S�������5T^L@�?��S�Ӫ��������Y�u����=��Z!��4������s�;3D��         ����S���9�N�����Jpp���S�T�r:L�<>W�D @� (     ��f�Lg��CA�7��QVk;�cm�r�-v�jV�o��m�*T;�2�����ӾN{������#|�c?<�~��)4(�>�[��c�v�rf;]���������n��W�yU�v+���M�=� ���~t� b3xټ��g�?�SW>eǮ�0�y��І|���6(�
y�mnPIa�#�Z��Fw�vhm�m�=��������ym�x�b�n�ƶ7z<(�o��y�0.�������_�Ř ��U2h���z�����6��n�x����ye83�qx��n�1�3@A�y�z��Cy.��oo���C�����l�r��z�e�L@�'m34�~s"��U�Qކ������?��!          ��СC*�RSSm����UW�|ysfx�)9�9 �A1      n���2_˭?�^���t5pҝ�y�f`��#=�^͐��߼�~���ʲ&՛�sO���֣[���f��KV�P��#����h�����2b���Lp̄!t�w����{W�	�mX�X?�� ����m�߯;h�����ϟ��Sw^���F�q�k&��PB��I�����W5�	.��9ll����|��W��m]A�!��D�ۥSI���j�u��=�������<��_��3�s�=��IC��虣=�xS�����٥��{��ά���1�j7�=��Y�9�N�d9�|L�n�V7_|s�:s�=�� }��[_1���6�ۮ%QK�	�{�G�w�.{WO���|���vS)���os�&���m���v�u���i����w����<C�Mhj^��          <�ԩSJI���%Qff��=j�+�����cL�Q���W�n�d����� pn�      �Ѫv�|-g����nT�X]�z^�S�6�h���x��Ŵ����\P�3�}��-�T�S��kY�%A1�Y_��J�v�=]�9��y���~���=���R�J=u����,�S��BC�2��I�H�����q|�`o�b��n��0�3}��SMZ;I(��V���z��g��uq����й��R2Sl1!.e�LX������.���Ԅbَ	+y���z��'<Ҟ	Ÿ���n�g�9[I�I�$8xk�[5q�D��רZ#i5�m�	>ȯÉ���m�+#;��+_��3(Y>\�ˠ�&(&�c���Y@~���1W��s�~�@��zD�d�����lCa\y�����~J�����׏�kU�7�TY�_�|�˘�4          �'==�{�yHMM�%:::W�	�1�19!2�q��;�  ��     p�e͖�Z���b��)��f�vx�pO>��lT�Qo�{���ڰ���Y��ʄ��Kq�[�l-TP��[�����f5�ف�9���)��j�G+�Tv��1�/��ɏ���k���=K�{B����W���Cƻ�77����A��W{�_?�~�������kގy**��R��T�DT�p[w��g��Fw��V|��1;����W>mC�ܙ��;M�������y}��6���yfʺ)j��1���S����J�JJsmm��Z�n����W��7�]D;�����k��������2An�����g�̾�����o_�����i�z���k^s[����OV}"x�9�M�yj���l�fl�!          ��!1�fd:d�_9������R���@��ի+  @ ��     ��	��\��e:3���.��<t�y��e:(����ݍ^i����Q�O��,2�]>G^��=�h�����0(�|1��M8�o��v����/�ߞ�n��6ŧ����PQ\��n�p�Y��A�'$��>]��r�um�k��n~��"�G��1���"Ŕw��ÿPH`�<�B�
v�7]���uێn���p�{�`�V�Z��x���֛ ����I�P+��^��r�C���{]������6��1�|-ܵPW6��e���.�GC?����V�nY����W����S|��[Ŧ�
8�����g��LZ;Iws��v�{s񛺷˽r�9\�_���\�c��
����?h?Gݙ�q����UYuI�K����|�6����sX��y���-ߕ��        �Ad�H��@�ԬPS��� �&N�Sqqq�DEE�>c�	�1�29��,"(     ���U�k��'���n���BK����z��v@�7�m�W��w��}+Uִ��Z5*�8�r���0� Tm ��%�%��'}5��jS���������׈�F��Pۈ��z�T{^9�G�P�O�k`Mi������������$�A��N���m͍����vY7��P]��*;x�0��뛑ߨ[�n�43������ͦo���J�F�տ���v�g���/�Z�Pw}sW���U��_��EA�An�7���&,�B7��a���2�m����4��B���G��56�Ǖ�G���{��G����ڡ��p���q���ƂgL^7Y�^��0*X��G+?p.�������s�i�iԌQ^�l-�=�{���/t�%w��7�O3n��~��Sjfj���yaO�>�u��ΌBn�&����\���,s�)���SFLQ�{乜	-~qދ        %[��̿��X�� ��IMM�%:::W����BBBT�F����"c��w P     �BX����v��¨[�n��1�s?\�ʢ�!55�Q^k��8�p�uz��O"�3�=?�W�n��e�fva�X�\E@Ip4�z��C?��ᬀj�����x��z��g���m��ڀ��]G����[
��.׵�]��E���TO]���`�k�_��u;j큵y��k�z��7\֙s�w�}�����������חÿ<���h_��$z���zo�{��q�%*r�&���w�9\�N<�y;��� ���=2�;�>���7լQ��][s`���m&0����{k�[
�1�W���}��S�OѪ��
��6ެ�}ކ��3����h�;g��P-�]��rBs�ŷ(�?P1'c�IJOҔuSt�e��{��G�jٞe��h�G����s�o7���Fʙ픯3�~׷����i������'ߘ��+j9Ȇ���6w�]���ۮ��������ž/�����W�w/.t�]�
�tO�{�x��U�B�s.o��&�          ʺ��,����yV���Phh��1�1&8�<6�z��
 �T�      �P9�r��;�|\�%"4�������ʪg{=����^���u.�a4fpYҧi�|-g	Vk�mG��ێ%"(&�������qPuG�;N��W�O�v�׆!�_>^o/}�#禰�0�p��]V�b��������*x�	�zu�zo�{.��g�	��ـ<�1�	?o�Y���wYo�q�>�T//xY�,}��[y1��/Pc��
�+�UgBC�D�Q�f}�I�6Л׾iJL �7����m�u"�@�ԫRO��x�#yz���+ә)O0�'��v��fxqY����OOj���y���������1�+�]��/&��au+��P��]N?7���}�k�O����phC�뛰>zd���L���<��cEz�����.�����v�5[h��v ���ߴ���|v���K�]�������e�.cӀ��s��;s�G��������s���bBȾ���ez^�S�ߤ澠Ik')%3��r&�ĜwL V^3�E���^������{h�����.b�v?��@�����v��Ra�
��.��)'�p�Bm��h�̶ޢ}q�\�g~��j4��c�u��m��u��	>{���       ��0�Pk��Vx���!�f���q��}��d  W�N������}ς��Oǘb�dL�L�����FP     ��f����'�/(�q��^���ixS;��,i]��^��gg�K�SYP�r]���|/ogGPLfv����8|�	65}��D-��!�U1���РP=s�3z��6�c���Z�s��$�w�5*����Ѝ�nT�f�]k��8������|.x�	3�֕k�_c��޿:�v��a���Fu�#���<��	���g-߳\{b�(6%ֆ���m�!���juk��m�Ǆ�'hw�n���0a+�v������s����z;��<7��|5ǃ`]�J];�ڼ����y���,���)�����6!Kgj�Vs�k��f�9�~�N��A=��]'��<1Ǟ9�����н�A%�%�
��դ��?�^k�Ѽ���z�=�d��^X=�ߚ�U尿�>����,���m�9S��j�rFL�_���"�ǅ=l�pf�߻	�1a5f2�|�kSL8L���>d�P�L��	�2
�b΍��M��r�_>:o����P�bu�����/��ڙ!�e�L>���{��m`�G�����=כ�
�z.�X6i��ӓ�)��ʫQ�Fk/�?����|U�*T�mo��L朚��`�9ט���UաМ{���:{.       �|1��M?���&W�Pzw̽as�����`{w!�  �����DGG����WHH��1�1&8&'P�F�� �'>�      \�T9_�9��*���\״�F���VP�ۃ�v;���L���׿���ܤ�����������k4Wq(� ?3H�"�A�@IbB�Zd�3�xV�9�mq�-Ǝ�;���'v+:!Z)�)6TÄ �P�Z��ԸZc�dB�2k�,=<�a:�x��E�E��߭;c��k>�&�v�Z�翨�~>��*VҰ��l)��;������ݯ�b�[Vb�'�߯&ݠLg����2f�u����6욫��5�ѴH��mMX�pWFN���Tês�u��ɖ�x��l،'�����5���j�9�7���w��������+(fƦe&�p��o�a0& ./!�!�b�-eBI���zℂ3p����E���?���>6�       ���ܓ}����9���ץ~[̄6_��J���_ �/���R\\�-QQQ��M�Lxxx��<((H �m�      �`��GyGy�U���1��H�g�TV���W6��X�9��p��6[S�MQif���>Q
;�9�	�AId�Z}>�
~���l�WLǜ�v�qg���zqދ�9G�OV~���|J�.��7�K�]�U�W���?��ӆ�&�\~���0n��Tf����x��YzV��|1D�]�6��x��w����~xL�v,��$��|��bad��������+?�'�s��IC���Okl����v�zk�[
���r�ޗ��&'�%�aY����_���|����q����.%�'	        #�?�N���S�i��^ŀ���OtS��O�f���I�����@��k (ݒ��lq"|:8�$cdr�+WN PT��     p�ԩS�Z��_��%l�mD[��h���Uڙ���_��y���!�l�2�ݫ���6�8p�y��*���qf;�dfЮ)& ���wk`ˁn;DJf�f�1K��H�w/�OZV�^]������eLF�O��َ���e�-:�pH�t{�#7�M���P�zX��Ly�)��ګ����|�������1'c�}Bw�9C�/�]���~��O��^\�ݦ�޻L?��Q�k�.r{'RN莯�Џ�(o0���濤_#�;���e.��E���g�?<�.M\3Qc��v�-������(�LX�u_^�g{=��z=�@[�6l�0m=�U8?L8�#���?f
       �3}p�����.��}�����c�
ӯw��K�]����^�o��a�=^  J���T[���s�9�����c�cre���U�|�M P�     �B~?{j ֹ%(Ƹ��]z��T����\�*T;/ۯTYߎ�V=�'Uژ]̠Âj�T?��Y
����|Y�k�-�3̀�ԳqOuo����y<RK��hѮE��ϟ����}��=u�S6 ͕~���s��Z�oe��ϸ�~x̆��q�j\�q�ߓ$��̇�~��o�^���^�����_��]���S��b���z�gl JqHHKP�O��.��~/��s��`�;H��#�������~^��x��JWP&`h��i��O��E޶��Zu����B�p����m�H�v3y�d-ۻ,��(8�Y�WP��+?���|�8�E}��;�g�ԧi�B���/�����?�pfg{��'l8�	��������=má6n����       ���۴��g�޲�<�-�'k��f{,$�L/�}Q���:a
 �	� ���t*..Ζ�����L_�ʕ+��1A2g>
*x�- �A1      .�e��k�
T��h^��G]2J��Stb�J���>dj�O.��#&k�C�}*[���6Cպv��g:\X�B�8�C�T�r�B����*�4ILK��Sm1*T�� ��6Rx�p�<�`��P���ǵ'v�v��,�!W��_�!G9�7�7�\l��\���6R/��v����|�7k�,���']��z�������IG5w�\}��K�*�e<5�)����2mo��h��^V��*6��z��b~f.Բ��zB3}�t��7�}������n�n�x������:�3�t�3�6��HK�,����y��n���:�yzV�=6�Y����~�6��9�aUL`�����Cn��}�3miV����k�_c��
.g�����&��O|/k�u{ܬ;�N��<�t�]_�&jX��ۺ���PZ|��3-��:�+>-^�&�D��}i����5Y�Yn���`B@��ϣڐ�V�Z���w�ϾF��s=smh���l�FS�M�ǘ�Ŝ�9ￗc��
��9O�b΍�+VW׆]���\����^1�u��k�y�\�m9�E        �ӱnG���n���~���5�-���[����z��r �Wذ�x��o˞={r���1�J�*��d�c4�� (     ��)'�\�*�T�D�)��A�As�=<�a�FW4�B�x]�`H�!z���򥁈EU9�������@o���_�u�ғ�H�43�N7Eo����oo�W�Rx�3۩�f�b�l_�_d8�bfK�HQ\j� 0�w��ps�����i&(���ڒÜ�L�)5+մ�G��++�?оw�d޿	�1�&�W$�'�Y�L	S�:�l�I�J5b�1��q����Vpc�����Rf0���^�%"4�ș�Z�j�XI��L�=�>�[[�lՖ#[ι��/���U[���բf�`��{���1��2!5A������)�x�"�Ez%,� �� �9�ڢ�TR��ҿ����q��*-�gsIr �@�ڗ��iIz��`B����-&t�e����_5����6�t��dB�r>����d��%��b�nr��r���a�y�^X=U(_A�A���2�S^N`������o�S�ګ���       ��Ż���w=���\f������������6��3 �+VTbb��▚�jKtt�c����
�1��Ǧ@��Q     ���fЏ���A�fPQ�Z��܎�i�֒��7v�J�&՛�ۑߪ���|Ř+����z�7��)�׮yMu*�)����u֤���M�6(�:�w e���l�2[J
���:[J230~ѮE��TщѶ̉���ĄE�!S��L���V�����C���K�i��	�ۘ�Q�7
        o�դ���M@��m�=��'�k߰_�Ä؛>fb���t��i��{]���̋���L"��� J�ڵk�������[\	>cʙ�2�q~�� |A1      .D'D+?̌еBjٙ���cݎ	A1����>P�O���ӏw�������{���גӧi�"�ӹ~gy������ w   ��{�ܣ@�@�u&�g���         �ӏ��.vY7�Y�>���\��:u����}��;=7�9m;��e}ŀ����-z��+���;fb��W~,g�S ���ׯ���H%Ijj�-�ѹ�N��1��Ǖ+W&D�Q�      �����|/� ��W�b<�ѷY_�|���j�W*�̍�w�U���U&,���Ы_UIԤzM�eZ���ߺvk{��d�Iy�i�q��^� �9   �G�#@�_v��zf        @Yզv;a�+�m��c���~�ai��1����<�3��>Z�~���~��:\���rf���M�j��� _תU+͛7O�N�P����ȑ#�����Phh����N�ȘǦT�VM���'��}�      �p4���ӓU)��9�m_��V�[���ɠ���h�����W%UNHLǺ���l(&Lh����tf��
լ;f�9�K~����S�N�m�o�K�]b�QP�   ���퇫N�:.��S�5y�d         eѥ�.u�z\j���f�Ж���s����9Cb�d&���i?-p���̕am��D0�]t�"##�vN�Sqqq�DEE媯T����$��Ք�+
��     ��Iy�zt���g�R�����}�����<S�B5ͼ}�.������Q��f�9�D��丧�=j�D7L�A�)��u&$�����5�{���^��\^����*   ��G�=�n��%��0         �'�I�\Y��c����8R~���֯ڿJ/����O>�ۦ�f�bʕ+��~@�r�9��v
 |]�^��k�.��e��ɶ8p W����BBBN��T�R�t�L�5l=���     pc����
����e^{��5R���o�mD[}1��8�Fe��VIѪV+�8�G5��@%͕��Ԛ����i������W��i��sԩn'��۷i_��?N�P�cp��u  ���f��έ��-��         |��O���k=�����Y�ܯ�:�ež�z�׺��M��V��5[h��- _��]�j����ZVV����l���:����O���6@&'H&�)����7�b      ��o����Z+���$��{�׬���x�D�9��1��Y|}��

UIe��%�/ѫ_��^��,.�Ҹzc}��j]�����\����K��h�A�A����^/6%V{��
   ��d�3����6L���         �U�6t��ڃ�	�1}���n�~á��c^��1~�x�A1F�z�	�Pb���S111ںu� Lvv����mq�bŊ�Ccr�dr�� �      ��$jI���uQ/MY7�����A1�moS�#@#��TVv�|�y/�}QO�|B~��T�9��G�����h?�!����៫rPe������M{k���m�O�>�
2?�S�N	   �_��m(dDh��z���          ��*�(��U꺬[p�G�a&�2��ܙ�aj���b�
�ۧ�a�sյ��B PR�+WNC���˖- �9y�-�U�p8lXLN�L�*UN��T�^]��b      ���S����^�z�\vX�a�	.�+_!o3�sT�XM7u�bN�ȗ���RSFLQ��vi/1-��jb~��ߩ��x�zRz��jMBCl�Z��Wo��K���pA�B���b����/֌M3����no~��{�o���|��i�M����xP̰v�
�ނ�  ��a�;��t����S��z�ި��N̫������;         PVլT��m��Lg���<�m�{wy��qF��a&���c����\uM�7 �$��C�^�t�j�6ԂI�r:�����%**�:sL��� �5'D�<PZ     ���;�k�%�ι\�z�Jpŧ�{l�=/�
�+�8����6i����|�XI�\�������N�3���%QK�1z����B�g�������uQ/]}��
p-u܄j9H��M֛����c�U��b�a���_�V�Z�l�o���+��S�iτ)]���B�;o�<  �x4��\��)��Wtb�����         �����s%.5�c�]�wq[�+f��x�6Gov��	����aÆ���;�������� ���[rgdd�w�k��c�sfp̙�2&`�ۓ��DP     @f�13_A1&�Ą}|��K�m�_�~*NT�@��_��{]//xY'3N����[:ܢW����ЈB�a���8j������|�ؔX��?2���z[�^���V��!��h��#tŅW���f��ۥ��ڏ��OW}�9�s�l/��;:ݡ�]G��j�8ըTC�u��݋=Ҟ�ه�x�?�����  �o3���7۹         (�*Tt����{��w[�t�Ry�G�p���� %YHH�Z�l�.++�ɘ����X������5S�sOp-55Ֆ���\u�Æ��Ș ��P��ի+ �h���FP     @�Ĵ�|݀4��
�q�9t]��T��;�뙫��moӘ�c4u��b�����GꉞO�I�&�j#Ù�i����oj��-*&��՟�Һvk=��Q�h?�����n�L9�rB36ΰaE��./RpOp�`]��
���v�����;���Ʒ��   |����?�_��"         ��s�������h�g�����.O9�|���� (����O�N4j�(W��A2���JLL��1&TƼ������l���i�5S���r��>�M1A2&P&�qa'�
��     �<�g�۠br.=.�Nu;í5E���]�:���|1۞2b������[��&�����d�o�E����5�Q�R�Pmd������Ϲ�ԡ�C:_L8ͨ���/��>/����V�
�t�e�ْ��e�+s�}�����S;��A5iYi��1A?a�a�Q��Z�j��m�.���7+�� _0��P��9����9F��&/36�   |������6�         ���E�X�#�w��c��m�����\!(@Yvf��+&�"%%�t��)&H�<7%&&F�����DGG�3�oHH�=~Mx�	��Q�����U�re��~L�A1      ���O�c<��I�<��ۼ����j4ӄ�&h\�q�n�w���l��1W'3N�=?u����h|���V蠏K�,�#3��C��+��u�7wi��	zk�[�ya�"�i~n]�w��s����p;k�/1nhs�>_�y����/�z+����#[   �s0�>[�����}K>&          �_|j���CC<Ҿ�$ϝg��8�<%)=���f24�W�L� 8���A�DDD�\ƄX� ���d%&&� ��PSL= ����:}�EEE�Ug����гBdrB��U����@�AP     �9�0�mG��y���\���שQ�F�:�ªZ���(_R%����N[ҳҵ��jm9�E�o�?���8{#:9=�._9�����T;��.
�HM�7Q�ڭuY��<2�Ijf����	}���:uJ�hc�F]�ᕺ�˽z��7�Mlo)i3��q�E
����U�դW���x�� �(V�_��f?�ń5�����n����D
���z��#          �%�%�|��7,�(�Lgf���\���:31��7�)�r��;��r�r
 P8�����c�,���l�Ell��1�s^3�}�_6PR9�N�!2�9fs�cL1A2&P&�q�r��BP     @>�����9�s�9�J�Wt�������dCV|U���5�f������<�fP���͒~�@�v-ҔS���ԵAW�����.*���C�j�Ǔ�k��� �(LP�) �/:1Z�-zM          
�L���OլF3;�[a���m#ں�_h�<�B��Iגғ(  /���?FѨQ�\�&�"11�Z$''��&<Ƅʘ����- ����jKttt�:s̆���cքǘ���c8<<\�˗�.�b      �a��z���T�R�s.;��0}��s����oǯ����~���6�[�ݪ��T�$ۏm���/ק7|�[:ܢ��$���b��O^�u�����P�.{���;             ����Lg��;r6!/E	��\���qgٞe����._7�# ��q8�C(�1�&4&��@���$�8&&F�YYY������\����gǘ�*��3�     ȇ�������7._˿5�--ܹP΂����6׫E�Bn�.|U���L��1$=+]#��=�{�l�gmXJY6��P�AaS��|�Ӹzc��+3�̄�             %�3۩�w�e����4�)���-�Y�x�byR�*u]���FP �:LaJDD����  ��������A&P� �a�7S���s՝"cJ�*Ul�L��>��4 (      ��/�G�=��J��\�Y�f6���9��}?���!�Gg=������΄ܘ}�X�1�;��2�V��C��]��U�Z�b@E}���X�P�3AOq�q            ��h��ͮ�bZP���xe��l9�m���vr4Oj�������	 P��ɸ���e�bLpLll��1�<6��`��:�(�K�
�q8
��1&<����T�^]��#(      ��l/��|��?z�C+�����~����]v���l.��韟.!1g2�C���z��7T�]��J��d�&��x�e?����ݺP�9�tT�^�o            @I�8j�njS���$\w{X�,|��m�>\M�7q[�p�ByZ���._�<) @����:��Q�F��N�mx���c�dL��y���) �g�3sl���ބ=���� (�����     ��pŇ�ut�7Fs���ӔS��펊:���6�K}_�6n�8���U�Fo.~S!�!�{�J��o��}?����V�[�mG��]Ƅ.����_c�URz�             ���9���*W�\����zZ��Mҡ�Cj��W�=���f��:������Ƕ P�9�<�(�y��$$$ؐ�Մǘ�9�	��&55Ֆ���\uAAAjР��7o�6mڸ�.E� (     � 2��������_�|Xp�f�>SW}t��'w�L�����+��
�3k�,=7�9�f/�{A�j���m�WI�}*[��,ӂ��t�R�8�CG��*+;��PӠjum�U�[V��}��؄�̹k����]{c���g�)Lǵ5�tէ            ��lO��>�Z�ֻ4W��5�����~%�%䫽�/�Y�/���X�1N�Iu*�Q��.�"�G
 ����ȡ���ԭ[��2'O�t ���` (���4m߾ݖ�˗k�������A1      4'r�����[:ܒ��[�n����M�>�É�Ϫ3!1_������"��	�m�m6��43����P��բf�&f���v����w��Ɍ��zd�-�����m�k�r����V�����Ճ�?�o6#g�S?����1W�)�{5�5ws�m             J�W|�2(�h�V��_�۾�M��7��Έ�#�ٰ��\f����'�I�\1�m>�Y  UŊmq^����+<�̯��ɥ�;�	ǎ����C��iӦB�"(     ���1{�2�Rx��7! �����kîzw�j_���?��0�|�jR�%�'��w����(_u$�^^�>]��R3��ofz��`;��\����V����2Mo'�mhWo���"��7����             ����S��>���s�b�b�<�F�o�^36Ͱ�����W�O�Ck�~�wt�C=.��v2��zg�;���+&$&>5^  x[@@����mq��t*%%EIII�����������L��	��׌����ot�m��nݺB�!(     ��'ם3�Ԭ;f�\�r�Z�I�&��}q�lPF��ZBn�.|������?5n�8{�ט�s����/)1-�Hm}��+���5M͐����C�5v�X            @ia�s��=FSo��v���ݍ�������nyR��uԣ�뀚Ż  _�p8bKDDD��S�N)99نǘИ����P�dP�deeٰ�|�1�x     PH?������}=p�Z�~X}��mG���/�,29C�U��m�+�\���F� O1�4�am��[Nf�Ԉ)#���.             (M��������-z����$;������V9�.�D-  %��d6'H�nݺ.�IMM=+<Ƅ�$&&��9y����ߋ/��W_-�b      ��ɟ���/W��vŲ=�2o�<ܱ��eeg)%3E5+�T�*uբfui�E�j���_����#�)����L=:�Q-�w��~+rf;��q����i����7�J���|��"�G
             J�S�Ni��QZ��
5���������:�pУm�A�#;�tY�}*�� @�lK�Z�\�gee)))Ɇ�$''��������0���l%ɪU�ԵkW����J�h!      ��������W�F�^ن	��r�����؀�����\��z�k֯D��,߻\sw�UY�p�B-ڵHW4�⼽��IG5���x��D��ʏ�x��=����޵�             �V'RN���}��E�V�c��W_o�Z�vM�kԼfs�u��`�� PV���+,,�W�N��1�1&@&���9ń� ���[�l�%�\"x��     �q���i�C���*�(�Ѷ��n�h"�Gh���8�a��/�=]��=��Qx�p���s�
�s�>�e.;/�^�o�ݗ�����w�����>��cf��z�χ�             ����G]���n�N]�w)R[�N�ҿ��K/�{A����ϻ��vӷ  ��p8T�J[��w������8%''+11�ɘ�9���m׮]��b      <`鞥��n�F]2�cm�٩��w����Ej�`�A>�ڢ�4���z���Z��|��C�m����(&���7���s��w(-+�X�w ��~��G]��:�����(+�t|             e�����>��������U	�R�6v���?>�Y[g��7�Nu;��35�o�^  �`���mq'--͆�$$$��z��I�v��{}W�\9���     �������t�4��!1gJNO�+_�+>п��K�_v�~���V}&�ϧ�>-֠�q���9��?����屠���1��C             P��ɵ^��u����N����]D;���s���h�<NY?E��N��]�_��ۺ��W���  �g�V�Z���t:������8%''��&@&66־fe���Djj�RRRT�bE��1���b      <džk��e�jc�FyC|j����&�����~�K�]��)53US7L�gƦz{��
	��vL0̘�cl'��a���JLKThPh��Z�oe��             ���K��[K޲�Z�jj_��Wo��A�U1��bSb���h��*%3���)�?P������  ����PXX�-���SL�LRR�}���UZ�b���	�     (��nCX�W)R;&8��/��L���/�SW>eg�(�(��������'9=Y?l�A7_|�׶aBUF��	�'�|1��,ڽH�Z*r[ff             �t"���o��d�����   
'88ؖ����'O�T||�r}5�͠�)EB~�a�      xH��l�ڿJ}��)R;S7L-�����,�4�%���͸u�Uk��67r����s���v��o����u���1�#A1+��                ��*V�hK�:u\�gee)))Iqqq���Urr�-�ÿ́ʘ�OA1      �bߊ"�|���uש��5�I�b@�n��B\3:���ʕ�h�&h䴑��a�|��]��܆	�Ys`�                 矿�����li�(���N�S���6<�|�	�1A2&`�<������     ����^���%;o�q�q��@���=��Y���u"J{b��I:��G��U�Vk����j����|��cە���J��
���Û���$                ��s8��d�IMM�29ńʘ��ĉJOOP     �AK��)�b����>����ԩSz~���}b�>��c8���-G���q���<��}*$�0�����ְ[���y��                �����DDD��7A29�1�������!2�)�#�6�      xPzV��휧!��j�u��|��K�?��w�TH`�׶���6��?��鱶���W|(_�9zs��bfo�-                @ّ$�F����ʲ�1&<�ɘPS�c�A2(��     ���.tP̦�M�w-��]�_��Ea�a^���c��<3a��k޿�v��]�u�'ת��                @�����*Hf���v�����'O�`$c�&$$(##C��!(     ��fo���S��+�W�u�NDɗ� �+>�B��J�o�P�!��É���ƌM3��̇�ˊ�����g{�                �_���P�V-5l�P*TP����W��i�dLxLLL����l�LZZ���FP     ��I:�uשS�NZϤPG'F��l�ޤ�����*,8̣m'g$�%�%i����֩��|�ʾ�}�^�3                �	��������7Vpp�U�jU5j�H��???egg�����d�Ή'l�LRR�}nƊ �DP     ���cf��b����._�1z��~�W�РP�����$���Z����t����̐�;�r�P�e�iN�                PL�KVV�-9ʕ+���[�֭k�� ��	�9r�v�ޭ��%$$��>P�      x����K}_��˯��4����Wk����]�*���6S2R�R2��1�C7L�A1'cTĦ�j���VbZ�              (I���T�Y�@�TtT  (�&�ؒ#55ՆƘ�h�"egg��b      � �D�VX�K�]��uҝ��u�v-Ҩ�4���
�q�b 7-�R)�R��{j�SZ��J��'���(p �	d            ���[�n�b�����tf�h�QM>j�Mn9�Em����Bޚ�4U��zZ'44T  ����Z�j�����      /�z��
��+秒��_�~X}��7��m�q�2/���,ݳT�.{W%��0P�����$��6[         ���;����?���� E�}�ZQQ����.W��^�.�k���^[�����jk{���*j�D�wqd	$�$�,��NO������L��p���w��y�O{f&�  �3��%6�id����c�?���a&]�  2�P   �Z2z���;WFvVv��w�����~�n�k��᫵OQ~Q��J
JZ5�zYu�:��hlj�L���Ԫ��M�/j��         �����1���o�o�~+~��c��1���  �eB1    k������G�ƾ�m���y]#S$o֞zש�Sߝ�_i�UާoI���-m����'.M_�%�6n���         h߶�`����w�+����>%����   V�P   �Z4�͑-����GIAIT�VD&(�.���~<}�ӑJ�Vi����*�j[�޲�s�@���}d���K-�^ONy2         ����=�8��8c�q�k7  �j�b    ֢{޺'�t�"/;�E������9��I<��3q��7��=����-�ky�3jMH���uu��
s[��g�=��aY         �9
r
�cnJV��O�:  ���   X��,�'>x"��շ[4�oI�xg�;�I.x����oÒ[�v�>�_��ߟq�����=�����U�GM         d�K�]5q���  �:B1    k��7G�8�E�-���LRQ[>ra�v�m�^ۧ�Ol��V������_i��kP�����_F&�ѥG��Ϊ��~�l         t&sω�'��A��.�%�K�?��q��#+�ժ=�>��x�7��� @gWPPK�,	h	�   ���w��e��7EWf����Lt�;�?����ӆ;�z큃�Y�7?�E��N�O>2�&=6i�ܻ&��M�        ЙL�5)�w���=J>��z[ƶl: ������k�dge����[��*�K �άw��1}���   X˪�V���&�^��ҹ۬�Md�$�q����S�?���6x���:h�Z4��'.�L׿G��}a�        @���^������[ґ�C�>4~���b����uw�8�������� @g֥��/L̈́b    ��;��ӢP̎��9���~id�q���sӟ����ݪuC���֏9���Խ�{��!+��������L�i�M[<w���        @���nI�|sd��8:���q��.����=��q�sפ/� �Y��P   @xg�;-�W�S;��9^��bd��>��������d��I��W<}E�O'�|B����\����l�g�ͫYV�L         ڿƦƸꙫ⽹��}'߷�XLIAI��N�׿t}  tVYYY-%   �&Ϟ��{��;cC1���hL�lB��N�Zw��ƈ�#���)����n��tά�Yq�[�D�K�R�Sߖ�{y��w���!         ����H�s�9�����O���  h!�   �6����xW<}Ed��^�.�����j����q�GƘ��Dgw���}�_�[^�%�5,�L���vo�ܷ�         d��_�>��������c{n�g���3T/  ��	�    ���3�g�&=6Y�ܽ��%%QQ[�hԛ���\����ZwɁ��}��Ʀ��R�T\:��ͽ��ۢ#H��o�W>y%         �<MMMq铗���c��XvVv: s���  ���b    ��S����8m��r�s�-��GG&�^V��q{����[�n����cw86���ߣ�:l��b׍v]鼗>~)>��At�lyH��>9��          3��6.fUΊ>�}���N}w� ��   h#I�%���w��nƆbwL��ա�Ĉo����{8*j+����5���U-�;��Q��e�Ű͇�h����1m��          3555�����;��Ƕ�`�   VN(   ��$W�hhl������Vߎ��ca���D��|-��ߣ��mX�a���ŏ��(:�K�]���t��7�������l�(.(n��$�        @f{z��+�lT�Q   +'   �Fʫ��O߈���ҹ9��׿t}d�$frפ��}/h���{��G���Y��q���h��&�'�>����]On��'�<         d�)��xr�9  `�b    �И�cZ�I���)�I<��C��I�R1򄑱��w�Y�����խW�>qtdge�h���>A�.=�m�j�ܪ�U���         �mA��/.(  `�b    �Н����EQ�$(���{����(y��QRP������tO��k���*'+'F�0:���k񚧧=�I���9�-����X         �m���b��#+��M�  |5�   �6�Y�g1v������?g�s26S�X㦍�#�9b����q��7�F� �����I�Rq���ƾ�m�e5��'�D�+�)�s�yn������        @櫭�]���3u�E��b  ���    ���^��š���=*����O}�蹏�[�PL�]N���8�3;\,f�!#�G{��Uk�h�����钿wߒ�-�;�|F<��3        @��ѥ�
�746Ĳ�e  |=�   �6v���Gyu�W���E�ٹ�����9=2ѫ����{$Q��
"�=x^���\:���ɐ��z�k3_�LW�_�wa�����-���
1         �W}v�zYu   +'   �ƒ73����.n��Sv;%F�-�(2͛��������z/C���s�oI�8i�IQ��&2U�}��a�3��J��g������^�z�h%���         t���^��Us  X9�   �u��箍���-��J��f��EC/�SF��&��|���ؼ�櫽���oG�rD�_2?2Miai����c�������Y#���>�������Ƽ�y        @ǰ��{�����>  `�b    ց��������9�E�O��=qt<���i>��fB1�o��FL8wB�4�xz�ӑ)��d����;�����GCcCL�?-2U׼�q��n��TV���5��U�
         :�!�Y���t  ��	�    �#W?su���Q�[�ҹI\��co���!�,��dM�y�Q�F1v�ظꙫ�G/JEګ��ܸ������.�����kV嬨o��L��G�wl�s�Ͽ��[��
W�        �(�v����������   VN(   `I�W��2���j����֋�'������Ɔ���sMK�9�9?������?��'���ЁC��C��m7�v����#S�h��	;������.�_>��         ��8}��#/;o���:��   VN(   `�ݸ��ɻ��nԢ�C6?�����'����b��=�l@�u�]���Oƅ�\o|�F�k�m�]��[��om��5��ܪ���v�h�����o՚��^�+g         ��E���]����U͋�g�  ��	�    �C�˪��4F�0��k.9�2oJ��8:2���Ek�: =�MW��2��hjj��4t���ɐ�ā��T*���_R�$2M�.=�!������:j���?         Cnvn�s�%%+|��w�Ʀ�   VN(   `=it���i��}[4?���r�-��O�/D{זo��7`��HB:#��&���羿��7�l`��1q܎��V�mkSu]ud����x������Z���G�5�         ��[~�����=�l6�+����  ��P   �:�����uJL��(.(nњ�������^�+�Ο�Y^v^��sP�A����fM���>�|�L<?��(�._�}���|��7⛛~3�;m�S��L�ZJvVv��/�7ܪuɛ����X         ���⠸��k�e�*/}�R���+  ��P   @;0�|F��s��cnn񚲮e1�G�b���׮c1���������>=~�Ϗӱ�|S�M�)��G>��UuUQ��*��-��y]�K^�(�/�^]{�f=7�e�����$��.$�'S\w�uq�և�jM�s9���        ��շ�o��1q�NǷ�bl?{�g  ��P   @;q�k��w��N��-^���:����X��>��hÒ���Je�c/������$���ޥR����1|��Z������t�        �/��΍ny����H_<.� [򙶒����j��b�������:�Zo��g�Z��o�g?z6  ���   hG������l��ܬ�k��I�b�^?4ޙ�N�7�t�$X}�)��"�Y���#���qZ�����_ċ3^         Vl���c��Xt��O���?;  �hhhh)�   �v���<���x���(�����/Z?^<��8�������d��	Vߖ�m���JcSc�7ɕjn;�8v�c[�v��Q1b��         �s��d~�C���2  ����	h)�   �v��9o�I#O�1'��T*��u������>�Ӹ����=�ѥG��g�`�u�����,�Ο�I�.=cԉ�b����^��goƩ�O����         ��^>=�s�wbʼ) �?UWW��P   @;t���Ņ�\�;�w�Z���W}�إ�.qƽgĢ�E�.0��Jek��[S�o?��7�1�=��ؤ�&�^;s��8��âz��        :���}(N��Ԙ[57  �_s���G��P   @;u��WD�.��}/h���v<.�'�:9���t�+���9�osx\�������I������^;�j^p��X         ����qѣ����{  �euuu-%   Ў]�ȅQZP��l}p�_i�;|l��ſ�ŏ_���іv�p��ِ`��g�}b�����缽ΞC��>�@̡[�J�+k+����}         t\/�x!n|�Ƹs��aY   �O(   �kjj�3�=#R�T���i�^��ʊ3���xl\���q���GCcC�m9Y9�ף��~ެ9���a��Q����N~���zJ\��+���t��XX�0��x��7        ��#���G��?�����)O�G>
  `��   h����1�Geme�d�OVi��]z�uG^��}N�xzD����Q�PkKٹ����w�6Gı;�&�j�s0���!���6�i���|��1��bҬI        @�3�~��h/���U.�����]9;>Y�IT-�
Zfi�Ҩ�k��+'ׯ     ��+m������fa\v�e�J�Vi�A�ō߻1.vI\��u�`̧���癗���Ĝ�����#���t�M1s��xa�k�\C6���:p�j�3�|z�aXL�?5         h��~7�|C�1�����h�
7�S��  ��P   @����c��iq�7G��.��φ%��ߺ<.;��7m\��8:���d|���Uگ{a�8n�����46�q�w�˪c^ռ�Mj��Dm}���_%%��ʊ��z�G~N~�k���1���q��+�7O�f�^��[~�8~����gŶl���=7��8�֣��o            V�P   @��k�]�Q�Gq�����/�#	�84=S�M��?�gO��f����Y<'��-Y�&	��-��{��7�=��x�����"��Es��ƄO'��>H�=��'�>Y�hI�.=b����c���6�o�m�]z���+�JNVN�l����=�ǟ_�s���m�ߪ�٥g|k�oő��6�Ѭ	{�oqƘ3���.            X=B1    ����ǎ��1n=��8x���ؾ�zJ���fYM,kX���-�Y��|5�����&Ifm(�.O�w?�K�%�m7�6o28����m��";+;֦���C��s�������x{��1oɼt'��%!�$ԧ�Ol�}�ش禱�;���v��{m�Tj�=�$,t�}g�-��           �?566Fuuu��Ԥ�&#9-%   ��� �!;$��缸���!���0�0=ړ$���{���>/~�b446��s�I�'�<�z�WQZX��/t@:�q������Zo��X�&͚��ql�?��           �� �xkVVV�k}}}��եc0�/�y���g�}�<������b    2X����㯌G�4�������v�����1�8>Ƽ5&y���Q>#ڻE5������G�b��M�	;���t|�EGR�P�?uyz,kX           ������I�$�D`�.]����dɒX�pa̟??�Ν����6	�    t ��y'�ip�5���Ձ������(>��,nx�����[��G�J�>�O>=~��O��]N���J�E�{��g���ώɳ'           d�����ڵk��0I�%	�TWW�{��/Na-Z��� X��b    :��Ɔ��k��	wƥ�.������΍L����c��#b���Q�PIeme\���q�����=��/�e���#2ʹ����G.�{޺'           �=�������t��{���Leee̞=;},��	�    t0�̏3�=#F��wa����-�[d���f�ŏ_��~[465FG��~i:sפ��/G�%������}?�x����;���>           `]KB0.L�� L���ҥK2�P   @5�|F�gx���y���?���1x���^555�/��?t~,^ڹ*�sω#o=2.zQ\r�%�J���I~&c�wL�#�M��y          @[hhh������,Z�(�����***���.���   �ખV�-�ݒg�uF\u�UQ�S�I�����;�-���謒�ʯ��u����%�.�������1w-�(           `M���_���������!��X�ill��b    :�?���x��c�c@ـh�������~�j�뱿��������^�O%�����>��XZ�4           `U|1��_�Lr��Xr?�;���b    :�	�M����s�x�q��G��'�:I$���G<=b��b�,�SF���}_           �ש��I_������2~I�'�9�>�   �N���2�w���ψ��:�s����x��������j]�s��{Ǳ1�|z           й%DMB/��K�5	�|1S__��'   Љ���?����O����ox����r�s��y��y�������.           �����:�I�/�H0����c��e˖|�.]�DG�J���   ��&|6!v���q�a��ɻ�ܦ�2oJ�e;�١��9�rv����#�=           t�����/����ͣ��"�I.<
����0:��hǄb    ��������?��G\���w��mr�n�݂/;~����|wM�+�sF,�^           d�$��^�Lyyy: ��N�%#�/��TZZ��R��hǄb    X����g������#�9b���[[|+^����,Gowt��+	Ü}��1�͑          @��dɒt�%��������R�~���!   ���[57����8r�#�G�1��Yk����ꙫ���"����ٹk�<wN�3�}�ܘW5/           Xwjjjb��GUUU,^�8}{���QWWОm��VA��   `��|o<5����+�=N�T*���ѻ[��������"N���8|����9f�ψ���x���          �����!***bѢE��H0�ǒ L22UQQQ4(hB1    |��ڊ8}��q���5�_�n��?Ǚ{���x<��Cљm�k���\k��,�����*~7�w��nI           �����ӱ�$�R^^UUU��N�%1������j�}������m�    �R/}�R�q���]��|ylP���;�J�m��{^�g|0��ʺ��C�>%%ke��'��?t~|���           ��jjj���"=��/����ɨ���6�`��y睃�#   @�465�-��c��{A���9�-��ٻ{a�xb�1����ӊO�3)�/�Ny �X�{'���=��x��g          �/KB0I ���jy &�����򨭭��
�裏N_@��#   @�,^�8.z좸��k���3�:#
sW{�~�����O���ib1Ih�>{n���w�g���.���{8           :�����񗊊�����OF}}} �STT�w\���#h[B1    ��yU��'�$�~��p���N�.�]Vk�-zoϝ�\�~h|�����zv������L�51.{Y�;���           Yyi�|1�|;��466��4(���oGqqq���b    X-�*g����=zQ����q���cÒWy�Mzl/�����۾�|�LtD�{�G���ؼ��kd�f�W��"z�!�          �è��KG_.\�<���(LUU��P�Z�a�w�m�Ql��ѷo�`��   `�����k��&���8q���o��n��*�Uֵ,�����1��-���ЁC������խ�j�S��:FO���1y��           �4555����ŋ���<I�0��d$��``����^��ѣG����o'���,����C(   �5���6���_�c�~�ǩ����pl��j��������c�M����;+��-�L�J�����<.9����^�}&|6!������	w��<           �U�I�/�h�4�O�0����}�����/�Hb0I��v�;d�    ֚W>y%=��ǹq��ĕ߹2�vo�'�zr�����ߏ�f�����q�17Ő͆����@\��%�P          @{��L2-Z���$c���QWW@�XQf��֋^�zEAAA�1�    ��-�[7�zS�5��x�'����U��E�t�Kq�s��=�_Q��:2AV*+��9<�8�(�/Z�}F�92Nyb446          @[hhh���ʨ��Jm�����oWTTDccc m#'''�����=z�C0�Q�$���t|B1    ���g��p`<q����dgeǏ��q��q���=o�MMM�^��o����]6�e��5q�H          �������ŋ�ї$��D`���ǒ���3��.��$#��$Q��۩T*�܄b    hS��|-������>������{�N�+^��B�������/E{2�l@\|��q�N'���7�rc�>�t�          ��jjj���*~i�$�d$ǒǄ`�meggGqqq:��`��Ks�gϞ����u�b    hso~�f�}����i���/�b�&��ų_���>�?uy��6.֥�e����<N�����Z��ݮx������          �P�i�4a��'a���� �^NNN-�����+=��%%%������b    X'�Ο��48�?��ح�n�����O��g�7�|C��8*/]m!+��6g>+�����U�X������^�.          �Ω��!����%��hѢ��d̟??���X7
���QZZ���4�N�Rk�P    �����1�/C��cn�cv8f���e�]���C���ߺ;�|_��:6j��Ě��X��F��w��n��ѱq����ދj�1�OLy"          ��+	�TVV�0UUU��I���<}���"X7������8~I0I��9
SVVyyy�P    �Tr9���b�g�7�&r�V�%�n����� =��U��)c�ُ��W?y5�������Je�������{�77�f�;`��[�7ִ�f�G�vtL�7%          ��V__�/NG_��K�I�7K�755��.��$#��$Q���Ʌf���   `�K����xi�K1򄑱aɆkd�.�]�ЭM�D}c}L/��,�$>Y�I̭�u�u��n�?��u�����^�=zu���ŀ��ck�M��g�wV:�          d�����>}z̜93����HG`jkkX���KIII:���/�`�QPP�i�b    h7���\ls�6q�!W�i{������ʉ�eӣ=�W5/~t�b�[c          ���/��ҥKX7���_��In'����쀎D(   �veQ͢~��7m\\s�5�^�z����=q�g�ܪ�          d�����뮻b����}ݺu[a&]�v�L�b    h�FO��x\2�8s�3#;�cT�?\�a�������H           ����!F��q kFvvv/����.��E^^^ �$   @���fQ�s�9q�+7Ư�U���J�"-�^�}�q��Em}m           ���G��UPPP���4`��0�ג����]hkB1    �{�gO��n=*��}:s�ևe̋�kƟ��S\�����          ��f͚o��F +VXX�/!������ �O(   ��1i֤8�#b�w��� �����ɏ�hʼ)q��7��⥋          �lcǎ������*'''|I�/��b&��<�]�+    ��ٛq��FIAI��aq��'����T*�N�WEmE<��q���SӞ�&          t.��ӧtt�����K���1�u��}��b    �XI�%��$c����c�?&����o����k���iŧ1n�x��G�o�#j�k          �X&O��B�tYYYQRR�<�D`�C0�������   �Cx����WO�*=��u�o��F�;`����ؼ��ѫ[��>G]C]|�ࣘ8kb��p|:3u��           :��3gd����(**Z�)--]��ݻw�q 3��   �gIݒx���ӣY���1���X606�i:&���%��u���Xְ,��VŢ�EQ]W��g��9���ySc�����          @�2k֬���!��L��]��1	�    �),�Y�~�jz           �TSSS��������(..^�)--]�)++���� :�               �
uuu�����.��$1�� L�5�ĤR� �"�               �
"1��/�`����իW@k�                �����t�%��$�$��Ib0������                |������d$1�$
�|;�J@[�               :����())I�_� Li��$�

�=�               :����(**�R�w��ѳg�t,���               2^aaa:��<�L�i��J� �	�                �^vvv��/I &��4Ga���"/// :2�               �](,,\IF�I�0ͷS�T tVB1               @���1�޽{GYYY:SPP ��P               |�����urss�ї�Lr���t����� ���b               �+����&��*,,\�IFs��v*�
 �,�               �]�v�����L�8N|�b�9����� �m	�               ���h���wމ�&'''�����޽{GYY��LIIIdee �P               |����gd(&�J-�$��L�����  s�               ���n��b�رQ[[�Mvvv/�����.�����E^^^ �1�               ��Hb+{�G�?~���K�.��/I拷���"�J �P               ���{�|�A̞={�������������FAAA �P               �Dvvv�p�	q��ǜ9sZ�>'''����% ���ݻw�q �:��               Z�k׮q�)��s�=���j,]��_OB0I &	�4�`�o'k`u�               @���������o̙3'#???���� X[�b               ������O�> mE(                ���                h�b                 �9�                �vN(                ���                h�b                 �9�             ����݆Jv���3�qf�I�E��Z��(V�|�����Kɦ.jC[(�鋢/��R�j�m��aq�!�I��c6�4�<h�n��&1���n��y�Ng.�U�Iv����|��̙��������  '                �8�                ��	�                 $N(                 qB1                 ��                H�P                @�b                 '                �8�                ��	�                 $N(                 qB1                 ��                H�P                @�b                 '                �8�                ��<�~����U*��fB1                @)�������3��2�z=��P                P
�f3:�Nt�ݟ\˲,VVVvb1�L(                �6�Y����/V*��ꪫ�ӧO/���׆�)��߿���ػ܄�~3&                L�޻���/��                �M妛n���q��T���j�����{�ޓY���Ї>�dL�                `������O]�����#��N�V�0<��Z�~�^��:�~���~$F(                �9��`4�^��×���q�R�7�x��z��sssy�С�F�b                 ~���g����8���7�x����ڿ����ַnM�{	�                 <��`?��|tcc��o����]s�52�`�P                �elooׇ��'O�<t��я>|���r}�              (�,ˢV�E�� 0M���n��� R��t�/\��w7�t�\}��o>p���^�+              %2
�,..���\  L�Q,fcc#��~�f�Y]]}��;>v���߾�뾵�k
�              @IT*�h4��y  L�Z��f3���v�1)���j�z��;��믿���\K(              J ˲X^^� J��=�ŋ���G�z�^����w=z��>|�n�#              %����J%  �f�YZZډŤ���W�����[^~�����XC(              ��h����\  �U�Z݉����HU��i\�x�߆�oߍ��b              `ʍ6M�b1  eV�ՒŌ�������㯻����B1              0�F� ����<R7bss���o��B1              0劢  Ұ���;��rK�����q�+              S��� @�M�=O��˷���hx���W(              ��h��`0�<� �����O·�=[����Xů�z�������P�������              ~���f,-- @moo��~J��n��K/�9��߿���s�t:������t��_��B1              P����z=j�Z  �I�ߏ�����̑#GF�ύƱc�^1�'��J��K�E�3~�(>�|�G�R�槯]�~�8��9#�{�śo���~���cL�b              �$���byyY, (�Qxeuu�Yc.����lxx��������U�^��N'�<����q�+              %1�@=�H]��c~~>�Uۉ��4
�loo����K��������xx�K��F�`?��?�y              (�N��3�,�J��s ����`0�c��xOL�����O(              ��]���=̖z�~㇣�U��3�.��'.<�����CO= �������Ȋq�{���`0����
�E�+�O(              ��[�[�5�-�v|�?���iT��]�i�����=(�[/���q$���Lj�,���s>�                �����EQ\��/|a��|��8��                J���?\�T&���������8��                J��}���o��3<�Ob��(�b                 �O�e�m��������
׌k"�                ���ĄB1Y��b\s	�                 �Uř,�&��Ҹ��                J+˲��Z;���q�%                ���I-\�Ҹ��                J+˲��(&��P                ��E�>���b                 .g�ɲl"k��                ��<��s0�ᄖ�Ѹ&�                J������S1�b                 '                �8�                ��	�                 $N(                 qB1                 ��                H�P                @�b                 '                �8�                ��	�                 $N(               1�۫����W `D(               1�A7y�xU�U 0"              ���|�3���D  ��               $��7��o�!^}ի @(               A�A/����/}�K�\h 0ۄb               uv�l���;����xY�e �.�              ��=r�����g���x�k�Y� 0{�b               ��ߊC�z(^������q�+����zt����  �O(              `J<p�8�/#˲X�.�Fw��l�ڈ��RL�(t \�              �)Sŋ�Č��Vw 0��b                 '                �8�                ��	�                 $N(   �	sO�E  �H�NU7�         �l�   J��F4��  �\ν�\���          �B1   @��?6��Db            ��&   �V�b5Zw�"�             �jB1   @)�<�w�#�f            0�b   ��)"Z_mEuͣ            ��   J�y_3��            ���   Je��B,�Z            �2�   J�v�+��            @��    ��o���r;�^             e#   L��Ȣ}W;*�             (#�   `���ھ���            @Y	�    Sm��K���b             ��P   0��O֣���             (;�   `*U�+�>юl�            @�	�    S'�g;��|+            �Y    L��{V�v�             �B(   �*�'�c��            0K�b   ��1wf.�6            `��    S��Z��]��"             f�P   ����E��v��<             f�P   ��"���VT��            �]vX   Ik<؈��            �,�   �5��|4N6            `�	�    I�=U��ݭ             @(   HP�ɣug+�^             �    �D�N����            �%v\   I�w���{b.             �B1   @2��K��            ��%   $�v�+��             �$   L\��G��vd�,             x&�   `��"��W�Q٨             �N(   ��}����z             �܄b   ��Y:���Y             ��P   0�s�h��             .O(   �s��J�O�#d            ��	�    {*�g;��|;             ^�   `O�ܽ��             ���   �L�d#Y             ^�   `O̝��ƃ�             ���   v]�b5Zw�"�             �%�   vU�͢}�y7             ^�   `�������G             W�.-   `�4l����            ���   v����|r9             �rB1   ��՞�E��V             0B1   �X��y��lG��            ���   �&+�h�hEe�             ��P   06ͯ7c��\             0^B1   �X,~o1���             ��P   p��?�Ǿ��             ��   ��T�*�:ъl�             �C(   xɲ~�;ZQ٬             �G(   x��}m_���            ��%   �$˧�c�            ���   ^���sѼ�             ��b��Y��۠�fw3  �r��W�����?             �#B1Dc�y��[o�� ���zY��hG���H            ��$   �`+w�D��Z             ���b   ����F,<�             �=�v�������J����;q��  �|���	�             0B1����?o�շ\�3��?��   ʥz�+w�D            ���    �)��Ѿ�y7             &G(   xvED뫭��y|             0ivz   Ϫy3��             &O(   x�������              B1   �Ϩ]��ʽ+            @:�b�sk�b��p��E?ή�  `z�[y��܎��             ��!���0;�O  �Tʊ,�w���Q	             �"   �h�ی��z             ��    �^���,             i�  �W�ͯ7            �t	�   ���W�}��              �%   3*�gѾ��V             �M(   f��=+Q�Q-             H�P   ̠��Y���/             �A(   f��ٹh>�             ��P   ̐�j5Z'ZE             0E�b   `Fd�,�w�#��            �t�  �Ѻ�է=
             �Fv�  �h<؈�G�            ��$   %7
�4j             �K(   J�z��{Z            �t�  ���;y��hG��            ��&   %���KQ]�?            @�-   e5             JB(                 qB1                 ��                H�P                @�b                 '                �8�                ��	�                 $N(                 qB1                 ��          `O->���� ��Yg�w6   ��	�           ���AY/ `����   0-�b                 '                �8�                ��	�                 $N(                 qB1                 ��                H�P                @�b                 '                �8�                ��	�                 $N(                 qB1                 ��                H�P                @�b                 '                �8�                ��	�                 $N(        ��c�nB��������ή%K��H��đ�(k�"BsU�Cq��=de�=$��D/S��Ň
���KC_�\�^JEӀc� e�4���tf��M��2�������`��{����
       HN(                 9�                ��b                 ��                HN(                 9�                ��b                 ��                HN(                 9�                ��b                 ��                HN(                 9�                ��b                 ��                HN(                 9�                ��b                 ��                HN(                 9�                ��b                 ��                HN(                 9�                ��b                 ��                HN(                 9�                ��b                 ��                HN(                 9�                ��b                 ��                HN(                 9�                ��b                 ��                HN(                 9�                ��b                 ��                HN(                 9�                ��b                 ��                HN(                 9�                ��b                 ��                HN(                 9�                ��b                 ��                HN(                 9�                ��b                 ��                HN(                 9�                ��b                 ��                HN(                 9�                ��b                 ��                HN(                 9�                ��b                 ��                HN(                 9�                ��b                 ��                HN(                 9�                ��b                 ��a�������Z���<�������7�                ��P{n߽?i�$�Amw����                `��b                 ��                HN(                 9�                ��b                 ��                HN(                 9�                ��b                 ��                HN(                 9�                ��b                 ��                HN(                 9�                ��b                 ��                HN(                 9�                ��b                 ��                HN(                 9�                ��b                 ��                HN(                 9�                ��b                 ��                HN(                 9�                ��b                 ��                HN(                 9�                ��b                 ��                HN(                 9�                ��b                 ��                HN(                 9�                ��b                 ��                HN(                 9�                ��b                 ��                HN(                 9�                ��b                 ��                HN(                 9�                ��b                 ��                HN(                 9�                ��b�Wt�ƍ��؈y����V�w ��c               0W�b�W��K/�͛7���b�                sG(                 9�                ��b                 ��                HN(                 9�                ��b                 ��                Hn�C1�$��fp�х��=Z{4���1�~��A��               `��:���_�����<����{��sq��.�4�¿|!ֻ�               �_s�                �B1                 �	�                 $7ס�����(6�{vvv�}O76�����                �0�:��v�����z�������?�eY               ��1ס                �i                 ��P              ����X,c����ȮSvb�� ���              �O՟��4?���cii)���c|{����_ ��	�               $�TY�k���#�G"� �!�              ��N�N����(zE  �K(               ����qu�j}� �wB1               	U�j�-�E1� �b               R�P���  #B1               	]�] ���b               �9T��� p�P              @2ã  �	�                 $'                ��P                @rB1                 �	�                 $'                ��P                @rB1                 �	�                 $'                ��P                @rB1                 ��u(������NpO��Ȯ��zn              �}{뭷��T*�LbvY�߻r��gǱ�\�b�׷������S�Nd����nM�s;               �!)��ceY>1���k���                 ��(�VY��=��=���b                ��U�ek���b                 ~��(ZeYNj�P�8|���X�S�˸2< ���7{7c���v                �`0x�(������Zs��տ��~����v���               ��(��㓚]����֚�P                0�>:��EQ��ZB1                �,;1��eY~\k	�                 3�wީw:�G'5�(
�                ��O�����bR�+���k-�                `&�ߜ��λ���q-&                ̪���_ׯ_�k1�              H��c��S/�Տbx�"�Z5v��4�T�S��_ f�����?��w/_�����CeY�����8�             ��j��h�����(�V�E�R�;�B �+�hY�1���G���y���Rr��o�\L(�*E%Z��G�����             ��(����z=  f�(s����v���nܸ�k��bB����q�'�S�P�R})��Vgk��             �t�V�����J%  f��w�v��w���o�}�,˿^6�y/��`��1:G�#�^o�z���?���F����l�              �EQ��  3��l�YF�_�7��d����������G���r?��A�0���0�U�V�'N܈1�             �0�8- ̺����t:?��������W��v���Y__����<l��ѥK�vc��b              `�E�z=  f����v����k����{�0T���a�k
�              ���V�{�� �A�V��w��^o!���믎{M�~�V�              �g� ��J%2k4뫫��4�u�b�s��/�W~�+             ��)�2  �E�w�F��W��P̜���+�^�/�ޗ�ZQ�             �F�~?  �E�w�Z�����O��A�=ס��}�s�x���J��F+����N�����#��ŧ�:��|L����ע�o             ��h��`0��3 0��nd�l6��g�9���P��G����g�����z��`��̙x�'���0MN-��g�>�l��             �ص��h�Z 0�F��N�---}cmm�/j����oeY���N̺�G����J,//              �cww7�V� ����ގ�Z��?^�z��/�������j5�|��8s�LE              ̞����&�` �,)�2677���E&������߭��=w�ڵ�5ס�^��~?fݱc�����/U��S�ܖ�             �h�(3
�4�8th�� 3`��t:�n���u2�k��������e^̱;�w���N̪j�+++q�ܹ��̂�?�w�L�s�Lw�            ��F��G�h�i�R�� �J�H���hii�G�z�����>��s��eǏ��/Ƒ#G             ��T�e���t �qi4�V���7o�|�����b#3c��j���Ĺs�               `��������F�O����$�A(f�?~<.^�G�	                ���j�~���^����^xᯋ�('y?B13�Z����s�Qr����?�3���&�$K���Tp��A*��b�Z�U+R����ފ�zzN�p@���{�-�
�E�mk�c-�F�X�AE
Jи���������|=��Ͳ	I�a^�9�3�������a~	�컻;���b�*                ��K͎���ʾ�ɾ��b��١���]}��Si��o~�bD��害�3zzz���#                ��r������XX?��o
�T���&j��ľ��|>�Ծk�---��v��o\~��b	�Y��}Ѣ��;����"                4�\.7��w���h B1�Pggg���DGGG                 +�P�2��磻�;���R�(                �A����p�\����]�v'&&���:::&�>����z�\.��e�}8�(��e���3zzzb�/                ����r�k�}qjj*�P(Ě5k�k���1<<�֭{����7B1�|>�����Օ�C                �-a���g]����, �\-�O� :;;���':::                �_�\�wM(�C*��GwwwtuuE.�                ��j��Z[�b��c�9&�?�����                �D(f�������]]]���                �N(f	��쌞�����                �g�YD�|>������+r�\                 �E(f�tvvFOOOttt                �|�b��|>�������\.                 ��P����===���                 %s���������r                p �b������鉎��                 8B1�I>��������\.                 K(�0��쌞�����                ��K(�*
�m۶8��3#��                �� s�tvvFOOOttt                ���С����=��y�G�P�W��Uq��gG.����ݻ��}��j               p@:S)Wb�<~Я?������}lܸ1�#�\.����߷K�P               p�:s������/�W�����                 ��P�ڲeK��/�rlܸ1                 ����<5�T�s��m.4��^����DSSS �cd�����U�=                DC�b�y���ΉO^��8�� ׽�{���               �H:�\Z����?�=���o�                �b�ُ�O8;n��8��                 XLB1s��rq��F��                 XlB1s��j�w�i��7�"~�����㘵�                �b�����h���o�u\}����all�                 G�P���ǲ`�����wo��                 8��b�De"               `ll,}�ј���|>�~��X�n]�r� �CM(               htt4n��������Zm�z=s�QGe�4�~���9 �`�               �Ƨ>����j�{���f.�bq& ���Q�t��� �"               ϡ\.?g$f!J�R6}}}��ZZZ���O
ɤ�L>� �P               <��o��yGb�K���ڵ+�g��r�nݺg�c��)���&               ��;v,�g��j188�ͣ�>:k=�b����蘉ɤ��`y�              �y�HL�R���T*e���7k-��g���I�z@�>�����'               �����Z��޽{��K�X|F8&Ee�1�t�����'               ���닕�T*e3�����2���c�������!               �Q�Tbbb"U�\�]�ve3�b���xLggglذ!�ʴ�� ��P               �G#Gb�T*e���7k��Iј4Oʴ��G.� ��C1m��hijY��5�5,�b��-˻885�Z-              X��^���/"���XL=$���1�ٰaC��,� �(:s�����N_��M�6����rE\��Xή��U145              ,}�\.8���jd���;k�X,΄cҤ�L
�ԏ�wQC�b               `>�$��T*e���7k�P(�ڵk�hL�ǤpL=(��ٙ��D�v               ��J������Z/�Y4f�ƍ��#2)*��� ˕P               �b�J�l���f��#2�����2��\. KUC�bF�Gb4?���,����]�}�Uk�              `yYY�����hooϢ1)��1��̆���% SC�b&�)��,�J���M�Z-              ���Z����@6����֋��L8&M
ɤ�L�XT8�:               ����T*e���7k�P(�ڵk�hL�ǤpL=(��ٙ�<_�&               x*�Jd���;k=Ed6n�8+"��[[[`!�b               `?��|��522��\�իW�d�s= ��S`&��@"               ���Ғ�b��j��0>>��Ν;g���^{{�L<&�d�q�6d�O�q�               �<���bxx8�HK�����lz{{�����b�ڵ3��\�ȤI�[`e�              �y{�B1,9�Z-�^��Y(��L���c2��Lggg�,/�Z               ��	'�?�p�rR�Tb`` ����g�555e�4)"S�ԏW�Z��#               �8�3���o�Z��LOOG6ώ�$�bq&���A�t���8�b               `���q�)���?�J�R6}}}��
��L@��y��u��pw              �s�袋�G�j���*�J�޽;����g�c:::f�2�8��pp�b               �9lܸ1�;Ｘ��;ؿR��M__߬����g�c��i֭[MMM�P               ,@OOO�ٳ'~��p�&&&��'������|���cRD��I�����b               `r�\��o�"w�uW �N�Z����l�R,g"2i���q�?a��              �J1��.�(^���׿��x��ǣV�px�J�l���f�
�,��1i��I��&              �:����+����������3344�M�Z �_�R�ݻwg�l)�v��g�d�q��X,,B1               p�����E/zќk)^122������٤�t-Eej�Z �O�ǆ���y���g�
���Lggglذa&&�nݺhjj
X*�b               �0H��H�u��Y��j5�W�xLz��cRH&f����T �O
:�{/Moo�3���|���g�p��ttt���G}t�Z�*�H�              �E�"�����J���E��I�t�w�ޘ����H1��Ed�b�8s�I!����r��CI(               ���H�y��9�SH��������,j��Ӥ�Z�����4}}}��R���=�ƤxL
�ԃ26l�����%               �T=$�q��غu��J��cR<&�dRT&M:Nׄd��V��=����w�z�o��4)$��2�s��P               �P�Ba&<1WH&�,���gb2�xL
ɤkCCCQ.�8�J�R6}}}���}�v������"PO�Ȭ[�.�����$               *��gA�4�7o�sO�Y�#2���ψʤ����D �N�R���~��g��{���=�ƤxL���cPG}t�Z�*X��b               ��*���/$���xL
�f��Z�t^��x����LD���w�z�W��4)$��2��\.,_B1               �A+
3Q��[��ZzHftt4����xL�ʤkCCC1==��W*����뛵��յk�f�j�ǤpL��ݸqc477K[C�bR%ijjj���?>��:��              X\O��%�����LL&M
ɤ�4{��r����{���w�z�X��WӤ�L
��w�rd5t(ft`4��b�R	X\�8W�lY3             ��|>�}�4�7o��^��btt4�]��I�������d �O�T�f���ߴiS�~��q�YgEKKK�8:               ,m�\n&$s�q�͹'�-�
�ԟ���8xO>�d6��ַ�~��/|ap�	�                �Z�X�fӦMs�W*�92������j�ott4>��ĥ�^�����%               �h�B!6lؐ���J�����fϞ=Q.��,���/})֬Y��zjp�4t(��o�ڦ��?T�_�� σ�c���X�&�=              ���X,f�y��9�GGG�x����̤����	�GL�H�����w�������y��hDu���T�����~"��z"               ��5k�ds�q�͹�B1�x�ӟ��)4+I�T��۷ǥ�^�               8Z[[�9�c�\�V�1<<�c����@����ώSPfzz:`9ٱcG\p����~B1                �Y>�����g3�Z��dR0&�c��)&S�J���� �w���8��s��O(               `��r�X�n]6���{J�R��B2)��ӌ��dG�#�<"s��                ,�b1��)��Y<�>CCC3��S`�V�J;w�̾W)v����9��!               ����Dggg6s�V�1<<�c����@������xjj*�@�@���x����
��%L(               ����X�~}6�S*���L}RT&Ed��޽{crr2��VJ(�V�5�&               @�X,f�y��9����bhh(���q�<�fh<�r9V�                �����l���T*122������٤�t-ej�Z N(               �C�P(����ٺu��j����31�z<&�dҵ���(���&               ����c�ڵ�l޼y�=�Ri&"3::���L
�LLL4"�                ��b���|!�z@&�c��L:O��k�Z�J#               ��Q�lܸ1�n�:k�R�d���IA����,��2����PLOO,7B1                ��B!֯_��\���lOSSS�)�JYXfll,���ٳ'��r�R#               @�H!���Y�&6l�g�qF���D{{{�j�,$SȤ�����#M(               ��W�¤I��ڢX,ƪU����#�?����r��磩�)�_.�cll,ɤI�ݻw���`���P                ,@��T*����Y�fM6�7o���B2���D�ٳ'{�,$�"4),355p��b                �I1�j��777Ǳ���ӥ`���x|��_���逅h�P�%�^[�[���Mg���=��x�֗�rv�c����d               И��b6�\.`�:s�Qg���N_��M�7��Ni?%~~���rv�On�               HC�b              �Hj�j���z͚��   �              8BN�{j?|�����=  ��C1ӵ阞�^��Z���J��ܷKQ-�]               ���������_�fM �k||<��~�.E��j                ���                 ,B1                ���b���,�P                ,��7
Ű`B1                �V�^�PB1                ���b�B	�                �"��r%                ��	�                 ,qB1                 K�P -ߔ��� N<��lֵ���ͫc�Q���?1��RLLM���P���c��c���S�O               �0B1 ,H[K[��/��oyy6��u�IG����z���x詇������|;{~���2]	               ���b د�Go��N�(.{�e���B��[�{�n^/{�˲y���Ȯ�x̿��_�~1��_��C;               ��YN�<-��į��W�P̑��1����lj�Zܷ�����-�y2               �Q	� Ŏ,����+�E,�\.�mٖ͇/�p������������(W�               �D(���t�I��s��<��Y,f�*4�/zm6�Fv�_��W��>{��               4���m˶���k�ug�.�M�XN�Y{L|�>��yo|��?7~��x���               ��L(�������揳@L.�;��"  ��IDATd����S��ȓ129��R���c�2���Y�&���Ѿ�=֮Z[:�dמ������s+�>�������ߟe�               V"��p�Q'���旽9�M��z�������ߏ��}/���w��]�����ӡ��De�ޫ��=�[w\����8��3�%Ǿ$��:Oˢ2�%��s���U��*�򮿌����               ��D(`+6����k_}m�Z�c屸����w�����1]�>$�kxb8�x0��|����\/4�ksW\t�Eq�)�y'�����������g�3>t����w}��}^               XlB1 +��_��cq�Q'.�5;�v��������}|��oFe�GR����y_67l�!V7���O�8^����/�u���=�Z}T�s��g�������w               �;���ӿ��xK�[�w�4��������{~|O�j�X*Ƨ���|>��|K\x����f�U�U���Ύ{�����/�7>���               ,gB1 +ж-۞s�};�9>���Xy,��r�_}��t;�]o�w���q�g��5��|��/               X�b He����s�����=�X�K�Y�&�E'_��?�O�0               `��h �j9���?���XI������柍��������Z��               +�P�
V����|�o�ۯ�'����������o��������\���               ����C1��R�O�/x����X\����߿��vI��?�����{��O|?�O>��ͥq�	�č��               �4t(�<Q�����/�J,����Y�}�$�P��n}]<��C���~������sqʆS               ���� �T�����j���               �;�                �%��C1C��X�[���c�������XΪ�               P���s��C1�T�����%�}`�|������7               �����j�P                ,�R��PB1 +X���Ľ?�7ƧT�               ��]�v,�P�
�+]������Ͻ=���;              ��cjj*`��b V���:)�����o}"~�~/Ƨ�               X^�b @.��w���������^w=zW                ˇP@���&��k{|�Ώ������L               ��	� 4�BS!���ڸ�E���>���o�}               ,mB1 ��M��=�{O|�Ώ���E�Z               `i�h`��B\{����b����}�             ��Da"FZF�5��|  �P�
vףw�U��*Z���{ɱ/�{~�����>��#Q��             �����@[<6~c� X���j������X���gS*�bzz:`��b V��v���������Wm}ռ{WV���\�;�uq�g����z(               ؿ\.�|>��������T�����x�'b�Ν�ux��b V�����q��� �>������<V7��w�Yǟ;޳#>���G��HT��              �HR����9Z[[�P(dA�J����1<<�E`���CCC122���j���I(�Lצ��{n���+n��x��wk�5�����������^?���               XIR&�`��ڢ��%�������TٱcGDLLL,6�������q����u_�
����	����?�����Ưߘg               ��R��E_ҬY�&�����O��سgO��倥N(��T�+q���~1n}ӭ��-/�w���_r}\��K��{{<��               X*��jg���b0�����ߟ�ki,wB1 ��]ƹ?7�9������bUaռ��;鼸���������D�j�               8�*�J���dїIA�4�L����g�P@�LW��7ė��Kq��ƶ-������7��x�������ձshg               <�R)��L����K
���4B0�_:���"��ܾ��V�}X���? ?x�q��ωkο&����XUX5���O�8x���_������              `R&�_�ԃ0�������5t(�_��;}��7m���zۉo��ν,����}UM�RS����o�/�Ǘ�+n�m[�ͻ]뺸�7��_��3���              h<O���b0i����r9�篡C1 �����9?'�9����k>-��y���E����q헯���9              ���R����P�??�xxx8j�Z��r�\�K��,�,��Jܰ�����_�[�tktm�wG�#nz�Mq��������9쟱\-�Xy,              ���B0###100���Y�%�ׯ�s!���իc���%L(���������mq���ć^�hɷ̻��]o��H��w>o�۷              �cccY�ehh(���g�/�<M�T
x>r�܊	���Y���5t(flb,ƛ��rr2��U.�c||���R4][��Y*ӕ�a�񕇾����x�^��ٻ��{���$!aH�L��xEq�Zg�׹(2*��[�Z��[](�hۧ�>�`U@E�Z��@���TGpDEP�B2<�y+<���$�|N���s����Y�`��w              ���KI���ˣ��t��E�i%��u��1���9����� @�ŬX�"V��b�)Y�f�PL#��������|I�9fL䥚�_�              ��*++cٲe�t��())I?�l׌d4��ݻ�E�b ��5�kb�������c�>��T               ���"JKKcɒ%�|��Q�ŋ��K����2�{�4� ��]��[O�U$            �dG�tDL�35 ��Z�re:�RRR�~��v�\VVДu��!z��4� �0�0�?���d             ��ާĻ_�o/x;2Mn*7�=���a�F�_� h����cɒ%�|��X�lY: ����~hΎ8����
�P tT������o            @ӰK�]⮳�Q�����12E���1q��8�ǁQ��,  SUWWGii���K�)))I��-UϞ=c�]w�P �jת]���_�y��W������q��������            `��s��o��v8(ν��(YYҨ��=N����� 4����t�e�����$��_/^��$��``݊���SN	�P 딜��}��ѳc�:Ϳ�����Ϗ�e            �,��yZ��u�8a`�6�?~��Vq���Ņ] �PV�^%%%��K2j�k��@Luuu �өS�8묳�u��A���[
rb�Q�㧇�4���78I����ńY            �\�:���/|>F=2*n|��=�!�b�n{ lN����	�|���+�|R�T���';�����P k��q�w�O��ţ�<��w^�[6/            �̗��7�xC|���9��I�HzK�gH�|��ѶU� ��*--]~��L2V�^��ӦM�h߾}l��V��v�E�^����(h<B1 �O�\q�q��/�Tvj��KV��������            ��9y��c�m��3�<#^��;~AnA��_Ņ] P����X�d�ڑ�_�8L2.\(�]�vѩS�t���8��������E(��ۿ��q�w�.�w���'�{"ν�����             ����o3Ο������]TWWo�u{w��O�]�������� �Seee,[�,�/_�~�	�,^�8�]RRUUUlY999�LM��1�Ν;���t���B�r㗇�2.;�He�68��e�ӿ�4���6�	            `˙����wX��ԫ�9y������О�ƈI#b�śt̑�G��+�-X＊�����+��i� MSEEE�����/I�%��$�k�K^�&FAA���K2�L������
���hϮ{Ƹ3���������s��9�Ή�K�            �4�5���{C߸��[�}�Z��w?1^��8��3�ُ����ڵj8�q�>gnp�g%�Š;��= d����X�|y:�R�I0�H�K�	�@�H�RQXX��$�$�R��رc���-�P@���?��Ob�1cҥ�Y�fE�yrL\���QU]            @�R��4�=8���d�|���&�M�s�+�.�:���f�51fʘ:_S��6�Ƥ!��gǞ������{�Ǣ��ƕ�`j�/5A���If�ʕ4����t��s����$�Daj�����b Z�=��#Ɲ9.}ҥ.����8���c��9            4m�g���?}9&�����u^r���G���v8(��_:�ֹ���ta�=nl��i���WTU�;@�ƫ���+V|+��t����d,\�0V�^@�*((H�_j�7c0ɀ�h�3?��O�ʣ���ɖD�����+����w�            ��w���n���q�J^�����.y-�LSfO������������:}���d�'q�g��< lk#0˗/�e˖�C0�/N�WRRUU����J����0}I0I�&ӱc�����B1 �خ]v��g���������D�������            @��h���^3?�7�rs�mնֹ]�u���},��zu\5�����L�߯{��g�=��V;l�xy�/qΤsbI�� ���I�/I&y]�^򺺺:��WPP�6���$�Daj�������f�?�G�"1++V�O\����'k            ��k¬	��ܗbҐI�W��j���N��F���rp�8$N�����#7�����k�F=2*n|�� ��������˗ǲe����u2j�0@�Ib0�:u�Ν;��/5Q�$����X�b Z�7�x#�M��{-            ��㽯ދn: n<��8o���;�О�Ƈ��a��6��_�'L_��RՄ`jF�I�/���E�bժU4����h׮����7c0I&����3Z�Օ���WǵӮ����hJ�v�]����L            `㕯)�������}<���?GqAq�s���0kB�����|�� h	�����s��MG`JJJbٲeQYY@�j۶��LM&�NF�6m�"�����oư����_��"9�t��Gǐ>C���'Ǥ�&	�            �f��?L_ot��{b������Ip�?'�g��?@KPQQӧO�_|1�4�T*�����K��7�sss������"~3�71��ѱ�bU4�u�-������v            `��x�������]�x��#++�N�{{��1p����Z���Ҙ8qb̛7/�-+???ڷo��$�5#y]TTT��@s!�B$'[ξ��x�ӗ#����A:3�ǀ             Fr���oN�a}�EQ~��/Z�(���1�t~ �"1��|+S\\��0��	� 4sU�Uq닷�œ/�kVD���ʎ�z��Ü���:�u             '���ˏ�<.;��v]th�!^���8��3㹏�����z���Y}�f �f$����kh��|5'�����'Xzv�g�=;��7,�-�6            ��׹m�sНqd�#������c��3⚩�Ę)c�7�h�>����?��w|+�R\\�6
�lgee��Zv(����UW�}z=�[F�;�[����!2Q~N~���	1���8����a            ���OGb�n��F������v��J@s3e�׹�b%���/��f&���ly-:S��$�.�[��I�
h\K�,��s����H-8��g�>�8̙���Z�            ��$q����*~~��7x3�E+Ōf�)�OY�#v:"f���t�x�����X�`A|��g�YNNN�k�.~���Ԅ`:w��4.�B ��n��bH�!1���ع�Λ�^�겘����[            �8�mO��v8h�s_��R�q������
�|��ѶU���=�G���W�US��ʪ� h��|�̀�m۶k�/I&5��}@f�`��K���;�>�s�'En*w��KN�0��?s|L|ub��*            `����q�wD���;���:nz�����KcM��{fM����L����]�gS٩}��8�_��w�y��@S�駟4�T*
׆`���׆`:t��Z�
���`�٭�n1�������ܶ�&������q�q3�����            l��윸����#/�����]X�0�N����w���jv�b��c�.\�:��<4^��z��x�������/2E~~���KM&yNFQQQdee�<��P�/D�׏�ZQ�"�~� ���QRQM٪��IQ~Q�{`:3�ǀM^���Ǥ�'ş_�s�Y8'            �M׽�{L<1�q����`F�u�Y�y���YY�2.��E���Oş�9���un�����s����).}��XS�& �����X��y]J�+((X�IFM�f[Z���]9�^�Tu	�q}Z�i|Z�iи�ZprBhH�!1���h��z�֛�l^����q���ų?���            l'�~b�6�ت�V띗\�Sߘ�_��K���+���P��b��0�w�g�yF|��� h*V�\�����|+S���~��O �l�;�������튷�,k���Mq�CGeUe             �O��Vq���ŏ�8jY���C&�'�{����d�'q��98.;Ⲹ����7��M�����K^�s�=7}�i�� 	i��(((�V����xm&����� �L(����ɏv?!F���<|���s~�|�            �.��Eq�Anp޴9�⬻ϊ�6�XUqœW�+����=�j�U�s����!��O���+W 4Uߌ�t��)=��$��� ��P �t`�c�~��{� 
�7i��K�F�T��ҮK             #'{���&7��rʕq��k���j���}~�O�=���c@��Z_|�ű��c��> [NNN�k�nm�����[a���� h(B1 ��u��c��cD��g�=7i��5���fM�G�}4�8�	�            �_.�2�=8�̞���Nn<}�͇�eG\�yydge�:w�n{ 4������d$1�$
S��� 2�P@��Nš;#�����8)rS_-L����|��9>&�:1JW�            �Y�͙����/��ŎQQUW<yE<���q�;�7��ƒJ����0~I0I��&
ӡC�hժU 4B1 -Ԯ]v�a}�����G綝7i���z/�y��?k||���             2Oo�f�51fʘ�M�B���7{ńA�^G l)999Ѯ]��1�N�:�G򺨨(������hA��b��chߡ1�ǀMZki��x��c���1��iQ]]            @f���8��3㙏�i�c���8�O����Y\��D*; �1


�ᗚQ\\����lgee@s&��egeǁ=�!}���>��un�^���2�0=&̚��~�X�"            ��6u��|��XP��ѾCr�����s_��Ϻ;�v��j��[GѪ�z}�C���R�(,,L�_� L���t��1����%�h�����{���^�}��y��Wc��q1�Չ�z/            ���T��+��2�LU�U�	f|0#���^1�qq��FK�ey�辬~�|�)�梠�`m�%I&���lgee �&Ќ}�_��ё�/�}��q_�{y\���+            4-7<}C:�i�-��o;>~v�����" 2]vvvPwI襨�(~�	�Ԍ�u~~~ �q�b XkUŪ�2{J��5>���_3�$            P7�|}Puuu��>6��?- 2]AAA:~���������ڵ[)..^��ԩS��� ��P 1�Y1aք�땻�5^            ��0�ә�鲳��u��QVV-I�6m����7��H O(��Jj�����ƭ/��/|?              X��ݻ�;��I*�����h߾�� L���:D�V���"�B�r���
�����c��Ӣ��:              ���={6�PL{���$1�dԼ.**���� ���h���cH�!���W��=���g��}              �?�{���S�Fyyyd������d��$�YYY@� @�Νv��G��ˏ�<����?s|L|ub��*             ��,///���4����t�%	�$��LM&�@��O| �%;+;��7�tc<���1aքx��Ǣ��"              Z�$3{��;w�f_���`m�& S3
#+++ �E�b���{�u��u��o�}h\{����M�C��UU��X������^��}���/������uzz�[6/��������y�             @K��Zw�uW|����lQQ����?�`�P lH�����ؽh�:�ߺSݣ2���O�}��'DS��',S��$����c�.�ư��b�~ãs���^�[a������o�������o�/�              -A~~~�}����K/ŋ/�K�.]�/''�[�d��uqqq�R� �MѢC1 -�;މQ���_>��8t�Ccd��q�'En*��k��e���q��k�������t�f�cu��              hΒ���˖-����t$�]�v [�P@SYUS�LM���m�#���=��Y�R٩8b�#�ci�Ҹ��{c¬	����Fuuu             �ka��١gtl�1rR9��bu|��˘���X�bQ�|�����K��;ﯪXC&	�����0 ��� �`�K�ǍOߘ}��#���3�93ڵ�����8��d���1�I1n��h�G            l9YYYq莇Ɛ>C��^G�6E��:w��91e���s֝��'�7�wܮx�8}�ӿ�~�겈�  �A��,\�0�YX���[��q����u��f�����D�>�?���q�C��i{�#�������I��ڥ�.1���q���������Y� �             ��눝���Ǐ�}�ٷN�w�Sz���1�әq�ԫ⡷
   ��PL�� �-)���9.=�J�}ſ���c��^+;+;����             6��T^���w��m�͢}����O�)���^s�	   s��P ����Oc���q�S��a=��}�Ʃ{��s[            �8�䵉�G<��<t��wd�#㕋_��rA��9>  ��$�UUW��9S����Ǡ}ň~#b�n{o���:U1�Չ�0            P��Tn<x���-S�m��1�qqx�����嫖  �Y�b ��E+�M�ܔ�o�{�3$F�7":��Q���a�{�ظ��k��O���^�/�~���j�W            |ۯ��U��-��оC������;N���  @��`��5���Ȩ����ɥ$sr�#'���dgeǀ��7'�&�0=&̚��@��.            h��������qzu�3Ο��阘�٬   2�P �lUŪx��ӣ[a�t0���ύ�{n�z��T���q˩��#o?���<��cQQU            ��$7j���"++k�󪪫��O����z(}���DUUUl]�u�;qܮ�������:�t�i�>-������G�  ���b ج�-�c��M�>�����GƠ}E�Vm7j�ֹ����NO�E+�o<���<��Q]]            ���穱��{�w�s?�9�?��O_����#}�Ѹz�ձ[��b�a�b���)�/���{<N��xr��  4.� ��Y�͊��ø��Kc��c�~���n�zZwH�g�q�s����            �����w��_�s�Z�ʪ������c�ġq�K��N�C��ԫֹm���C#�3�<#���_  h<B1 lq��J��oM��;�g�sf�7<�w��5�            Z���o�8����f����;/�����S<{�f�}�����?����u�k��*�z_�4<�ug   �C(���W��O^c����z#����81�Ry            |ױ�[k����^P�HL��+���"^���wƸh۪�:��d����kx�  4<� EUuUL�35=�����:=~t��b�n{            ��%7l�ͨGGE��M>ƃ�x0�_�~L>9zl�c�s����SnI�4��gn
  �a	� �薔/�?�����}��cH�!q���F��            Z��n���W������f;�_��~�/�r�_b@�뜓��7�xc�r�3~  @�� ��5���Ȩ�������-����˿F*;            ��$A���/��7���QU]�Y������?��O��w:|�s�X�oN�M���W�U   C(����bU���}�mѶq־g���#k=�            �Q��������}3>��E�Y��,���������]��u޵�^��Ō�2&  �-O(���Y�g1v�ظ�����Ɛ>C            Z�$S��_��b�]Y�2N���8xb����Z�]y���&�M����  �e	� �dTUW�3=��U�           �9).(�uߢ�E[�ث+W�&� nx�zo���C��T\��  l9B1 4II4            ��6ymjݷ�b�?~eUe�4<�|�~g�:�'��I�d���]���  l~B1 d���!�j��w�_�bq|���            ��l٪e���ئc�]:w��$3��Q��4~|Џk�w��.��܂��?r�h  ��b �hWsU���Y�y��W��w            hΖ�XR�Nm;5H(&Q]]M�(*�*��/�u���##������� ��L(              C-)�=ӹm�hHI,撇.�U�b�a�j�wN�s"';'ι�����  `��             �P�W,N��Zo��}������}����/�E��)�+����9����Tn�8,*�*  �tB1              ��y�ǡ=����pP\7��hc���kV���__�A���T^�kP   �N(              ��6�ZC1�Y�QU]���O�:}�_�����Z���<-
r���	  `��              d�$�.��G﮽��y�Gc���FEeE�p���b�����w�}  �4B1              lڜiQ]]�����6j(&�g~�k�����>����9�ka�   6M�Ŭ\�2��YZ��:t�q����ҥu��f��             ���K>�7�����ξ�}���_�U�ј��⟢���N�C��  `Ӵ�P̪����G]���и�PLII��I(            ����{|���m����z���X4�[_�5V�^����T   �W��              4I槇�t����wNF�bw�zw:s����bj�E�/�,��^��ئc  �P             @���������ئh���;i��b�λĻ_��`¬	��bU�u�]���R��e�/ӣ>�
�� �yj���^S�&*�+�<�*�*��U�U�Yu��f��             �QU]_��r�w���Sq����Yw������M�Ϻ;rS�  l����zb�����8���x�^����ʿ          MWY���   �玙w�3�����z���΂w"S����Q��<�@��i  ��iѡ             ����o�_�{v��;�R٩����c�]�"�<��#q�'ǃg?�9�  l<�             �&�����T�:�U��D���Xv�aѻk��쫨�  �n�b              ����e�<���?y>=  ��'                ��b                 2�P                @��                �pB1                 N(                 �	�                 d8�                �'                ��b                 2�P@3�K�]bۢm�)�Z�5               ���h�~|Џ���               �i�                �pB1                 N(                 õ�P̨]F�n���y�6]�	�q�nP��h�.x��(]S                uբC1�S��MN�:��O�и�Ry���f��                �ѢC1                 M�P@36��c㶗n��h��               -E�ŬX�"����<���4�5k���w������Xs��M               �ikѡ���(�.����+Wи�`SYY����!C1               @�ТC1                 M�P                @��                �pB1                 N(                 �	�                 d8�                �'@Z��n���ѻk��ѾG�o�>��I�+]U��ǋ?���/~�b,Z�(               ��!Ђ%!�����}�F�m�FVVV�>WYUO�t���1�Չ��ru                [�P@�a��wn\{ܵѡu�z>���Cv<$=�3&.y�x��               �2�b Z�����0hB���	�e���������m/�<xA��X               ��%Ђ$��'G>�����k��7"�-�6N��D�               �̄b Z�Tv*&��E"15��uT�6�tנ             ���m;ǀb����V�������ͧK�K�E�+���/|?  ��K(����ῌ�w>z���}Ό'�{"��            @�P\P��;'F��u�m���.�w�rW���ߧ� �M'���a����h��]��1��ɱ�|i             '?'?v�ctl�1r�sc٪e��|>Z�Q��\S������.�����h�צΟ�^�=~q�/⒃/��~�����/��5�  l<�� ��$'x6��E���=����ļ�y�hŢHe��C��}���О���;[��z��tj�)�?���_��W             [�6E�Ĉ~#��v���g�}�����+���_��oN�q3�����\7����a��!;��߭UN������rl���k�Z�n�ݢ�����L��  �b ���Zo����9I���.�{^�'���j��� J�3��?/F5:}��6� �N�U�            l~�q�1W���t�e}������s̘�n�uq��k��u�ҮKL9%zw�Y��]v����8��c�W��%�T�)�/�^��V  � 4s��>u�'yf|0#Nwj,Z��N�%'~nz�x�G���n]v[�n��ҥ�is�            �y�تG�m��b��w��g�Ryq���1;G���X�b��'�#=v�c�-S#��<~�������9&  �aB1 ��q�W�7���zl�X����~���8���ū�]��sNr�H(            6�m����/x:��)�n�7��d����b����>���g�}bK�a����!Nz  ���{������˵�Isk�
��B��r�# �P��eDgG8�Ł3�=��3�KE��((

3xA��P�S(��M���ٹ�$��~Wz�씴�ms�|��+����<OX������2B1 cXaAa;�؜��ޞ8��s�*3`m����_�]��S��9?�]�            �?�E�q�'���H̀Cv?$�;庸��Wg_��e^|�}_����ύS�95~���  �P���=�6U�sv۳��������{�w���'�șG���Q\X��L             ��ړ���]���]�~�۱�uu����{�X�9�-y(�\�d�k_�]�QV\��'ǾS���>1�������Ӿ"  [H(`K~�2��?����'�V�P̄�	1kҬxm�k            l�ݪw�+��2��-)*�O�����?��:?�9+�W���>n^x�;�b���8<���/��sN�$vs̬c�7	  `x�b ư�����ؽ1�Z�T����k9�V9M(            ���#.�TIj��m[�,�'}��X׾.:3�1�bJ̝67Θ{F6㰜_wּ�bEӊl4�o=���8��ψ�tӰ��'W<�������+�}%


r�w��  ��ê˪s�/\�0zz{�v�7[ތ����^5}��            0|Il�C.r�������7������y���>N�sr�t�M���z���]���?�k^Y�J�������zK}��_͆g�?�����������  �;��jR59�W�����V�����{             �神G��HB+���'㖅���u�{��8���C�=s��ٴ_TX��9e�u?q�'�*3 �ל���1���fS&N�y�̋V�  �;ס����x���a�_^^�����o�9��vD��q��.�ι��є�{5v4n��             �IsNr��'~8�H̀�F�g�'���l f(��v<������L|����mݖs~�G
�  �0��PL_���c����ع�簷w��툴C1�'��O���~��������T             �f�n�s�o�����-��ӫ��[��5.9��!���?�|��Ż���zR��A��v�/  ��ס             ���������_g#,[�gO�l����_�?�+����H�5�A��&�  ���              �`�*c��=r�������>�����{cT�V��l^6n�|yf�39C15��   �g\�b��<+
V����� v�e�ˢ��7F����             ��Tm�=�����n�/��.��f6h�ʺW"���^uYu   �3�C1��n���T�V�s-�[K2K            `��,�̹�����/ަk���圡��ts��P׫N	�  �p��P             �HW5�*�~{W{���lӵ�;s\Z�Z#�Z:[r�W�	�  �p	�              �`'L̹��ն��n��}�Ξ�ȧtO:�~q��� �p��3             �VXP�s�+ӵ�����}���~   #�P                �'03�����z����s����ǔ�S"ߞ]�l���m               �P�8t،òkG8a��+�n}�V�               ��                �N(                `��                �b                 F8�                �N(`��tS�E�7               �B1 c����.               `t�             �f�̈%W/٦kԖ��ܿ�K��}O�|)-.  `��              �B%E%1{���r���  F�               �B����aÆ����O�4)R�T ��"               ����O>�d<��c�����YYYY6S[[�i�������� ��5�C1Vu�u�>����`�ګb��c�1�=��H���              �KWWW���?��˗�wvvF}}}v�����������۠LIII ���P̹������]v�%���S�g�}f�fi�K���              �G���2�Nz{{���!�r�����I^WTT ��P               ��?˖-�n�okkˮ+V����f�1ɪ��y�q�
��O(             `[ټ2~��c,��t�h��d�G�i����5k�d��J"1���Q[[�)��.++ ��             �l��E�;> �</��b����������)��.]:h^QQ�)�րL򹲲2 =�u(���!{�}~�@`�������?�#Q�/              ����z�V7n̮7�|sЬ��8������l��L�2%JJJ��c\�b�2Z�����?��+y��ed)+.�y�̋�����Q^R}�}�a�Xָ,^]�jt�t             �H�+�2d2�hjjʮ�K��mVPP��՛�1IH��eee��5�C1 l�T��zI�2�8jϣ"U������xj�Sq�swĭ�����             ������M477g�o�1h�J�6�c�USS�)&�'� �K(���:�;�����ˣ��tX_��w��Gg�WN�J|���ė��r�u���y             F��������.�NgW}}��Yqq���1�z�q2`���'�8�[�n1�xB�YSGS4���z�#�8"n����Y;s��Q^RWU��������O�x2              v4��-��dbÆٕK*���I�[�2�qAAA 0�P�W\X/\�BԦjsΏ���xh�Cy��I{�����̆^�a֤Y����1ι������            �h��zU���l���U��X�N�����~Ь��8*++�ј�S�F]]ݦ�Luuu�x%0ƽw�{��ļ���xx��y��>S��_]�EbT�V�]�+N��	���'            `�ڐڐ][�+� �E&������Z�t��fEEEQUU���$񘚚��q�&O�&L��L(`�;}��C�n|�������}jR5q��ݓ��=�JRq�E�Ł���h�l              Ɨ���!#2�T*�)��$$�e�

`4��Θ{F��������[�v��O�>���;����3��o�����              ��J���U__?hV\\����hL�I�1A��S�f� #�S�a�V��M�/���go�tO:/�I1���a�ۜn�^{ �[�\4ll����V9-��6?N���(-*���_z��G���5              `82�L455e�ҥK�S�TL�2%�ykD&�ʔ���H 0���C��|�μ��+�}%J�J6{N�����M��]����Ԧj��]WՐ�K�2�9���3            �X��{��-��q1m⴨��������?��7[ތ��ǂeb��E �E:��+Vd��J"2�d%!�$ 3p\PP ;�P�v����߰qC�i��r�i���C|h��,oZ���i��ڗ7{^S�)���ڸ������C6���/�+�2ں�            ����uL|������yL�0qX_�F��~�]��h�h ���L����͊�����*�I�1I8f (SWW����/B1 cؑ{�s��E�D�/��{\x���
�P�=�8��������Z�ra|�G��?s�JR����N�{z����            l?�U�7�sS��ߙ[���&͊�O�>�x�q����1��� ƒ���hjjʮ�K���R�M�d%!�$(3eʔ����-!0��{��s�?���y�����f���{m����-��c���xC�A�$?X�           `<9|����圭jY�y�7y��������cw�����t�������k���iq�-�EKgK �&���[+�NgW}}���@D&	�|�TUUEAAA ��P�U���_�'�-|sa^��=�]r��p�{������C߈K��4v��}�콳�            0�|崯�I{��s��w�c^�u��c��KⲼ]��9'ǃ�=��t�X0����fc1}}}����LQQQ6�րLr������K`���fM��s���-�[��{$?�ٜ�.�ntf:���=q�S7�5']3h6�vf�R�K�i[            0�U�U�~��������^�{��䎼Fb��m~��_�i�~Z����hPPP�T*6n������FSSSv-]�t�| "3�8NVEEE c�P�5{�����?}��)Vn.����x��|�۞�-g(&1w�\�            ƅ���E�9gI$&���Cr����Ɣ�Sb{I�Y�x���� �Ŵi�r�:`gimmͮ�˗�Gee妈LMMML�:5�L����QXX��$0F�Z�k��5���l.��ʧbY�m�ǋk^�խ�cת��<s�̉_0            `�;}��s�'���;�~'o�����]����S��_<�Xټ2 F�3f�0jd2�hjjʮ��s[TT���$�$$3�^���0r	� �Q�*s�7t4���uu�w��C�\��������:qj            �xp��cr�/|sa��ᵼܣ&U����9�s_�x�����`ق�/���tf����>g�vT�U��e�e�{}�W���`�����~8`���������%�J�- SSS�)"���� �Q�9����y��!����#K�|yi�Kq�>�گ�P            0�M*�{M�+�����}�p�br��͞��}]��/�.~��׃fk����_��x�?b��)q�Y7�G�t�k]t�Eq�o���/�؞�M�ӧO������,�NgW�?륥��2�e���ؾ�b ƨ�	�C1I�7�q�f�O,"�%��Q.�*            ƺ��8<


rΒ(K>����f�y���8�{�Œ�%�x�����[/�W׿_:�K9�I���/�o?�� N:餸�[ƫ���X�vmv�J��ј)S�d�[�2eeel;��1���?���҉y�����Yָ,��֮֜�UeU            c�{�s��/�����r���u\̬�9�<ӗ��z��"1ou���^w�͇��P0j̞=;�͛/��R ����쪯�4+//[8�Ǖ��CF���Z:[r�WN�����qؐ��W=���՞s?_�,            0�͝:7��c���=.>������c��[u�+�2>8�1�|Ҡ�{g�7�>���� �:�hhh�5k�0|ٵjժA��������������������� �B1 cTK:w(fת]���3jf�nջ9f�3�OE�E9��2]            c��ɳs�/\�0o�8y��CΒ��|���n��:�k~-�v��͊���=�^{  F�$Xq�����+V�`����FSSSv-]��m��������d�1����T*0�� �Q͝�9����m���3����/o�%򩢴"�~kWk            �X7kҬ���zϻ&�k��X��E�ě-on�=n}�����_��A�Cv?D(U***�c�X,X� {����`��������Z�l٠yYY٠���quuu64c�P���}}����3�6UM馭�����r����-{,�i�ĩ9�[;�b            ۪ʪ���.���5/����>f��_<�m�Ǫ�U����|o�>S�	�Ѧ��(�=��8�#b�ҥ�|��hjj�����J��lI����>��V����l
��mP��Xr��g\����ꎍ�.%7�������n�s;������I���yg�-o��k`���=���h�l�|�Q3#�P            c����9�7vo�tO~"��:�����ro^�����s�bfO� �Մ	b�ܹ��V�L&��ڲ����hooϮ�8�knn���� �����hhhȮ\R�ԦpL����@L&9Nޗ#͸Ť�ұ�mðϟ<yr ;W����܎H};�6��Es�9jR5�fy�G�:3����=��?���ȷ���˚�            �e�9�;�v�#�8b��S+���������/�ܯM��XS\\�)>1{�� V�hmm;w6�<�IB2I`&9���	`�I���U__?h�<Õ���g8��$��x�ԩ��Daaa��0�C1 cY__<��#q�~g����ǡ3��+n�u/;���x�ȧ�8p�s��[            0��iJ7����N�w��#K�|Y�>����˪`�)**��J�H2�J�2I@f�u����`��d2����K��m�Db���Ed^���l/B1 c��^�]�PL_��Yߊ�w\d�2þތ�q��9O*���z_�Ӽ]���	sΆ��            �C�b
����w�E�ECΟ\�d�Ks�9�~eYe 0X*�ʮ�ӧ�'!���L�inn�F-���J^����_}}}CFd�s;�IV�I2���{�P�v��wƷ��v����{?8��_}jX�O�27�sS���yί��Ut�vG>���	9�:b��            cYg�3�~���U����Ο^�t�K[W[���	U���L�2%fϞ=h��d���$f��d��L���dOH��$┬���A���⨬��Fc�xL��$�rIII���P�/{~%�HN�=5.����<��h<��_�vg���ǎ��}]���q�A����OƤ�Iqٝ�Ś�5C^���:���3枱�����E������f�3            c]KgK��ʲ��b�qؐ�Ǝ�X޴<�;�{�J�J��,;ӗ	 �'	R(r�dz{{���cSLf ��Nֆ���;��IN��ҥK͓���s���S�F]]]6*SVV0�C1�}��|W�/�����]�]��}���Ǉ���(,(�9?{��ㄽN�;_�3�~��XҰ$ֶ������=iv�����#>uu��ςe��7���>�rZ�4礜���<            0�5��s�O.���%�I�e[�g�{����ͿD>���~ssg�S$`'(**�����>}z�s�����E{{�ۢ2�����9����,y�U__?h������l@fภ� ��u(`<xf�3q���}b�s�(L2��9����]�v���%�\�b            �
�$��e����?m��w��%f��r��P��҉9��:���)	S$k��L&���I�1�����{����� ���"2I����*�I�1I8f (SWW����� 0\yϕq��'Ō�����y�7�В��~݋�8�~�'O�|2            `��ؽ1��MQ��4;|�÷)sҜ�6;xi~����ܑ�֮� `t*..���={���[C2�����ښ��$Q�d���%����6����g*YK�.4O�O�j���L�x��!04v4�G~������GyIy^���eU|��OF���1��9g�-{,�2]            �������=��ށ��7��V_����r���Ă7D>�Q�G����O �Mo�%�No
\$+	�$q�dmذ!����6�s�����A��9����>�S�N����M����(,,F��q����y��w\rG�JRy�f�'�Ьk_�v�qW9��Ż            Ƌ�V>�3s،�bߩ��+�^��kVN����=m��3������ȧ�w�?��k^ ƯT*�]ӧO�9ooo��cZZZ6����^ggg [/��l
5-]��m��������Fc��sϘ;wnL�<9�y�b Ƒ߾��8���㗗�2���#�����q֏����)��L���ќ�������#            `�x�����|a�~AAA�p�q�����k~���gc1C���{#��~P���� e�ĉٵ���'���x�[?������`<��퍆���z������:(N>��(//v<��q��+�~����i_�O��(-*ݢ�OB-�={[\��bU˪��=^s�5QTX�s���ǣ��>            `�����cc�ƨ(�4;k�Yq�����1��U�U�U�_��s~���#����g��䜽�� ��UVV�]ӦM�9�d2o�$!��5�Ib�;���g�y&�-[\pAL�2%ر�b ơ�Ζ����!����㓇2�9�������,iX��z_|g�w�5/m��mﺽゃ/r~��w            �'I$����0����4��M��k�㵊��sn�ݫw�+�=�2��Q���9�`{*..�ɓ'g�P��t455mZ���ـLr���]]]�?ɳq�-�ĥ�^UUU��#0��l^�����\>9��u��5iV���g�b���x��X޴|�|OI���o9�����            �77>r㐡��������o��������͙2'�}����}N��~��'�og�;+�~[W[,Z�( `gJ�R�5}����7Fsss���FKKK�8	e$��JB30�$1��n�-�)((v� �:��%g�δ�}]v            ��S+��߼��8c�9��/���+���q߫��3�����k���*��1����gŅ�k�-oƏ����~���/:����o,�L_& `$���Ȯ�v�-�<��d�I<���1��۳+9N���L�XS__.��;,�1�b              F�+��8q����l�s&O������������ȧ$R��=s�^�s�5 �Cqqq���f��ٳ�{{{���%��h��~nmm͞��C=|p۟P             �(�x���+�;��v��S+��?��_��C/r���
 뒀ƤI��k(�t:�������=���6�nll������ _6n��/����/���b              F��.�n����|&��m�h������ۓ��V�UŹ��s֜n��i ��T*�]ӧO�9OB2�����Ғ�sGGG�βh�"��D(             `��]����~|�=����ںڲ��e��"�>���GuYu��=���{� ƪ��̮��s��d���-������=Z[[������^�����V�X�B1              �Ho_o\v�e�\�s�3��[}�$s��=3^\�b�[UYU�ӱ�4�����  ?������6�r���͆d�xL��Ǽu%��I����3���b����/�L(             `���ߏ߽����/����ams�9���oƷ�V�v�n�������T>)笭�-��� �EEEQSS�]CI��ـL���۳a��׍���e�ƍB1;�P             �(��iy|��O�U��*>��ǉ{���~H̨������խ��%�����^��l,f{I����}"��M9�w�xwtf�� F�T*�]ӧO�9OB2---���ܜ]���$��5�BB�1�	�              �r����w|7�e�eQUV�������;��I��c�� `����.9�L&��ڢ��)��ۣ��5�ill��%1���� �޸�|�]��9Us�}������u�ng�������?bcF            �~:3����  ;Jqqq���f�P��t63����@\fÆ������u(fZٴ�=���ϯ+�`�)�٢�v$*.���              ƩT*�]ӧO�9�$����hnn��I�2ɂ�L� `��������ڻ�c]��               Ɔ���P2�L6��c�!���L��������b ư�O�>.?���n}�ָ��              0>Gmmmv͞={м��7Z[[���=�y �De��Lr���0Z��PLWOWtww���,�\�s�%��H���               �WQQѦ��P��t�����Օ=NV�I�2�}��u(�uck$�USS�Ε�G5)��fB1               ;G*��+V�m���2�M����QRR���===و̆�!�丽�=;��a\�b                ߒ LKKKv��^{�uuu1{��(**ʮ���������l4&��$_�~��lL���YH��F(                ���_2�Lv(((�����>}z��~ِLqqq���Fwww���l@�7ވU�Ve�4�-�b                `�mL&	ɔ���̙3�+���7n̮������_|1��0B1              ����:c�����:�  F�	&dפI�6�-Z�(z{{�C(`�џ-y(ƢM+            ƃ��c�n�c$��tEGOG�������cm���������0�����k  @(`{z���            �^��84����2}�Xټ2��.��6x�xb��}   ��b              �*Ņ�1kҬ�:{���S���ts���m�����˛	   ?�b              ț�TM|�=�ͮ߾�۸�w�ĳ��  �m�b              �.N�{z���)q�o���_���'  ��#             �vS\Xמtm��Qq���Ds�9  �-'             �vw�^'ă�=�}�h�l	  "������7`8�b              �!�~P�������L  �wS�N��+W�P             ��p��8�'�HP[^�Q^Ruu1w�ܘ7m^�3u�(-*�5�������k�?\  ��ĉ�K(             `k�h��_�?F����8�]��G�4>����&U���9隸�����/ �xV^^0\B1              l��ޞ�������;/�ˏ�<�t򗢪�*��Ņ���ӿg���  �
�K(             ����tƿ>��q�w�ݟ�;�����}p�Ɯ)s����  �΄b �ٓgg(�G��{��1�jzL(�5��(,(����H>�:��+��ZWŪ�U��iE<���x��             Ƈ��D��t|,�����}�

�3G~&���   ޙP CJj����8e�)q،òA�mєn��V>�_������+^��z             cWcGc�s�9����Ң�A�s<G(  �I(���8ab\t�Eq�Q�����kצj�љd��3�O<W�\|��ŭO��7            0�,Z�(���w������ڙ1o�y�Қ�  �<� �&O�<������T��继�;~p��3n��>�ո����;            ���[�|+�p����p�쨙G	�  �0� ��u|��y�����r��Tm|�_�O���W��CK
            `�Xټ2��.��6�,�  0�P�8VPP����g~#�w����+���������r߿D__             c�_�c�(�>S�	  ����*  ;EQaQ���?����I���K�|)�Ý�~qd�2            �~���h\�+��^�{   �L(`*((���q�!�Hu�A�G\�󋢯�/            ��mu����*�  �΄b ơkN�f�"1K��ӫ��V�˚�Ś�5���m]m���d�)),��&Ɣ�Sb��i1kҬ�������o����h��������s             �[�^�\�K�  xg�:���6d}2��'�s�������nG���{�S�ןz���l�c�ӿ�4~����F��t�$s�>��E�\G�y���暓��'V<�}��            �^s�bJ�J���x�/�  rס��޾�����������-y����܎H;1��ux����p����������w}��楼�?	�|���g�~���>���w����'�����ܯύ���             F�$3����   6o\�b ƛ�O�:f����9K���~�X�l�v�^�]�����柾7���g�>C��{��q͉��տ�:            ��ir���]�.�  ��q���.���/n��{_�7���y���;ʟW�9�׃��o���?{�������1ִ�	            `�����s��{ǽ�	  F�q�y��h.h��e�e�\k���b��1������^~��Q^R>�����#�ӻ㿿���8��s���q\|��9ϙP<!��迏k�6            ��g��Y9��[�  xg�:�x��[t~o�7���ޗ�-SZT�;�sC�����q��H̀޾���/?�{�%g]|�73{�lvs�$�%\BJ�R.���@Т�
U+ڣ�ZK{<mEO߾�}{U(��K�*o+r{=h[���P�\� �����wf�}�ξ`f�&l��3�Ϝ������>τ���r�|w��e�C�V�O�����[����            �.'/?����=�  ���:P/N;��X2wIŽ�сR$��+#��8������>�v�_4gQ��u���            ��rʊS*��ݴ6  �W'P���'�����Y<����z7���~q��9�Pq�G}@(            f�c�;&�/Z^q��  ��b j\:���W�]qoKߖ�l�eQm��������Q�����z�Yєi���H             �ß��O*��Ÿ뙻  xuB1 5�}���sVܻ�Ǘ���@T�$��;�_zϗv؛�<7�����{��            T�3^F����W�{d�#�|��  �:��w��*�'��k�6���y���_��Wјi�a��U(            f�7t�!�q�7&�����-  ����qo:�M��{�xf�3Q�^̽w<sG������r�[�o�o            @�z���U��,�.��?<6_��  L�P@�[չ������~T�۟��b(��            P�������;>�un�R�I���+K�p  ����N�ce�ʊ{w>sgT�;������Eˣ)�#��             fVkSk�~�����N���I����������
 �zW(�J(��-��,��ي{k7��j�<�b��C5�!�+���7?            P�^xp�{Թ3�4J��z^v^�5��ܦ��p��R &y~�ޮ��M��s/ @�
�*������+�o��z7E�������لb            ��.>4����;jŕ�\�x� @���@�T	� ԰��Ί����l1Y(fi��             f���)~��	  ~a۶mS%PÖ�]Rq}S輦-&{�K�
�            �lrُ.������B>  ���������a��,���R�K1[l�m������            �./�^�߹�w�Go  `�	� ԰����냣�1[L�\'��            աw�7.����;�.��  xm�b jXSCS����p��c��ksCs             �e4??Z�����k�3���  �B1 5�)S9�/�c�-�V\oih	            `f�s�5���<�u?��p<��X����{l�c��?ۥ���v�o��  �oB1 5�1�Xq�X,�l7ٟ            j�mO���0�A�H��G�ݗO�#����h  @]�bj=(��v�x`f�ӲOt���짽?�|q�~�            ��h~4��  �ou���bռUS>���3��uz��z���.����	               �O�X����(�a��:                �%�N����|���D___lݺ5�l�2���r1��                ؉$ ��dJ��I�/I&��ݱiӦ����a��               �n�R�hii����hnn.�`��Klٲ%�n�Z
���00S�:ӝ뎞��T���0���g��j�/�              ��/���ҥK#�����XEwwwlܸ1�o�^zժ�C1�c�1:::��80�
��.�n�QR�              `z%񗁁���닮���H"0��d���K1220[�u(�^���q�!'�l�O�>              ��`z{{K�\.W�'!��۷��zzz�P(�*��:��mii               T�������+E_��K�I�ג��b1�^	�                ��F.�+�_�!�$ ��r��P                �Y�)�_�A���m۶���p �O(               ������Kwww�����/�}2�k�1��#               P����J!�$ ��墷���پ}�D�P(T���5�����                Ը��`��K�I�ג��b1`w̙3'jA*��G��a��P|�oE-�wý              �B)����[�/��������l���D-�`�\u�U�              �nI襫��4r�\���M<޶m[̄8 	�{�P               �����Kww����陸OFrT��+W{�P               �466V
�tuuE.�����Rf���$S(f����8�#��C(               �5*�^��K2������Ԣ�;.�����C(               `'��K|��흈���0�}��z���'�|r���                umpp0���&F.������|۶m1<<���N��}�{_477{�P               P���|���Fwww��������H��&�Ĝ}�ٱ|��`��               f������Ꚉ���0�����b1�׮��-�����!��}B1               @����$������9�L&���8����㏏���`f�                3fpp0���"��Eooo) �<NF___i {VCCC���łb��x���Hϛ7/��t0�b               �=��)�$��_���m�bxx8�=/�͖�/�1��R�<O�RAu�               vK>�������K2���c���d>::����d����~I0I�����舦��`v�               *����r�������0�b1��#��N�_���`�(Ly�J���%P�>����5�]{7F=;zߣ��e�Ǖ�\              ���!�$���_���5!���1�ŋ�F9
�aZZZ��%P�>t���S/��_�����E��D=Y6Y|�����~�cq��
�              ukpp�|��r���[
�$��#������hkk���̟?"�dɒ�>T�o@���8'���A|��/ƕw_�Q��m�7>���ƅo�0��             �֕C0�a���J�^z)FFF�����D�%I&��T*`W�u(ftd4RS�&0��oDj;v2��]_~ϗ��~>.���q�Kc����%-<(.:���~;���              ��|����r�%��ݱ}���Z2`��d2���^
�$�$�R��tttDSSS�t��P�@�@l�MU��fVR0ܺu�۪T���v�vğ��OKA�����+?�J<�환��t����o�t�{Թ�Ig             `6���$��������0�b1�����P
�,Y��t��`��Dy�J����� ԣ������>x��mO�W�}E����1��������ѿ���8zߣ             �Z�<��_��K2O֒!3/�͖�/���L2��� Ԡ�}�sq�{/�e�MzL:��SW�Z��6���^7<zC���]�/䣚�i�g���x���իV�O�}����uI              �)�\.�{�R ����IF2
`f544��/I����d>o޼�>���Ԡ��)������}!.:�h�4���ζ���[>U/�^�������w�g���	���?޾�����q��gN9��6��˹Ɜ�P,             �t[�n]�z뭥H0�Z[['�/�L�q[[[@���P̷G�M�SuZ������9��kc6(����������K�{I���wN���]�x�'J#��<�����S?����I<��xz���_inh�UKWő�'|b�|��qȢCv�<c�����������             �n�b1�����ޑN�c޼y����"���P�:�]�ޣ��/W�E�����/�<N���8e�)��g�y�p�	S��t*��wLi������n�il��{7�=/��ͱ}`{)"�=�]�O��!�m�mєi��sƾ���~���e���G���+�!��oI�T�?z}|�?�Ol}"              ��[n�%x�� �Wss�+�/�(?N"1I,�]]�b ��mO�o��q��S�W�u��ѻu�9�s��eǗF5��� ��;<�*             `Ϻ��{Eb`7�R�hkk{E�<OFkkk ;'Pg��ʱ_:6NYqJ|����Y���M�X������[�w��;              �������~��2�L���O�`�ϟ?���舦�� v�P@JB+I0&�-;.��?����h�4F5��+�2�~��ǆ�             ���v�m122P���D&�L2okk�T*��!P����8����wo����Q���x�Ao�j�Dmn{���_��!�G�             `o��{,�^�c0�dɒ���(�`ZZZ�B1 �tv�w_Q�:W���`����_��W�z�o$?k�]���w�����ػ1              fJ��MMM��$����O�g2� ��P ;x|������|it�uƻ^��8����W��j��X1��+��c�����I����>uk�s             P֭[0�d��W�`�!��<�J0�� �S��6�5�]S��q��������C:�X�? ��wz���Xߵ>�m_��œ[�����?��p�             @5z��M&�)_�!�r�<����-B1 쒮���ޓ�+�_���--1/;/���͏���p�����@i             0��r������mmm�dɒX�xq)S�̛7/��t �C(�i�?�_��             @-�����=!�J�B0I���I���l6 eB1   P�F�����   �UŦb        �����^�L&�����������舦�� �
�   �QC��            {V6����$#��$Q��<�J�k%               �*���b��ť L)Ga��---��	�                u�����)�_^�Y�dIi`&�W               ��lv"���$�Da��T* �J(               �	�L&���K�$ ��_�Q����hjj
��J(               �5���D�%I&��T* j�P               PU&��,^�8�����u(�#~$V�]1��W,�������zK�f��?���`              @�jhh(_�L�IB0�(L�ill ^��C1��=$�w���������v���5���b              f�T*����R��y�<�� �k�:               ;���\������2�L���ǂ&0�<�-*��`��               �$�H̜9s���?�QKKK) ��`��d��$�N�����C1�c�1666����| 3+y���C-             `6��쌧�~:jU6����$��a�d��r �yu���uGw�{��'53`fEw��_��(_�             �M>��Y�ihhxE��)�d���_k               ؉��:*n������Q����+�/��ϟ�$�T* �nB1               �mmmq�G��?<c�!�NG{{{)�R�$#�'!���� ��	�               ��8���㩧��\.�Ǯ���P�Ҽ< S�,Y���@��.                �"���?����7�����}�$�`�L9S���� LF(               �`����.� n��X�~}�c2�L)��`��� L2/���� ��!               S�x����G?�7o�6���h̙3g"3o޼H�R �M(               vQgggi ��"                P�b                 ��P                @��                �rB1                 UN(                ��	�                 T9�                �*'                P�b                 ��P                @��                �rB1                 UN(                ��	�                 T9���{o��X�juԢ�������"               �� ԰Ö��<5jі�-               �B(                ���u(&ד�-�-S>���=�����[�L�u[��               �K�:�����Д�	`f�������_�UI(               �Eu�                ��b                 �\]�b67E!U����o����m��fc㷽������=���               �zQס��|����?�3�������\����                f���                 �B1                @MH�RQ,+���̈́b                ���������c6�                jB{{{G�P�a��av�Vf��                ��p*���_^lll�d�lْllhh(,Z�h���}��NX(���	�                 ���Yg���QG�b                 ��P                0�
��/}�K�]��T*U�/444������L&������;���n��'>1UH(                �y�b�|�i�&c��X>>�1>~?�����񥆆��������yST	�                �q�|>5>�Oߕ���u�e��477��3gΟ������s�`�H��q�>G�qˎ�%s�Ģ9�bn��͏�������gc����E��               �i���M�㔁��{���u��������ߙx.B1 �Q��8%~�����<5:Z;^��ޡ޸�����{��5Ϯ	               �i�B!��������zfΜ9g�w�y���� �q�����s.���]�������q.��?����M��'�>             �t:]�T*  f�$ʒ�������[>00���k���o��o��޺�P@x�o��Ms+�=����нaZ��D^��D�1���sڡ�Ń�`\xÅ�/��K             05�������L&  f�$3<<CCC�8K���󩮮����ꪓ����|����k
� Ը9�s��o������7�#���i�ޅo�0.��˧�.�<�k~��X�]_���            ���v͝;7 `6K�ӑ�f���)r�\f�j���w��������j��?���{�ZB1 5�+�Q1������͏M۵N;������N[$�,9�ߝ�w�B��G�             T& ԚL&mmm����b1����P���}��_=��h����P@�;��gN�w�]�N�u�/Z���7�!�g�Z�X�U�*��po��Z             �RKK�H P���t���F.��j544�p���rO]��C1��G6�ݥす��qA�e�b6{n�(�ީ�%q�3��yv��q��n��k�ՙ�bOjoi��~�X�ϫ            �WJB1  ������)
Q����V\}�՗|�c�̞8]�b>��ӱjު)�����z�~�տ2�#!�wA���k-_�<���Ž}�_#_�O�u�z�[�}G�oJ��d�O�;?�N<���ֿ-2�L�ӾO����>+;vG;��J�[��             �J� �e���1<<լ���S7�x��<�s�M���:P�N8��I�n\{�]�����-?�o�0�x�����z�[q�_\
�\�k�Eg��q��N�H(            �eDb �z��d�����tWW�WƧ��s� ԰��Y�}]<��r�C'|�N����YW�]�]�z��!�z殸�w��V�W�]
�l��               PM���W��Ը�t�W(���p@�P�͏��o*�r����s�t?����s��){1�b����~��Xڶt���tC)s��W             �B!  j�l��gxx���k�}�����<o]�bzr=ћ������̬����������v�UKWU\_��i9��б��1���3��o�.�{C���ܿ.�>���g��L�            ��666V��;���  ������|����l6��P(�7��1~��*244��!3}F�Fbddd��'� 3+�����%?h�K�.���s+������r�7t�!��_6���Mk��G����_s�5q�I�����|ЛK��bo��            �v�/k�f� P��HL�(K�R����'�I��b1u�W��N�?><<|����1�FFF���s�u(��-_�������Xߵ~Z�q��'�t��_�ba�ϟ|m������^GkG��xv��            �/B1MMM��d �����t?�J����#����}|�{����J
;~�=9g2~��c4�ו�{���������.8���b�� Ԩ�\q��M�N�5NZ~Ҥ{��Ѹ���_�5�{����:yc�a�%�	�             �����}}}���& Ԍ��8/����|�#W}�������ȵ��{A�<��866V��v2���7��B1 5j��%׷�o��k�,s�3wƶ�m���u?W��,_�|���V             �_�P�����f����\�x �Ile``��=ή:�3����555�c����Ò�J#��ښ�-��k� Ԩ��s+�o������}���t��g��v�ڊ��E��            �W*��T�>��N�c �Y#�^&	Ì����Ź�;x��7?0>}G̀���t�O(�F�6�V\�잖����;ݿ�;c��t�O�=�޳�z{s{             Ժ��P�yqMP_2�L�츝F~�����'f�����6�- �=o�x���t��]v��T*������H(f��+��|B1 5j�PL�����'?\N&_������e������-B1            @��銿��_�eava<v�c;=fӦM�q�Ƙ~����Ԫ����Q����^���<�P@���>�i��e�O����'��?�K�p_����               �ɤ�駊��L]~�뮻���s��i P�z�z*������J*��c�?v���^x(��dљ����              �6���=��df������e��OO�Ʉb j�d��������%���sN�����tj�4W\�,                ��n���)�O�3�
� v�{����:���}�'�t�C1s��T\��               ��������o�y��t�L\?�N8]���Q�z7U\�l������<���>e�)���Ž��O�>�{�z               ^E��	�
���\B1 5��-�O�w��ĥk.ݭ�fҙx���=��=��)�b���+��uv               �L*��T,���k�O׹�b jԦ�M��wc�۾�{�s�n�b�v�ۢ��c��;��3���K������               v�P(lJ�R3u���u"���ç���y;��p�	q����ۏ{�����|j���{�{1��2M��sUŽ����               �W�=�מ3]'��a��������߮�۸�;�{p��g��wL�>|�����Ǐ��(��qˎ+�b~Y�X�'�>               �3�t�?���i��	� ԰o?����bn���Vt��o_��8���cpt�U����W��ՑIg&=�_�ט�7�SV�Rq}c����               ؙb��?���������?����{o����'|b<xу���>?Z��I�s�>G��>��8zߣ'=&	�|����t;��*���ܽ            ��c�ރ���D�  �*D\jAQD�hA�^�`��n���[w�;���ә�gw��O�Ut��p��#��h�(JѕZQ��E֘r!�<�sH�ےh~O~��o~�����.O2��� �'�d2���-@����M�dƒ�[Է��	b�_�����M<���QY]��vEYIY�:.�~fn�w�y�+��c�����iצn}���3�����3o=               �	2�̝G���v׍�b z���[㟞�������c�M=vj�y(��lܰ��nW�vu�s�z�W               ���K/}�����	� ��?>��q�c���������iצn�g&��ŧ.nw�vomlܱ1                -�b R`_v_,\�0����b��Q�z�ׯ�>�۹�΍1Cƴ;��[OE.�               H���x��8�����%���A����־�/�<�Z���}{�;�{�Շ               �D( E6��g�rfܳ�8w���u�u[����̏��ދ�6k̬������5�4���V               ��P@��س#�.�v������:�K׿_�~|����mkn����O�[߫#On~2v7�               H�T�b��l�߿���[ZZ8���oi_>���_�;��_�ta,8yA�3���1Սձ����7~�m�/��?�w��'3���p~�++               �&ա�����Q�������8�v��;vt~�&R.�%����X��j@�3xL���G&��?������5.s$lؾ!�|gH��{��               �M�C1 ��=M{╝��whjij;              ���                 $�P                @¥:�D�����Y�fύk�ѳ!�!�ny;
����                �T�b�˾ץ�s8����Q��               �4Iu(               ��Z�"��G&�	 �VB1               	Ӹ�1�ox?*�* ��P              @���}�_ @+� ��~C�؁�Fi��X:0z���|>r�\�6�F���رgGT7V             �u��xk,>yq�?8  �b �X�!��Ǟ�GO�ӎ;-�������E};u}����Z�5^��j���X�m}��\�-�             t�~_}\��5��G���4 ��� 8HI�������K')�?���_����կ�_L���v�޳U}s}��ݪX��X�ʊؗ�             ��^��R|���O��$�� �^B1 ��!��ķ>��Xr撨(��ԞSVR�,h;w]�+�|����3?���5             ���﬎y��Ž��� @:	� }z��o�������m��I�ˇ�w��N\7뺸a����K�%�             �G6�l�?�_������b��� ��P@ʍ8*X�@�=���C���.�-��zE\yϕ�}��              >���㮍w��c�����F�޺(�]ک����G���q4T5U px�b R�1g�#_}$�����=vv���^��~zY�ݲ6             ��m�� @�� �Ԭ1��_���1�t@$MEYE<q�q�ݗ��7W               ��P@
M1)�mɿEyI�!]_�\[k��κ�Q�X�M������2�L*C���#��A�GYIY��ѿ�<���b�m�b㎍               i&�2K�C�P�"1�Օ����/��elؾ������$�����FM�Ϗ�|\��℡'t���X̊?]�8=j��               ��P@��z٭q�?q]K�%��p������r�!?�5(��o����`�ج1�bəKbѴEQԻ�c�7t\ܾ����+               �J( Ef���O]���{�����]�����{<�并�����ޅߋS|���L�J���]����               i$��L&n�얶�ٻo\��u��zD��ͪ7cᲅ�hڢX�pi���u����7�)7��|.                m�b R���BL=vj��{k㒻/�g+��#������/��_bXٰv�L19.�xq<�ڣ               i��P�e�.�1��tz��c'pt}���i�9-
��o�M��#���Ϲ�ù������,8*�����/���B<��D������s�V(              �TJu(fڠi1i�N�1pD G�	e'���ΎBv����x(f��q����p���|3V��:���������=��iw~���1q��شkS               @��:���ry�s�����/�����{�˧|9.�tI��s�}�               i"��,lw<��Ƿ�V��$�~���œ��{�>h�5z#              @ڤ:��e#��uz}�B
�F���+�6��qd����8uԩ��=��ظcc$���q���c�i���8|b�4:ޭ}7                -R���S���N�/++��jll������$j�TI��ΎL&��ܝ��Iu׺��Ŵ�5fV<�               �"ա�48{��펿_�~<�'"���|6�To�1C�47���B1               ��P@7mԴvǟx�hɵDR���x�w��_�����:�L               �S	� �p���l�����H���|��P�I'               ��P@6�t@�,��܋�I��;�;(F������               H���!'D&�9h|v����t[j�D}s}���47���B1               ��P@6�|x���Լ���"���|l���FM;h���               =�P@6�|D��;��B�s���C1eB1               ��P@6�lX���ս�bg��v�+�*               �B(�+/)ow���.
EG���g              ��H(�+�]��xsKs���M펗�)	               H����P̾�(EmJ�J               �B(�+�S��x.��B�?p���               �DB1 =X&����W�W               @Z�                 $�P                @�	�                 $�P                @�	�                 $�P                @�	� �Љ�N��O�<
���               �N( �.�xQ�	               ��.سgOlܸ���KJJbȐ!1t���ݻw                 
��.����u��}�L&�w\L�<9F�                 �K(�������1�                ��"s�&L��N:)JJJ                ���:�X�U{��ڱc��ԩS�"1�L&�#���!��m�&F>                �$ա����������KJJbʔ)q�YgEEEE G^sss[,��	�                ]��PLWd2����c���P(nXuC�����'�o�               H��N������ǖ-[��K/���� H�����               (l��T8J3�]����E������+�F�Њ ���LCTe
;|�=p                tE�C1?o���]X�����X�pi\9�� ���[��盞               �4Iu(�p�5�Ţ{�3o??��Qڧ4                 >B1��_���Y~��4bR                 t7��n�iצ�y�̸c��hڢ                 �NB1ݤ��.����X��Uq��ۣ_Q�                 �B1�l��e��������1iĤ                 8\B1��M�6ř��w,�#�:��                 8B1�����X|��x������Dߢ�                p(�b>e���c��u����1�bB                 t�P����W���O���q�iW                @W�!���q���ē��l��/�                 �!s�-[�,^��B,�zy�<��                 �$B1G����z̸eF�<��X2cI                 |���d���q���6�T����ѿ�                 �G(�([�~Y����X~��8y��                �Ǆb���x=f�2#�����7��f                 �wB1	�w����G�&^��R��EYIY                 ��I�e�źw���k�ǔ�S                 ա��^�ѧW��k���͍�Ǎ�Y��#%�J��OQ��lC���                ��UR��o���4pR$֮�����ԩS�O�T���\y��q�G!�ڋ_���w               @g��$�֭[���&�8�8p`                 �#S ����駟�ɓ'Ǹq�                H����fc�ƍQ]]ӦM�>}��                 -R]�k�����QH~�������cΜ91x����inn����ڷ,��               @W�:Ӵ�)����д��C=3f̈ɓ'�IKKKA���.��               @W�:SȲ�l�]�6v��s�̉���                 z&��WYY���1o޼:th                 =�PL�{��x�Gbƌ1y��                 z��"���ڵkc�Ν1gΜ(..                �g��a*++���*�Ν                >�����.V�\3gΌ�'                P؄bz�l6k֬�m۶�9����                &��n˖-���Ƽy󢢢"                ��#�����r�ʘ1cFL�<9                ��"��l6֮];v�9s�DIII                 �A(��ZC*555��UUU��͛c���1jԨ                 �O(��r�\444D�~ΥK�Ƽy�b��ّ�d                H.����f��jժضm[,\�0���                H&���{��"��Ǽy�b���                $�PQ__+W��.� F�                @���&��Eee�P                $�P                @�	�                 $�P                @�	�                 $�P��e2�(..                �����>}��ȑ#                 i�b                 N(                 �R���r��f�������o              �4Ju(���.�Uo>4r�Ȁ�����m�
|��               �KR�                (B1                 	'                �p�ŬiY2���Jc��������A��(d�               ��Hu(�����GNϞ�t�s�c{��                H�T�b                 
�P                @�	�                 $�P                @�	�                 $�P                @�	�                 $�P                @�	�                 $�P                @�	�                 $�P                @�	�                 $�P                @�	�                 $�P                @�	�                 $\�C1s+�ƨ����:3 ���db�����h�5               @g�:3g؜�4pR�1��$�䁓��QG!{tǣB1               @��:                P�b                 .ա����H�               �T�b�j��jU�c�9& ������m6�       ���+N�(�p<��Sq���"       ��Iu(        ����cXٰ��1��        �I(                 �b                 N(                 �b                 N(                 �b                 N(                 �b                 N(                 �b                 N(                 �b                 N(                 �b                 N(                 �b                 N(                 �b�0�x㍱{��H�g+��6<�c��㢡u�sƏ                i#�骫�
"z��W<���PL��~q��s               ��#                �pB1                 	'                �pB1                 	'                �p����5�j�566t�\DM�=v�|                tI�C1���Ş�=������S>��={챃�                ]��P                @!�                H�T�b��ث1�оt�l&�{��                ]��P̊}+��4�o�/8��|�� ~���                ��:                P�b                 N(                 �b                 N(                 �b                 N(                 �b                 N(                 �b                 N(            �����o����߹�>�9�/q(�H�D�Vh*�Ũ��a5�Q��J(h6�:,�/�RUQeӑʂJH��ĂQ;�tjK��R4�����v��>�3�}3�$��㜘�������^?'�mE��5    ��                H�P                @�b                 '                �8�                ��	�                 $N(                 qB1                 ��                H�P                @�b                 '                �8�                ��	�                 $N(                 qB1                 ��                H�P                @�b                 '                �8�                ��	�                 $N(                 qB1                 ��a͛�o����tp����bk���]�˙_                ��Pk�8�F>ܢ���8��;��               @b�bȍ�Gb�4@�?�ؚv�gd��z��ڼ                �P��?������
�_bG�t;Q�'�V                M�                 qB1                 ��                H�P                @�b                 '                �8�                ��	�                 $N(                 qB1                 ��                H�P                @�b                 '                �8�                ��	�                 $N(                 qB1                 ��                H�P                @�b                 '                �8�                ��	�                 $N(                 qB1                 ��                H�P                @�b                 '                �8�                ��	�                 $N(                 qB1                 ��                H�P                @�b                 '                �8�                ��	�                 $N(                 qB1                 ��                H�P                @�b                 '                �8�                ��	�                 $N(                 qB1                 ��                H�P                @�b                 '                �8�                ��	�                 $N(                 qB1                 ��                H�P                @�b                 '                �8�                ��	�                 $N(                 qB1                 ��                H�P                @�b                 '                �8�                ��	�                 $N(                 qB1                 ��                H�P                @�b                 '                �8�                ��	�                 $N(                 qB1                 ��                H�P                @�b                 '                �8�                ��	�                 $N(                 qB1                 ��                H�P                @�b                 '                �8�                ��	�                 $N(                 qB1                 ��       �M��X���r��lD�݌+�+       �LB1        �	���oƫ�?��lďN�(���       ؙ�b                 '                �8�                ��	�                 $N(                 qB1                l��阪L������:����b����                6�w��n<��#�����n��l6��j�0��F#߳�ެ��l����r�r,�c����y���G��uR'               ��+
144�O�Z����"1YH&�z���Y@&��~��ɑ�b�����4�^;��\h]��q�}q�v�׻���                ��,(322������e�V����fee%�B����_.�czh:�c��>��Rg)�\l�@�\�\,4b���Y�b                ؒ�����p>�y��`����y8&�W�w��u�Q+��9X9���P�Bs!��y@&�ݜ�K�Ky�I(               �m�X,F�Z�grrr��,���bV2�,//G�ټ�3F��q�r8��tW�l�l�����\>�?�(�                6���(Ky��Bq��/
���t:7�c��L�w�ݛ>�Z�����|���]�����\�Z8����1ߜ�F��Y�b                �4O���|2��ɘ��;F�=�=���7�T������[�w�sS�2�R)j�Z>�k47�c�^��VkCg�G����|V���b�b�Y���6f�R�R���b                �\|X�0�w����)���/ľ]�b����Wۗ����v��r���Ǒ��|��n���1����F�k���|�=���Jw%��1S��'��,4�;�P                �jw�1�4�ϯ����犅b�Q�#��S�'��'�������;��o�r��Z-����n����xL6�fs�gT��8\9�Ϫz�gg�h�l}6��6�F���?�                ��,�rv�l>�9���*��C����C����/����^�x���x>�:�N�����c��L�^���b%�T��vF��[�c�>��c�=�V�l/B1                l;�n+����|��Eb��7�̣1G&��ǿw���{(�JQ���Y�n��h���R��ng�m��B)��+���W~F�s���i�ğW��5ދ��B����K(               ���i�;����z��Z�92y$ߏN�C㇢Z���r��w��gU�^_��d���Jt�ݍ�Q(ǽ�{����׮�ѭ�lcv-3S��K�K��!               ����Z��^�m>���b����<�O�Ǧ��Tej�gW*�|��ٓ���W����1Y4&��v�����J��g�rg9�s�~���k�řƙ�o�G���#       ����P(Ķ�����.��W��Y�ta)�{� ���Q,��+�W�P������_g       ��n��Wf������=���7Ƭ�c���N���gī��u:��pL�^��1�t����hi4�T��s���b��gb�1���Xh.���ϏP        ��D剘�M�vs�̙x���o�9/f�_".^���W�X�/��O?;M�Ўg��      @J.�\�s�s�X{�v�c2�R)j�Z>�[��\�z5�d��D]����ڗ�YU��c�9�d�"2��`��                �-��x�������<"sh���ϮV��LMM���HL�^h<�R�����|V-w��Z��k�d���>��t�x��'���P                �����N�S��=�����xp���5�k��
���c:�N�YZZ�'���vo���h�=�Mvf�\��'O�ۿ��c����_;q��!             �⾱����|�
�Bz�  �AZj.�O�秛v�ʕ�8}�t��9��/�q`�@<0�@�>���]Ã�d����R���J�&k���������`>�]>�ng��.����=|��?��ɦX,��s�=w��l�z���{���	r�N���K/���5B1        ���*M�v�����������4�+   �s�������w  ؞�������,7�j��^[[ɹ8w�3^r�?�穉����N���oś�F(       �u��Vblx,����р��������,�n=        �                ��	�                �c�J�����L�v����               `Ǫ�j���l�F�Qx��go��                ��	�                 $N(                 qB1                 ��                H�P                @�b                 'C�{�}/~���܊n�                �P����                H�P                @�b                 '                �8�                ��	�                 $N(                 qB1                 ��!�Jz�W�O-                �EB1D�����;�P               �-�                H�P                @�b                 '       ���K�(�J���ŀ�
�m���YJ���o      �O"       ��M�O�de2������ԍ���������,�n#        �                ��	�                 $N(                 qB1D�o`�|^      l;'�x2Fˣ��\�����]�]<�gb�iw�       Ő�       �uy룷b[�( y���W�*       ��I(                 qB1                 ��                H�P                @�b                 '                �8�                ��	�                 $N(                 qB1                 ��                H�P                @�b                 '                �8�                ��	�                 $N(        `��N       �s	�        �n��F�.�����������=v������ ~���b'i�Zq�y*       `��       `ݎ���Do"��������x���}8N�:�f3v�v��B(       �b         ���z(���/��B�;w.    ���Ft:�   �Ai��7}�P        ��w��8q�D���+���    ��Rs)�F   �������F(       �u+��1�_�M�&��}��Gc������/G�� �_��L��\���}�(U@����أ"(F��u��$�S<����x4&�$�ģ�E%�1���B�PD@@iK�]�|�|����.�����\�{��<�����      sy�        ��z���)�Sd�u��4V��Ot��-&M�˖-�LSZU1'       `�'        ���	'����J���       d�        �������;�s�=���       d�        �ҽ{�hݺu<��S���Gc�����       �K(         �������'���^z)��m�F���       �_B1         (777�=���޽{<��CQZZ       @�%        ��z���:u���?>��        '�        �WTT�{n<�����/       ���         lrsscذa��.���?�ׯ       ���        ؎���;:u��ƍ����       �8�         lg�����΋��~:^xᅨ��       �a�        �egg�����k׮��C����       h��b         �c�z���.�(����?~        �P        �v�U�Vq�y�ų�>�'O����        �         ";;;�8��޽{<��QZZ��K~~~        _%        ��H�bF��&M�ŋ       �0�         �͚5��;.fΜ3f̈���        �-�         j��Ύ~��E�bʔ)�nݺ        ��         ��ܹs�x�1iҤX�xq        ۆP         լY�6lX̘1#y���       `��        �keeeE�~��cǎ1y��X�n]        [�P         �֩S�8餓bʔ)�`��        ��         6I�&MbȐ!1cƌ䭺�:       ��%        �&��ʊ~��Eǎc��ɱnݺ        �P         ��S�Nq��''c1,       �~�         �E
c�С��o��/�UUU       �-�        j�U�VѪ�Ud�f͚������ڵK�b֯__'kT               �&��ˏ����4���Fu%�<xpL�6-�,Y���U�T                @+((�A����o��vTWW       �e�b         �sYYY��{D۶m��^����       ���b        ��wKލ��>�L3�� ��;��~hLxaB|���M�YUY        B1        l����ia ��ia�8���⦩7�'�06Tn       `��         Pﲲ���.��#�-�(       ���        `��e@̼lf����1���       ԎP         [U��V���⦩7ŏ&�(�+�       �8�         ���������c����ȱ#c��y       �'        �6��̾lv������       HM(        �m�ea�w����߈?��(�,       ૄb         �沲�⒃/���#�s��       �	�         �`�۩_����8��1nָ        ��         �gĆ�       �/�         �����x`�q����럾       �W	�         ��,*Y��|{���M�lݲ        R�        `�+�,���k��?��bM������       HM(        ��.?'?��G�&��nY�2       ��b                 8�                �N(                ���                h��b        ����m#/+/2Myvy,���v�g7�9j�����UK       �wB1        �ڈ�QT]�擜O��/>�m�ov��;��񊬊����       ��P                @'                ��	�                 4pB1        �ZQ��h��>2�ڵkض�5k��׼��U�E|       ���       �����0�02M~~~ �Vnnn���T       B1                 �P                @'         �Ԧi��ܪst-�Zt���(jRY_|TUWŪ�UQQU�W/��+���Uc��       [J(         RHD`uG�~d�۩_��y��ز�&�����\83�/�O��T�2�����       �B1         �O�qH����ql�c�M�6[�^�V����z?=���lݲx������o���       ԆP         ۽���oT\~��ѳ]�zݫmӶqv�����������o�}QU]       ��P         ۵������]�����{��a�{��d��G/�g>x&        �         �K�
[�u�]�p��~(�Wǽ�������>|a�.[       �τb         ���n�;&��=����dT�Q���㸿|�A       ���b         خ��Q��YF��V�������/ǉw���|       @�P         ۍ#v="�h�n�}+�*��eƻKߍOK>�ū���cu���,/'/��7���M�C�ѱe��ٮg�h�#r�s6i�6M�����{�mpL�75       @(        ������o��u$���:^���x��'bʜ)1}��(�(��}����?����sh��ZݯY~�x����[�Y�f       �7�         2��v��g���Ϳ�����-So������x��[�wiEi��ы��5O_=���s�?7�s�w��I�F�۪�U<t�C��w�b���      ��K(        ��7�1ѥ��F�)�(��\�={]�)[So���e��"~=��q�7����,�r�Ҟ���1�~�� ��m�G��mR��Z�V2"��z��M��8^]]3�      2�P         mdߑ1�琍�3{��8��S���ޏ����$��������z0z������'�9!&�9!���ڡ�&�?���=6�z3nԸ�ӡO����QpyA      �لb         �X����ύ�3���q�}gǺ�b[xk�[1��3��z������x�'c���      ��G(        ��u����N�vJ;�o�}q�}gEEUElKk���Iw��F�������m�G����[�̗�Z_y�=�G��(~��       �B1         d��윸蠋��_���(W��#1_*�,��ƞ�_�|�2 �9?8�����U�Af���F��=6z�^       ��         2�q����m�������)cN����hHJ+Jc��#����՘'�!����A��ӡO����k�;r�#�kQט�r~       �O(        ��t�>���]��U�`Ղh�>Z�Q����o��M��){�"��F]�󲳲��g�5O_      @��         ��İ��R��,�?���h�����C.��-�ט��񑗓*7�'?'?����Z�_<�8~��/���:      ��&        @��S�hY�2��o����h�J+J��7�5�\Sc֦i��۩o���kA���ر���>�{��qh�C�ٹ�      �لb         �8�|`�����q����1�g�=���?������(�����&ߧx@�P�v�ꧮNƢ�UUuU      ���b         �8�w�������Gc���b֢Y�o�}k�vd��-;�1=�I9[�ny4�o�5f'�sr\4�()-	2����      �/�        j-?/?���#�����m��䤼�TUVm�z��k��/|�B4&/|�B�P�.mw	2���ώ���o�g�=ѹU������yM��}N����       2�P        �֪E�hY�22MӦMض


�e˚ח����Z�[�n)�O[0-�W翚�x�6݃̓Ť3f����2u(&�x@�P      d8�         2Jana��l����}�I��ۮy�(�-���� 3|c�oD�v=S��Y�NL�dZ�ʞKV/��-��8g�΃�W�^�s     ��$        @Fi��,�l���ј|���ǳ�����PL�(X�v6f���U1n������S�wN�s���/       3	�         �Q6�Y�~U4&%e%igM���/>h���S�95嬪�*�N�?�뵻҆bF�?y�'ɠu�EA���ʎU�����5�,l9Y9��|Ml��      �/�        j�o�"�s�#Ӕ�/`�zj�Sq��j�����
rR����Ҋ�hL֕�K>��¼� 3���)�I*��L���ϟg,�o.~3�t�S�܎-;�1=����~�^g�摗��r���$�6u��I*+֯��Х�K���8r�#����mvNFb��lݲxk�[ɯ��o?�}��V�l��$a�f;Đ�C������m{D���rN��:o��x����?���k����      uG(       �Z[\�82R��F@FZU�*毝_'k�U��?%b+��C]�,�S���$��<i|�����6�Ʊ����y��<�����ypԃ�M*��KV/���^���ث�^5�WTUDޏSk6W"
��c~��>>r�sҞ׶i�8��!�ۥ_�������q��[�J�j������W�G��#Y[�]����,��������s^�[=��Lގ�����}��r{��ҭQRZ      l�         2����ig��Ū�U�X4/h�v�~C�ϓ�c�v����r��lM<���5��3����_����h׼],]�4�z�9���!������b�٩�Nqð�.���F��yS#$b/:�Oq�.�n�:=���_�U�����"n{��F�     hh�b         �(+֭�ʪʔч�M[7�PL��mRO|~+ׯ��ő���r�����5�Z�i<���qL�cj��r���Έ��1ظ�M��c�~,�v���������L��</�L�ٿ�o�o�.
r�l��MZ�O�c����1r���|��     ���         �TTU��5K�cˎ5f���%�-��ŮmwMy|����ϓ�-3:��Yi���5����D|F(f�vl�c<��g�w��u�f~N~�9�Ψ���{g��M"X����|i����ݾ�\�J|���lT�b     ��B(        �����R�b��q�����h,v�q���篜4~G�~T��j������ٹϦ�����[�*]�
[՘��q��e@���kAMM�ģŏ�*SU]s�͍OK>�E%��y~��ܪs�h�#�s����1⎘�lN46�{]�#1����d᪅QZQ훷O>/EM������nʿM��o98�Z      ԞP         ��O_�A;�q��nĭ/��E��!a���A�7z�贳���&#%�߰>��@���y)����bҸ���ׂ��d�'q�s7Ľ3���|Vc�����8$.>��8��	_��ĝ#��>{/�s�?<�_{���<���N�3%��W����3�=#�3�;Ѧi�����f�x���[����      �v�b         �83�Ly��]��$�He֢YA�ֶi�8~�����L�k$�I���ȸ��ˢ��4�_C{��`���2����c?�u֥=���2KI܎��ȸ����C��3OSv�q�hv�a��u��Z�p������|7�%�ĕ��2n|���É���==���k�\?���      �v�b         �8��}6��E]c���Ō�3��KD:��r�������Έ�܂���?~9��콯]c꼩1w��إ�.5f�����:1�y_�����Ǎ�߸�s�z���k6i�g>x&�q�7b���~%���8ަ{��[�I^���9�ω�o98�^\�5��[g�sF,\�0~t؏Ҟw����c�ƽ      ����(         ���~�_9?��W��wz�Ō�;2��E%��ݥ��[��ⴳ1���j����3mL\=����G����s����������ɑ�/}��������w��-����nߌ�v?*��ӒO��ێޤH�?����c�f;D�ԯ�DL�C~�|�      �zB1         d��^(���k?g�9��'k��FC�4�i��7*��7	�};�};�M9+�(�q���z����?;�g���UcvĮGD�������.;+;���K|�A\2�-�c�q�߯��N�)��8�?6:?��s��m������/�����Jyΐ�C�'�      '        @F���)�m�����q�ԛ��:w�sc�f;��=0���q=pt��co?��-��Z������8��,G9��Yq�����.����i�=zY�W�o�>��?�y�{w�;���윌	�3������Om�>*7�E.�g.x&�9�kޅ_      l�P         ������E�c�N�Ԙ]~���_��W�-_M���Ǘ����/~�b�x������v>f��M^�iw��$$�H�x�Q]]۳S�95�,q�Hz�BeUe�������GCw�~gDVVV�Y��r�㩯C�c�����#��yL��Ⱦ#�	�DEUE      4V����z��X�n]�]�6��į_�֬Y���ӟ7��xB1         d�?������q|�V;��q�?�����#��N-;���<�横�
���m��I9�l�g�ĻOl��_7�xS4�kZcֽM�8l��bʜ)�=�sH���c�t��oM��떧�:7C{M;{�����e��~�8W�PL��u`�4�      ��6lؐ�|z�2��ϡ�T��+WFUU�~?W(        ��uό{⪣��n��՘��ƃ�?�͎��o��q�����-]�4Z�q+P�vv߬�bC�M^���$&�9!N����{nϡ�D,g�6;��UVUƃ�����+���7�s�?7�-�a�t�N��xN£o=+ׯ��&E)�G�v�P     P'6'�R^^��-_�<2�         2VYEY\���qǈ;j�
r��3���6��m�0�0Ɯ6&��R�vҵ��lM�xu)ꒌa�3fژ�^����J�9i��{�|/�����?��%o��Ջ�|�g>x�A�b��w�f���>Q�{�V���9�c�^�S���i�      ����^�<?q�L%        @F3}L|w�wS�"z��>��q��gEuuul+YYY�S�{u�+����ދ?�������gENvN��[�ߊ��o�ړ�L���F�V�k̚�5��}G�m/�ۣ=��v6{��zٳ�֭+}:�I;[�zI,*YT/��\83m(&�     2���^JJJ���"�I(        ��VYU�~��1���#7������wf�Y6'�~���V~z�O���H9Kl���w���,h�1�s���v�m������ď�q��9��nC1���%�l֢Y�����6�KFz�mz���X8���M�b��Z�5RJ��    ��csc/�V���J�޿�	�         ��^���h{U����I9���c[����߿�����c[�~eи���u�]Sξ��l���ݕ6s`��W�^�Βwb{ӡe�����}T/{&���ϋ��{GCԱeǴ�����۾��~�Y"Ӿy�XT�(     ���.�RVV�?�t���+WFUUU�p�        Pk'�����4K���_| �N�ܾ1�`t��������:٣��$*!��W<�8�lҜI�p��-���%oǴO�E�.��>�?�:$��vl�c�YIY�]V�����mӶig�y����d�f;�  ۅ�8?����ǧ-��M�.   �_���|yKzIKܗ�!       @���jE�E�i!
`�j��G�/>�UEVE@c׼�y���Ii�c������L�6sV���'O�$6Tn_���$�I�Y}FQV����j[='_�)�+ ���~���S�9������    3m,�R^^������\�2����b          ��Ⱦ#���T1�G�x����o�}q���#?��`ھE�8f�cb��c{��������o}W������ܔU�EyeyگIa�P     ��b/�[��KIIITT���         �z4z�贳-b��/V�ow����ʴ��Ed�TC��TT�3za^�=�����K;�P�!     �����~%���˸˺u�|���Kb�~����@(       �Z��Ϗ&�M"��m���F�&5�/�������;�t= �a��E�b��ű�(ݐ�"Ҳ�e��۪I�h��*���Z��s�X;+++��    ��S^^S�NM��͛K�.h�b        ��VmZE��v�iJJJض�5k��ռ��V�F�
h��=��clm�ٹq�~��o��m4t9�9u���ҕig�����ʖZ�>���^���Y���?�    �媪��'��{�'֬YSo���.1r���s�=�y���������ˋ�����_�bE4m�4��������:�����?N���H<Ɯ������I|߸>�JD�JK�>X�nݺؚ��:g}����?.����c/���>2t�й��#         PQ�Q�FECS<��Q�bZ7i]'�|Z�i�Y���th�!�OW�N:��Xo�vj�i��E%�     ��ʕ+��k��w�}����ҥK\y��P��~`@nnn�y"��X#�IHcnH?� ��V(���J<��Y�E����������M�����������8q�3_�~�o}��>_(         ��9�^���O�>1���xu���t��ʲ���yM���iڦN��d�'ig{w�;�C�퓷�jc�I�N}�m߾�ӯ����c���     �k�ҥq�UWŢE�&?�������j��kGfggO�8q����/
�         �Ѿ=�۱ێ����)[���˨�����Т�E��a��߈���G�fm�I^��KV/�9��$�/|�B�1��GCU<�x�C1%�%ig��x]JDV
r�d����v�O�}�>�׺u��%o����n�,�Y�-_[����yߴ��}�     ��lذ!~��_�k$�.�SN9%�����D���>�h��?�'_         ��T�[7~�ƴ��L�M�Fb���/~z�OcH�!����o�[�a}<��#qó7Č�3�ƫ]�vq\����=��1�������5<���)g#�����,����U����Z7muiP�Au��럾�v�����Gyeyԥ������?'9�9���c��u��A;�v6kѬ     ��u���ܹs�m��;,N>�d���/^wWL�8qްa�n�         c�cp�H̚�5q�s7�˾���m'ߖ�qlʛE��5���==N�{Z��16.�pI�X�"h|��wf��䥜UVU�M/��J��'Z&,\�0.?��d��_5)����μ��땔����j�+���\ԕ��ue���lu�kA����ķ'F]�ψh��Zs>���k��i��V硘�:����J;���     6��駟���sss�?�adgglC��0a�?�b         �X'�}R�٭/��������R�%�h���w��H�eF���rh��c���o�K�ⴳ)s��{$&a���1iΤ8z��S΋oR(f��yig{w�;�JAnA2TRW*�*�ٹ�ư��R�{�e(&�w�{FC���O��$���{�{QVQVg���?*�,�5�2gJ     ��x�������ֿ���I�&�X������b         �H�9�q��ǧ��-_�?w}��٢�E<u�Sѳ]�:Y�kQ�x����?��
��]F�}���Q�8˖J�.sĮGD������j�g���cp2pT]][��}O��-;F]�����������6��:���C.������w}'�u��q�����So���ڷh��x�S�=+֯     �T�@̫��Z�{z��B1         d����
[����5.>[�Y����S�Rg��/5)�'�{"���/�,
��1J+J��7�j��7�?n�c4ɫ�S.�������O]]�����(�,OF��U��=��n�K�^ڢǛ��l�Ϣ�MxsB�.[��9���s��~��=m���e@��7*��?|>�-�;��9�����<�u|���-���C��z�p�;     6�;�k׮���;u�-[�h ��         ���%�O��{��u�߈�#��}N��СE�������?���AÕ����;2�����U�����))-��oOL��<���q���DUu�׮����Z8+v�r�ӣ�o�E�7[�Z�5�Z�y���;⒃/I9�ψ��;������=
s��$<�A�k~�s7�M'ޔr����|��q�=�m�ugH�!��Y:s�͍G�x$     `s,]��^�?���#+++���         #�㐔�篜��|��W��V�&��V̋%��$�שU�d���G�zD��ߙ�������(jR�v~ό{bkK�.ӽM�8l��b�ɵZk҆b����8�ߙ1v��M~�9�9qˉ���G}IDQ�;�h�״�,���z0���1}��M^;���;��e@4&}��q���N�vJ9O��^�����Z�΃b���7��D����"     `s�\��^��ܹs@C"        @�)�-���r��fTUW��~����=v�c��,]�4��tm�?��d$�u)�y\~��c�Ӯ��!�L�C冠a=pt�ي�+�w������#��[m��I9/P\�P��c�Q������;N�#J7��������%"%>��1��ШO���$����ꨫR�[������~��:oj��mݤu�v�mqB���Y�a}\2�x��Ҟs���$�V�=zY�W��z��5-�uM��ҋ�c��	     �\���wכ�y���P         g@�Q�[�rv����|��q�F�͊!��ū��'7<wC2��_#�+��ul��A�}G���c��g�6;���v����U��֖�{<8�����R·�=<����bU骯]+�ZMĊq�T�F=�f���=��x��Ү�g�=�~g�E]M�|e���W�Ua��ٮgԥD�)tٻ��)�횷�g��l�<�����ߤ�;�������?��ѩe����mXo/~;�w���o<�μ7N�����$�q������b���"����_��s�1%�%1z�訮�     h�����         2N�}R_�zI����:�+��S���D��;��hp�K���,��9<��cq��G�<g��B1�9��I�Cҹwƽ��$B �B1M�&D��|[����?IF@��7K9O�azdߑ�������5��Yk��F�fm�C�ɀJע�)�b��8m�i��E]K�zN���x�{/E�)���΍K�4�;�1eΔx�㗓��OW-ZFǖ�1�c�8&oJ�'�I��m�F�I8�����t��ĵ���L~-'ϙ|�A򺶺lu2��S�N1h�A�o�}��M�U�q��g��      ԞP         g�v{�<��TWW��^g�w�F翜��dd���+��{ψ���hUت����D����D ���g��'^��|l+/|�B�_9?m��x@q�C1���	��_N��מ����'o�UZQߺ�[��򏢾����8��Sc�艑������������mS�7������{�m�0ЦJD|���Q1�;S�w��=�]�v��檪�����	oN  �*�Ϡ�����,��i�|	�ٻ8;�o��3{&�e��&��"�5)!�j�P"�S����E���M��.��Ւ�U���Q$��Z��ElY%Dd_g�Y��y��Й��d�̼���{9�}��u͙��q]��  ꆠ         ��AU��������N��*kɋ�~���j���-����7�O��i�ZzZz���x`�A�1����ծW��dxH2 ��$��{����?��~H�CR!o}�V�ֻ뵻bP�A��#�_k��e��;el*Ԧ�=��Sq�'��	S#73���}�'�Ϋ�@���j˪8������L���¦m���Ί��z,  ���A�ƺ����lʬ)1�O   ��b         hrvXi��sku;�:��5����Gc}���Z;0s�W�O�Q��}�ח�42�t����q_4��>T�t�s����������Ćm�c���D�.���5c��1{ŧ�e'  ��IDAT�/O��D��}D���ѿC�]Z+s�?�K�$J�Jbw�f�8��G��'?����ȩ���_�|����+�[�^      �s�         ��tiݥ��Ek��vF��D����o>��k'f�~��8�K�W���y���hۢm���)U��\�f�Y1'ڼ���܏���.�+��}��qœWDqiq��K���0�xn�sqǩw�~]���>ĝ/��<uM�y}{�����: ���ÿ���5^㭏�J�<��3�$�n�s�����8��������J��s���3      �<A1         4)�陑��S�?P���ku[_��*k�e���{O����L�4(���A�|��s�9U���݀�]q���F�}��'�R6�n�њ/-})���Ձ_��<+�xL��m_���򲘱|F<2{�ݱz��J�}���G�m*��v��֢�q�߮�[��5�=��8m�i1���HOK�rΚ�k��w��?���ۻ�t�n{�xx�Õ��h�G;������*}M��im[�vq|��o��O\c�M}��h��f���2����pz<0��xu٫b      j��         ���٭+��V�-�jӡ=�����oņ�������U��.�]�x�ܼ2�Ι���?|=�j[2$��l�D"���]Zu�-;DǼ��1������O��ز}����AK5��`m�칟�Z2e�=����zG��V�z2P&�Ϊwbنe_~�����Zm���$)�s�?�L��DZ�j�+�����:E^v^jLIYI�+X���.Z�(6m�      �>A1         4)�s*�),.���d�eľ]�����Wwy�@���f�FVzV�46� ��k���j㶍u���++/��k�      �OP         MJ2Ƞ2�i鵺����+Zd���^A1k�VYkӢM�޲:       h�         Фl޾������H$Q^^^+��m��3����m�Gaqa��4��[�  hB�����<sr���<?   ��#(        �&���������̍�E[ke;C�W�w����
�)*-
   ��k�O��i    TEP         MJqiql+�99j=�{���]+��{D���+f��cW%�h�Ӻ�ږ�[      ��CP         M���ӪbP��.�k%(�m���_�����\>3jC��֑�V��~[��       ͇�        ��}���.�]45�[��a�h�"ڵ�����l�N��|��أ����<0���U�����DZ�������]n培�J�EQiQ       �|�       �����R��I$4�����>_>��٩��YC�Z����O�˟�<v���������6�n׻��e�       ͋�         ���͍38�B�^{��u�/欘��k��m�}�*�ɐ��6}����Vڿx��       �y        @�����TY��+bܔq;�����~�d�TY�ǢDm�*(fɺ%      @�"(       �j{a����M��u+hX��,�gV>S�{���Z��e�FAqA�f�V��<6��sG<����ۧ}�����p����2l�a��/\�0       h^�        Pm,����FeE l��Y��ſ���
�������>�B-�H��g�����.���99��)���lò��¿Gm�q`*��23��      �nĚ5kvjnfff���UY_�vm�l�2u��S����re��M�V�"==�^�������m۶Tk
�         �$�a�*�I�ҺK<��g�?��-{���вC��ܿ�A=��)3�DYyYԆ1��T�_RV�>�      @�J�������ܴ��(..���\7Y�lPL��n���S�>$�uv����u��g������         �$=:���p�ѭM�J�}���^����+��I3'�k�_�pr`��=��C����4�[��p{��Uk�_UP̛+ߌ�E[      ��EP         MRqiq�0�����;����va��޲:�mX����V٭�k뮩0����s?O�Ԇ���ƐnC*����+      @�#(        �&����>.<��ط˾_8�c^�T�m�(n~��-zA�����       ��        @�U\Zg���x�ۯDNFN�m��?�[�o���r3s���ί���d{L[0-       h~�         Ф�Y1'&�iB�����H������o�s������zv��mWi�م��֢�      @�#(        �&oꜩ������'2�3ke������+��/�:jӡ=�Y̪�v��       ͓�         ��?���X�vqL>cr���o��Z�eu������[�Em�x��       �'(        �f���_��?va|���E��]k4C���+����~S�9       �A1         4+�Ņ�_�������~G�1��/��r���?�����u�bنe�ܢ�b������gck��       ��&(        �f���4�~��T�Tˬ����i��X�um���   Ԧ����q��W�/.+   �         ���E[S   �JAqA�   Ԕ�                �FNP                @#'(            �j�ݮw��mW�m��X�ni    uCP            @=9e�S���W���b��ɱ;����Ψ�?e֔��	   �A1             �䘁���^P������rP�y�i/��`Z,^�8   �ݛ�        �m���"�GS�%}K,��4��i�「*��~�[27   �/�˓-�ZV�?}��b   �	       @���m��FS�<m��h`���ű��V�/I��      �               �n(;;�N�߾}{@c"(               ��N~~~���z���DP         MNFZF��u�h�毜�J�      4g]�v����y�8���A1        T[�N�Kf�hj�o�@�jݺut�޽B���mKj�^~n~̼df4U�~:(�]�n      @s֯_���Ϗ������o��F���EZZZ@c (       �jK�����M����%�J?_�M�3      �����vX<���u�~yyy,_�<z����               �ni�ر1mڴؾ}{����_�"n��ր����v��                vK�ڵ�1c��}��W'�Z�*f͚x`@CI$�w�q               �n���O�w�}7�R~��ǭ���:u
h �dgg��|"(               ��VZZZ\z�q�7�ܹs�d�����n�=��3��QZZz��ѣ7&� (               ��Znnn\{�����6�z�(//���KJJ��.��.�(9�HOO�C�?i����]9r��m�v
�        ���X�1F�ft4U�7,      ��222�[��Vy�1y��?~���q�q�}��\����H$�d�'�O޷�>����{QP         MNQiQL[0-      ��gРAq�7�ʕ+��W_���?>���زe˿ZII�N��~���馛R�۶m����.]���j>���{�g�k,[�,���S!3YYY����ڧ�EcѪU���̬�u�>���g%_˺�VAAAlݺ��g���Q�>�f���{t��'?i+�����p'�                ��t��9N:�Jk��ũ��͛7�BD>"�lɾ�jɾ��Omذ!f̘�3z��EP                �Jfff���ZM�V�Ԕ�                ����)**J�/
�Y�n]м	�         ����=Z������{cŖ     �jWBf�*��l�*df���Q^^���          �B��Nq�~GF��'��)()�[߸5     ���l�L2`��1�(���֒�

���0h�         �����
�v�I}N����M�8    ��S2`�m۶��3�A3�(�����3���7FiiiP;�    �f�/_{�ݳ��[��gN�����1�w����O�5%毜�Sk���'���E%E��hk����-�j˪�x�Ǳz��X�~ٿjm��qT���5�����ݯ���{��q����=��'�����o�uN��+��?8��x���   �ҳRA ;�UV�8�ױ��     ��d�L~~~���Ά�����#(     ���<;�qp������z�i��>.yY��W�u��b&��w�?�ʲ�R�+o�|3^\�b�%�d�����w�~V2�fꜩ�y���|~��-隧�٩�����n���  @�1=��v9�`g�0>Y�H���     P}�2���A37n����hJ�      �P��=RmT�QqɈKR}�P���=S�N�y͋ƦeV���ظ����|[�D"�zN   @c2��� �}��!�ĬU�     �?�4��!3ɾ���FP     @-ػ�ީv��b������<��@�6�D�M���������   h,w_j�� �U��     ��]	�ٶm��d��?�炂����{�Lrn]     P���L9cJ�x�qœW�_�c���7�n��^ã_�~�p��:�N2�   ���@m8���5�k�ز"     ��-'''�ڷo_���ũ��dx̦M��.���mÆ��#��h]A1      ud϶{�c�y�7��Ώk4��$��p�������l��[�i�O   h,:��#���ڐ�H�S��w̹#  j[ˬ�ѧ}�]Z#��+���i������    ��������V����     �X�vQL_0���f�FvFv���j��֦[tn�92�j~xeD�1�qΟΉG�?i��	q���FYyY����I��
   �Ř~c"3-3 jK2(�w�~EeE P�F��._T'k�~��   ���      ����3�?_�Ss��1�:����#���QFE�6ݫ5�MN�xd�#�~'n{ᶨk�6,�=���D�s�=�{��~#���3&�X���h�#   �>%bN�wj Ԧ��m�^��c�     ��$(     ����l�9+��䙓S!,#z�H��|}��#+=k���q�/���4n�n�طp���`�qX��*��zN���m�7�zT&�z]9��   ��4�Ǩh��> j����      �NP     �N*//��?�j�>um\s�5q�sS�0UI�n;��X�vQ<�Γu��θ�Ҡ�S�=5.z��ؼ}s�n/�S�Ͼdݒ�Ǣ�  �ލ0. �����1�����fn      �A1      �`نeq����}o�SΘ]Zw�rlZ"-&�19��bH,߰�����9ƭ'������o��2��76�~��Z�V�g�0tB���3'G�'   �O���>��	��2~�xA1     @�     P��/����x���c�.�V9�C�q�)��I��Tg��q��xd�#��!_�P�8lb������ѶG�����4sR�i�' ��!7'7Zd���&;;;�����-ZT�|I�%vƙ����td�#�Sn�XU�*      ꃠ     �Z�|��8�7G��;�r܉{�G8:�~��:ۗdHKeA1�{����Ƣ��je;����<��X�n�� hBZ涌�9-�����	�aeeeE˖?_2ʜ�F����Ǩ��.e�e�)}O����M      �G�     ���-���{N�Yߙ���U���c��N�b�/��6,�m{|�?�H�9Cω���z���&�M���)�֒A5   P�N�{jd�e@]�oL���=QTZ  �������z4E�,   ���     �#�z'�x⊸��[�3l�aqH�C��_��}(+/�)3�ďF��Bm��	q��צ����;��0�-۷�C�
   �O���L ԇv9��=��'�>  ��R   ���      ԡ;^�#�uطb@�U��谋�,(&i��Iq�QWD"��\���1��Ș�`�.�?q��J��Ν�
� ����(���Ԕ~� V�'��>_�ˋj��=��N-:@}7`��     �^�     �C%e%q���c�S�s�>'EVzV���>,X� ^Z�R�=�B휡��RP����^�UZ�wƽ 4=ߙ��h�>��=������W�d`@}ڧ�>�w��c���     P��      Աg?�8�ѡe�J뭲[�}����{���a��I�Ŝ��q�����wj݉�&Vڿdݒxa�   �i@������%C��~Y�     P��      Ա�Ң�:gj\x؅U��꠯�iP̃s��N�-r3s?��2�e����q�kw�x����8���+��;��(//   �O����0�����[cݶu     PW�      ԃ��}j�A1��V��ߴmS<4��J�]�v�NŌ0:���V�?3e֔   ���:�u��� h�i�qJ�S��5��l      �%(     �<���(+/��DZ����%�ԕ{g�[iP��^ã_�~�p���7q��J��?�uK   �S2�!'=' �i�O�IoO����      ��b      ���m�RA,:�����}���k��><��x���3�����DL8pB\����^+�E~���I�֒�4   P���c��	��ԱE��}d<��      ��b      �ɜs��I�ߣN�b���b���q��*�&��>}mjLu�?`|�dT�K�����y   ԧû][v��6n�8A1     @�     ����c���e[����,Y�d���m���>L�9)�ue$������#�����Wk��C'V����ck��   ���f h����n�x{��     P��      ��2�e�i�'�m�h���������.���_��
�s��S����;��8��ڽ3�   �O}��; ����c�W�     ��&(     ���ڲj��V9��e?�a.�Ō<&.~��شm��O:����k�KK_
   �O���D" ��1=���޸-6m     ��$(     ����"�E���ԹS�'�2��>ן��c���^��ʹi��!_��6i�(//   �/��Zű����$;=;N�{rLz{R      �&A1      �d[ɶ�[d�OP̖�[��yǄ�*��v��b�:�ѥu�
�e�e1y��   ��tR�����4@M�06������4      j��     �zR��cG�Dԗ{f�SiP��^ã_�~�p��J�M:����/�{,۰,   ���%�bl���u��_���x��g ��]2�8�K�ES4�i��g   @�     �����W��U�l�s����c~�INF��ŅQ_����dݒ�ݮ����a5�='���U��m'�}B���;��   ��4�����- ���.( �ԠN�bT�Q�}��    ꎠ     �_��[�}�����ɏ�-(�Ef���3(���<&Ϝ�}M�����<uM���}���!gFVzV��m�G�=   MI��O���+�W���z���y�y�2�忾mض!��l��E[S�%�[����X�~il(�ԝq�@c6l�aѯm�X�aa      �A1      ��cˎ;�o)��i��Iq��#�H|�?y��~#c����8lb��<0�((.  ��UzZz�6$��9,��94�v{�Wd���)v+6����gƌ�3b�3��_SKz���qP 4vc������I      �A1      ��k��;���èOK�-�,�G���
�s��󹠘}:h�2�θ7   v7�:������/�-�k}][w��>1ՒJ�Jc����?o�O<��c����GyyyPs���|
�����c���hS      �*A1      ��G�;��wPLR2䥲��1���ŏ\����X�?��J翷��x���  `w�:�u�6��T8��#�=h$=-=�~`�]s�5�t������)����_Q=������ANzN�������     `W	�     �'���a}���Q���P�~�푗�������;xl���]���gpf��'͜���  И��72�q�7�}N��-���ծW\9��TK�p&�<�0�QP\T��>'F�̖��8}��q�{�GYyY      �
A1      � y!��N����5��mپ%�Ν�;�BmⰉ�����:.:�u�P/-+��3' мL̞m?y45+2Wă�<��sp��qI�%��?yܱ������_���Ѩ��=���О�����ߜ
���[⃍��H$b쀱�;��=�rX����  Hz��Gbɺ%�;��̉�:/z��   @�     PF�iU���bN���DCH^�XYP����c`ǁ����L[0�E� ��&r#�<7���O@������'L���D;+%�:/<����W���t��M��6���ߎ� �{㾸a��h���:�ˡѳU� �݌0NP �/O��T���i1f���q?   ���     �zp���wX����h(�/~>�]}���P���ߍ��Z��3   �Efzf���q�諢k뮵�fQiQ�ܼ2�oXo�8
�
��� ��l������r�`����h��:ڶh��tKԴ�i�K����N�z�5䬸뵻��g���VDs7��� �����պW,ݴ4  v���������ep    ���     �:��`p���w8�!�X^^�
}��1?�P��!߬tΆ��7�   -�Hę���Nӷ}ߝZ#�2gŜ��r^�]17�\�f����x�ǩ�L;#/;/�?�t�'uA]���m��ܪs��I��ǡ��N��_�=n��M��p}4G��ǡ]��Q��Wc���[f�  �]2 �Ư���V�y�6,�?��s    uGP     @�ڠ���(_����L��4y����k"-�V���~ �� @��27Z�����e˖4����hݺ��K�'��V�����w�zG��mk[ɶx��W�E�ų��W���K�Gmڲ}K*|&�����S�:�#��j#���Ny���^nfn�`�bⰉq�㗥?w6�fwu��ӫ���1:��	q��;ck��  h���0ɀ�dPLM�-X�<{K���m���   @�     P��w
�rԕ;�w��ѐ��[��@��~GVk|�D �yj٪e�g�GS�v�� VNNN��W�|�V�-b����䴉�z]|�oEFZ�N�K^�6�i1u���˛�M�6ECxg�;����
=9��qN�3���;�����`�{��vQ|��oŌ�3�9�Iω�{ ��܌�8��q��� �1I��^w�uq���R�7�kk�ָ����'��m   ��	�     �Cɓ)�q����ҝ��;��j�$/h|���  �!�e�Ż��{���ǖ�����=~������5xH�++/�Y�J�?��ԝ�'�_��h��z�s��94^��/ǩ�N����k4u��9>Zg������������w  @C�ަ{\5��8��ĚTTZ�:�x�S����+   �?�b      �H��;N�c�c������pz4�{8�8��h��j��&͜   %+=�Cb����s��/_�e�_9?v�P�ז��j���wㄽO�o���T�s��ң[�n���� h
z���qP���  h(�s�ǥ#/�o�v��lQ�yɰ���>?|⇱x��    ꟠     �:�<�����:�p��O]���1�Z�5u!e�UI������   ���uK��n�߾��(,.��ն�m��g�6���l�eq�^�E"�����E�����7`�� �A��j����ˣMN�͝�`Z|�ߋ��   ���     �e�,�?����|;����Sw�kL�q��b�~��X�ay   4&�>�?�������hJ^\�b���e߸�K�Έ���u�_2P�)�ux�h�#�m^  �!+=+&�?>��ѹU��}i�Kq���K^   ��5���      u�O�>���Ɓ��ḭE[�.���ť/F���UYO��  ��X�aY�0��������hʒa8�4!n�~c\w�u1v���ti�%Ft MI"��1���/��E  ԥ�DZ�<&n��M��5��z���cꜩ   4�b      jAvFv\��R��j�����⭏ߊƦ��<��  ��l]����ٛ��n��%ۣ9yg�;q�������[N�%����Ǧ.lhjN�sb�zޯ���0  �¨���g'�,��_�潻�ݸ�oWş��9u�   h\�      �Ny��ϊ�|�;ѽM�j���s?��3'   5�y���sc�ظmc4g/��r��cD�k�.�����8��I���j��:6^�p  Ԧ/��r�丟Ĉ�#j4���\w�vw���   �8	�     ����ط˾qD�#Rw�;��Q��V�C.�|�q��\   �����XڼCb>����ڂ��T%�d�	��j����ȢGR��  �j����գ������Ѽu���goN�,,.   �q     4+{�W\6�j�M$ѶE��#o���)�v�}���Q0̧�w����?��z��   �b��?= ��>m�ā���� ��ի]������#�i՞��hk����q��o��   �=�     ���]�����6��[��/~>   �/6�Ӑ�?  ��q�	� vJ�6����W�y�W�]��=3�k��&Vn^   ��EP     @),.����9~��OS�  ��I' 4�w;<���+�� ��h��.~0����ߎ�-�=���,��P\���h�    vO�b      jٚ�k����~��Í   P}[tL' 4i���L���� �i��2.�����#m[����i�ť�]�W�   `�&(     ���o=�y0��(,.   ����iNo��S�������V�-  �]fzf�;�ܸ��k�K�.5��ϥ��˟�<�_�|    M�#�      ;a������7S'W&O���|�p   �EY�Yqrߓ�9i��:��yt�u�_ �Si��3xL�x�ѯC��MǼ��bꜩ   4-�b     ��I�l޾���܏���~l-��L���j˪�^���_�5[����Ҳ�شmS�y�u�^�=�/������W���ߏwW�[�kX��]\�k8���ј�+X���wYy�N�����h��V   ���{�r�@s3~�xA1 ����?*n9�ؿ��5��t��������;}�   h��     @3����,߰<F�ft����G4�fNJ����Q'��k��}  @�;}���h; ��_�Y3' ���О��O���8���5������n�_��WQTZ   @�%(         j 737z���[u��Dz�m�6�D�n�7FIYI�ܼ2��_�A��08���K�\�0NP 4S{w�;�}M��ol��+X7?{s���_Faqa    M��         �B�6�cԀQ1�ې8������[�W{~��Ϗ�?x=^�����޴X�iEPQ2 �9;��Q��N��pU  �C���q�QW����i�՞�%���;n��M��pC    ͇�         ���z�;7N��ؿ����V��v1���TK*//�7V����h���������-:đ{ �Yz"=N�wj�zޯ h�:�u�����d�%���]�yť�qό{�ڧ���6}   @�#(         >�>_���8f�1��H��m$��mH�]=��x�'Rw����Fs6�ߘ�L���.�yx������( ����c���������⡹�O^�,   ��        @��o�}���n���j�n7=-=N��	���[��e�_o�v47iqrߓ������sT<�� �?��������Y���a�EeQP��%5��b.����nݛݮ[ei�kj7���e�e��i)nY�"*����"�o�����?�����03g����<f��s��sf�0G��: ��~mv\~����   �(        �6)]P�|)�q�7�0��YK�,愡'�7�f����7jjk��8��qQV\ ��s���( �w6��;.��D2��1}�Dk�f���ڿ   �4�         ���l�3~���Ƹ�㢥(�+����1q��8�3��-�F[��! ������w�?�Y @�ս�{|��Ek3c���r��    ���         ڔ�F����?�u�-ё�s�}n��ӓ��w^�\6��8����>����kk�      �HQ         m�=��>�Xt-�[�WTWĒw�ĊM+b�ƕ��jkl���5��.�]��dF�g��1���(�+l���:(����}$^Y�J�� �u\���{�~/֔�	     ���        ���:�E��n�kV�^@�*))�n���/�5�K�>ҥ-_�p�Jb�o\|��ؒ��eO��k^��ښ]>>?����C�O���)��=���ٗ̎�o9<�\�f��E���~� u$�����O^�I      l�(       �]��=*�h�����$~s�ov�����:�YtO�䩟��?���ݾ�t��＜w̿#�yq���Ӈ~:�qf����۱o���_Ǆ[&DEuE�3���� �~g>+��8-�o	     @��         r�-g�#z���ۤR���ٻ�~5�X�F�<��ښx�Շ3cp��q�Ǯ��F���ǌ�;&��/ߍ�ͿF��K�ř�� �\��nq��G�Co>      i�b         �i��{l\x��z����䙓��%�ƞ���%1i��8q؉1�iѽ��No{�a����'�x2rA���{q� ��}|���      �S       �.��[�����#׬]�6��h���덻��W�Vg�[�W�?��z�9oΉ3��+7�������A�=(f]8+��S�m�D���Ę��DMmM�v�� ��Q�F�����5/ �;��w�W=pU�ʚ�    ���        v�����&�f��W��5z��1�c���t��ן��o?96Wl��������[��?�`��?��ی�=*�}N���]њ������9�ǡ�b  �l�ښ    �(        ���H$�G|a�믮~5N�vZ���l�~��8�'ż/̋A]�{��'^3ΌT*�U�����o     �)�         '=���kd�k�5�q�gf�YZ��[����ώ���T�'���_��9b��
       �E1         䤳G��ӵ�~�ㅕ/DK�������9����w=�q)�      h{�         �s�yq��׻�nۺ���%����qE��u��qF�������       ��P        @��{t���ջv�[cSŦh��o[�ν5.;�:k�:�zϭx.       h;�         �s��Nצ/�������-�I���      �6FQ         9�~��;�x��xi�K����x���cX�au��E1S�N       �E1         �!eC�b�њ�i��-�ٷ۾   -M������w   h�b         �9�:��w�鷞���eO�E�.�3?���   ��b\�q�c�붭�)wO	   �i(�         ��F��=�]{m�kњ������+
�
���*   ��l/�9y�ə�3�   ��(�         ���+�D"Q�ڛ�ތ�dg�7�HFiai��  `O�{T� 欑g��98   ���         �SJ
Jv��ڊU֗���ZqAq(�  `OR   �KQ         9���h�k���њl�ܲӵ��   @c�kd|�د*�  �f�(        ��RUSU�|*���(���;	og'   41   в(�         ��W��;�>����$6Ul�֢��t�'�m��   �F�W{��   ha�         �S�o[�T���:wjUE1��[��Tmlض!   �]ú�c�=&�����^�{Ei��(�+�<�]�um���՘���x���c���Y��в�q�I��i���[1��   4E1         䔊�xw˻QVZVgm`��������ا�>�ί޼:*k*  ��R�WS�N�;��bd��;�]ג�1��8x������̥cnz��Ţ_d
T�G��������O6����}��o��/�   @�Q       �.;���(y�k6�o���]���?�UpT����.OV=��7׽YoQ̐�!���b�n��;ߚ�n   �5G�sdL�45��ݭ���=6�����	��)wO�7־�O�I��\v�eq�1WE�v�|�邘k�6~���\N   4��        v�ؼ��)�)r�[���@3�;�w�O��3_��ޭ���W>�9A��wH�䩟Dk1���z�[�\   �;��.7�zs��%[�<<����8�g�Ŝ7���v�:�����Lh�}<���񍇿��x    {��         rγo?qp������&;{���/
   r�g�6n9��F��^�=��q���WW�Zg�̑g�m�n��ŝ��.����k��/�>   �=OQ         9牥O�;?�lhf����h�u���w��7�   Z���?��M�ݩ�S���{������_v�eq�I7F"���y��ŵ_��@    �GQ        �,��4���"?&h��g���;��ɼ���{�q�C�DKwށ��;�f�X�|Q   к��O��i�'����z������鉛2�?s�g�['k��O?�����W��*R�T    �KQ        ��[�nѻ�w���� �Wǎ�_�~u��k�#�4</}�ڬų2'�}�'�d�$����h�
�
₃/�w��/�>jS�  @�v�aǐ�!>���<��v��_9�+���8F�?:�G�t̼e�2%���`    -��         r����ޢ������G<�\pg�T�x^��ԯ޵�?��   �u�K�ťG\�Oo�|��c�1������b��5QS[��ѣ}��0`B�8��8{�ٙ���t.���8=�x�#?�᧓������_�{ߛ)a   ZE1     9�}O�k&\�UƼ��?^������K�|)��G�=����0��џ��G_�U�C{(.���.;�8��Y�����Ƶ�v��?rc?���ro[t[�p�w���q?�	}&d�����;�z��f�4#F���*7��M��ѯO�u�4(���>�٘�|�s�?>;�w�*��.�E�,�a�)OE�d��rO��)�֦�޿����S�G����X�u���{��3�0�YeV�V����an����ݧܝU�-+��_���\��6����%��Y����ܱ���oO�vV�/�}9���9;�M:)�r�W�ʭo��������\V�.}0���U;�5�^v�KwǍOݸ��uG\':)��?����[w�����㨽��*���w���ɺ�����q��e�{�S��/^��s3O�û�*��=���2  �����k��>]����壿�x�QUS-M�ľ����޵�	��_�   �nG<���ۥ�`����q�7Ƕ�mu��s[��̸뙻�k�Z������X�y���7wZH���bs|��/Ǐ����}   -��    ��.�(�+�*�����(��oA� ���^m-=�mn}����7?Q77��mn���>�]~���L$��&!7�cn"��:3��ޥ�s��$߻d��.�n�N���"7����ސ�{|����^��ɺ���yS쑍��%��s�oHk�� ���M��-�%��/ߩ��_���s�?�9ᮥ��_��eC�]��_�"�m   h�3F��ӵ��I�'Ŭųv9/]��/?�����[��.���a%1O��dL�99�\�f    -��         r�O��4�|̗��^��]s�5����/��b@�q��W׻��bS�:��   ���8x�N׾�ǯ5�$f��ښ��o?#z��	&��1�������ʚ�    Z>E1         䬍��Go�o���:k�:�]��G�����t�-�Hƴ�O�E�]��7�   Z����=�׻�x����c����������3��?G"�����\83s�T*   @�(        ���ÿ�0.9��mp���םx]\��+��]����#�>R�����'n
   Z�a݇e�B���(jS�Y忴꥘���8n�q;���5K�S����   he�     ���c۶mYelܺ��ܦ�M�*w㶍��n�'wk��鏹Ir+��nښ��w[e��7o}����irKR%Y�VTUԙۺmk��e���յ�;\O��d����r�j��έ���3WQ]�un���A�c�߻[�~�n���$�M�Gn,o�=���M���s�5�^��i����#�_�:���#K�f/��K6���  �}���WH��G�}5�+&^[����9���/��'^���Kg]�y�  @�7�렝���_6�}ܳ�-��ʃ_�<_   ZE1     9&]^��+~���dM�����8��ߢo�=�1�Ϛ,7�ڥ���$�5�ho�ֵ7�#[~nS�e{r�l�� ��<���1�;��0����tqgsZ��1������\���    7t.�\���5Kc��Սr����Z�����   ��Q        @����磥zn�s  @�о]�z�_X�B��ǋ�^��&�:k�_����   �>�b             ��E�_�uM��Gumul(���;�Y[�|Q    ���            �=dgE1�76���߶�ޢ�e�   �:)�            �C
���W�T6���,��i   �=GQ         9���,���1}������c���   DTTW   �:)�         '�1<n8醸��k��W����o��mT�V       �6�b         �i������OΌ��ǌ3�'O�$���$       ��P        @�ѻC�b�����b�ܩ1s���\�9       �%S        @�4���[��So��_�?S�ȒG"�JM�6⡇��7�ѣG�5* rպu��駟���۔�      i�b         hӊ�cҨI����W���ϻ=��_4�DM"n��z�q��)�r��o��K���Dt      E1         ��в����~=�>��xtɣ1u�Ԙ�¬���       hN�b         �95�5QUSy�u|2��c�=63Vo^w>sg�>��xa�       �AQ         9g�ֵ��q�����1����D"�ح��Ҳ��_̌W���O����i����   ��r�����>6Z�ޝ��w��N�����K�)�~uv��؍   4E1         �u��eJ]�#}r�#Έ)c��A}����=��'��m�n��bƂ���DMmM   @6�w�Mmt��M��b�    ���         r�[�ߊ�=���ؿ��1i䤘<fr��u���k��.&���oox;�|�θm�m����       ���         ڔ�+g�7�F�0>S�r��s���l���t�WL�".;겘�朘>z���]��rK       @cQ        @�T���?���̸�����a'����pz�%���L$c	�q�I7�ϟ�y���że�       ��(       �]VZR�E��k���h^���QZZwɯ�3�VQ]��pof�����ѾGVy��;�%�]�/��rL{zZL�?-VmZ       �;�        �ˊ�����(rM��h^�����/��D�vú�N�!�;�x���b�ܩ�B����       �]�(         v������^�=�=���Zҵ���%���}�͌��V�����gO�,^~��   ��H?�����E�W.   ��(�        �]�h������ť�.���&�E�.�S85
�
�ճ}ϸ|�噱��bƂ��v��    ����͙   �P�b        �e�+VG�K�YW�.�浥zK�*_Ug���"Z��ښ�+��G��Nq���c��)1���H$��wLf�p�q���b�ܩ�ȒG"�J       l�(       �]v��k#'�@3{`��g����m�3�.�1���8g�9�Ҙ�]68�(�(&���o�+f.��ι5�X�F       ��         h/��r\��5񍇿����c&�y���J��w��㊉W�eG]�.y4f,��Z���Z�5       h��         @#�M�Ɵ��sf\:��8y��1e̔8q؉���kPV2��c�=63�w���E�dJc��       �-�b         ��l���\����ש_|b�'b��)1�lh��:w���]�Co��~5       h;�         ��l����#�̌1}�d
c�}n���58+��      ��EQ         �a�� 3.��8~��1y��8��S�0�0       �>�b         ��T�T�}/ޗ��;ǤQ�b��)1a��       ��(         Z�u���mO���~%�y�7c���       �)�        �f֯S�8��s�3�>��
       � E1         �:u�S85&���>&�D       ��(�        �=$�H�у��)c��#Έ�
�
   ږ�z�}:��3�z��X�|Q��M�-�yf��{��'.��%   4E1         ��F��� �;��աWVYsޜ붭   Z�/���������Z<+N��iYew*���.��rKT�TFcI�v.�\g���$   ���(    �����K�5����a�غukV��'�07�thֹ]���ݧd��s������+�un���ur��w�:w��}��vNv�:wX�:�%���sGu���G�5�Y��<6���G��TlMe�;���_�����I�d�{dّ�������_>��A��cKՖ����f�[����PV\�un�*Y'���Y禿�>�;�Ӡ�s�j���o?�I���%���M�<4�^ַ]�:�=
zd�;�dP��.�.Y����`n�DǬs�+�/�zW�0W\[�u�莣c��^;NVFl��r�rh�k�/�����1�ݹ @v�'�M5)���L�*k妕qϢ{�O�4�[�\   @}�~��3%.t���㗋~   @�(    ��]2�(L6�cذaCVǗ�w�ܐ�5zn߼�M��/�_����n��wȾ��{`�3��s�w�;��>���?�;�|/�2��Sz��P��Z"��3��Qgn��-�����_g.��m�'~�Ir��g"�ʃM�[�ޥ)rK߻4EnS�
4I����1|��F��~Lf4v��N�3��s��rDf젦i���m��e�/ۓ^���� ���.�]|t�Gc��q��EA^�ng����c�?S�N�{_�7�j�      ��KQ    �@�;���zC:�D��>QZXE�EQ�_�lK�.�T*m����cŊ ��o߾ѣG�hKF���?�b�rU�VEEMEl������77���xf�31����� `�ڿ���r��s����Ҳ��^Z�R�1���6Z�ڴ*        MQ    ��z��S���>4z��3   v� Y�����#�F��V^]ϯ~>�������Ǧ�M 4�>��Y#ϊ�0F��Uֆ��g3̈?���       �R    �h���b��S�̡gF���  -A"�Z����8����q���������/�y1 ����=e�Sbʘ)q°"?���W���9oΉ���]��[*�       쌢    h���q���a�D�v  �)��k�<>>:���7ϿYa d�ʣ��;ϻ3ڷk�U�k߈iOOˌe�       �
E1    ���OҼj�Uѽ�{   �	�D"�{x��3>�}�޸�cS妀ݑ|����5�D*j߻ �'���%��̧R-�����������q���b�ܩ�ȒG2       4��    �C����?r}���   h�D2�rF�����+c��9uI�%�)�)r�[�oŌ�.@�7!�(���|u�:�U��=�8ڷky��7��91��i��g�7       �.E1    ���>*n�xS�.�   ͭ��,�?5n{���3?�T* Ж�%�b⠉1e�8��ӣ�]iVy+7��{��ϻ=-_       ��    @;�����ߎ����:>}�fmm�����[  h
��7�����+�Hd�����d�3�'�_2���ip|��/EU��9 mϘ�c2�0�>'��v�*���&{���:wj��½�m      ��)�   �&4i褸z�Ց����WSS��r��1�.�| ��.�{����g{aL^^^fl/��g�plL�����ß���[ r�����Qg�'�|"u�u�K�^�;����O�U�V       4E1    �DNtJ\3�]:93]S]]�y  �;҅�ۋ'�ҥ1����Tsh�C�o��0*k*>L��K^��56l�yG�.u����.�"��>��Y#ϊI�&ń"[�7���.�ϟ�_�       �'(�   �&pD�#⿎��z2f����*sB'  ��RvH�W[[���[��.�)((�Я����L�N��#��9
���(���\SRR@�*,,�����/�廕��̏�0�?��8b�#"�Hf��jS���G�g�~�}ᷱ�j[       ���(    ـ��;G'
�;�MMMM�M'_  {B��2=҅1��w���G��|!n�s @k׹�sL�45뜿o�{���]1u��X�fi       @sQ    ��0�0�3�;�W�^����a�1�  �=-]�~>�.���˫�6���xz���� �V�W��}��f�/?5��{       �OQ    4�+�2�uV�Z���tI  @sJXVTTD~~~�0惒�d\����_��*7 �%�� Ss�;c��5       -��    h$�w�?&�T�Z� &]  �R������F�v�"�H�֭�[|��/�5�&  ׭ݺ6~�ܯ�G�Q,Z�(       ��R    � }R�5���d^��������	  ��&]S^^�)�I&�;��5��������W? �kjjk����s�ƽ/�U5U       -��    h'<!�����	��/  Z�T*�)��`YL2��K�^�z�S ���w^�iOO�i�ŪM�       ZE1    �>5��-��   ����b��#�F�s�� h�6�o�Y�g����c�k�       Z+E1    ��#�û�a���2jjj  ���^STT�D"3�~{Ѩ���? ��l���������ɼ       ���    �Ҥa�v�^]]�   ��?��lw��GD�α�|] @k��bs���]       �BQ    d���4�s���kkk���2   Z��󚪪�(((�\/H�)�O��/L         ���    ����������+�  rA�(&///��d��	OP        ���    @��������Q[[   � ]�YT��Ř�w�?��c[��         �y(�   �,�����T*UUU  �+�E��B����(H�!��'�z"         h�b    `7�ܫg�ثG���ɓ�  �\�.�LŤ�� E1     M�#�|$�_:?����z�o��q��+���20   �=OQ    �};�����  �\�.�L?�I������    �R��N1��&�ާ�>   �~�b    `7�<(�6}�d��I  �\��(��� �IQ~QL;%r�=�����       m��    �M}J�dަO�  �U����ѣ�G @kҾ�}�z֭���x�	E1       m��    �M{����	�@˔H$�C��QTT�ڵ�d2� 4���P555QYY[�n�M�6eF*�
��I��         �GQ    즒�ɒ@˓��={������� �<����� S�.�J����ձjժx�w��5�t����s����(�+�ʚ�         `�S    ��(��	��u��=z�� ���Ϗ>}�d���~;֬Y@ː~�J����DQ        @3Q    �)}�dMMM -C2�����G�.]�֭�� ����lٲ��]@�K��$޻     ��g�~&~�藑��-�   @�Q    ���VI�������FIII �;�u��ڵ�%K�d
*����    �qL�;53    JQ    ���� Z��*��Q�۷����z �KQ �M��y隥њ���;��       ��    �n���	�����ѡC�  wu��)z��+V���T*�A�/ hm�n]���M��Nq���c��)�O�}       �S    ��6U@�*))����  ���b֭[���4E1l�����&�Lм�D��K^"���J&�q��3�0g�<3J
J       >HQ    �&E1�����9��ܗ��������z �CQ�u��%:u�\Ӿ}� �Wqqqt�\w����\5���8g�9�Ƀ?�;�       �0�b    `79I�Wii�9ژ�;fN޶m[д��3
3 {��;�9����8��!����|cl��{1      @[�(    �V��W ���K:u�(���L �=�D2�|tL;%�yf��48#]�6��91}����pfl��       �-�b     h��E �=��Ŋ  ��в�q���c/�]�VƲ����w�ԹSc隥      @ۥ(    �V�]�vQXX �=%%%���555@����(�/�\�i٦ ��_��5��2��|Mm��ݯcQ�8��Sc��q��c"�H48cc�Ƙ�xVL�?=Y�H�R��%��T\u�U��v]�v�\֯_�]������     @Q     �O�(�����(�l� 4��6<9ic ���o�Sk���(�H���3�0�t~�U�W�3jS�1��9�r��g��͑��vX �u:tإ�p�s�      �b     hu


��+?��� �eR6$�;�`�1�ˀ��X�~Yܽ��:wj,]�4       `g�%     �N"� ڮd2  �\:u��8-&���>f��;���1k�>z<��H�R       ���         ��D2��)�9���c�½�Q���9o�ɔ��\836Wl       hE1         P�~��Ź�vq�2p�2��_w/�;�ΝK�,       �]�b         ��ס�C�v�i1y��8f�1�H$���|c�Z<+�ϟ�,y$R�T   �v�=>F��h��q���   �4�         Ц%�?`|��ϋ�v�ΨM�Ɯ7�d�af.��+6   ���N���8rь3�   @R        @���#��>�ۻu�w������,[�,       ��(�        �M�O6�O�6�o�Y�ge�aY�H�R��y<��c������M�4)�;��e�^{m���K>n�>}�m���=�P�����+c��ё�������n�qݻw�[o�5      ���?��ή�>����̝=�d&+� �����BYd���b�
J}���
�>�}����>�"}Ԣ��He�� �
��HX�0�d��r�9c	������~���5�s�����ef����        `zs�qϳ��q���N�v�c/������~���1ٵ���c����dr�����ٍ�����     `�	�         �nԵ����4��qC       �X�        �ݨ)�������o����uK       �X�        ��p�㊷^�=��~W�{u���i<       ����������Ҳӟ����۶m۱.7�}�         � ����I��������o�W�sU�y~M   �@}���c$�~�5�
�vY~�΍U�
   `Ϻ���zihh����?�^vD^����tww��c�        `J{���hlo�����gz�����q����?������       ��+c/����V�%	��r���b       �I&�	 �����^7��)�ZzV����8uɩQ�7����X:�p��'��$������� �{G�jq       ��Pc/MMM�����P         S^gwg�zhU:�V̍s��<⃱lβ�QTPgxF:^l~1V�vU|��_��^x(       ��W_�����Z��dYr?v&         ��B��;����V�����z^Ԕ�x�9s�c�~,��[�Z���v��Q�V       ͫc/����V𥡡!r�\0<�b        ��d�y1ټ�})~�w�΁�9E�첼��vC�1V��K2.��8s�q�����%�FA���Kb3ɸ�W��a����[���;       FK{{�N!�$����Kss�n�3>�        0`��GU�*&��0����軽Zwf|�T:�;b�C�ұO�>��C�<�q@�1PEEq��s��|��q������Z<��      0P]]]��2�R__�,߱mr?&6�       v��� ��K"/W���t���".8�x�!�iE�<G���Kұ���q��W�w�|7Z:[      ��v{�1�e��KB0�񚺄b         `���˅߿0.���8s�q����%�E~^���Hb3_}�W�K+�?z�G��ߊ[�%zz{      ��{ijj���2xB1        X~~~d3٘l

Fc-///�ى�����#V=�*�*��y��~�����x���8g�9�x����ߎ���?⩺��=����e˖�v���>uuu1-Y�$jkk�]��|�=������c��]�z��hoo���������~�566��?     L<�|���Oǫ�'�&����       v��d`w�Ϙs��d����ؚ6mZ̝�����ގ�'cBI"/W���t���".8�x�!�iE�<G���Kұ���q��W�w�|'Z;[��%a�O|��]�W��w�S�����8���]���!�.�:���?��ݮ���?<eC1]tQ������m����]     0~$���k���O?7nL�.���;E_��5��<C�㸭��$�{<�c�r�ܘ�k�یB1         0B��˅߿0.���8s�i4���O���Il���j|��/�MkoJ�1w<yǄ9P      F[������;����a�?y�o�ʕqꩧƼy󢰰0���<_CCC������*�3���ٙ��&��e�nݺ�ߺ��b�s뮾�?������O�����        �����Z��y���Cϋ��X\�x�s�dK���cɕKb��u      ����E|�k_�@L"��|�#����aT��\.wP��W�X�n��o�8��^��P         ��皞�+ve:V�[uA��!�E$     ��q����5�\3b�_z�q�I'E&�	a�r�܏���k{{�_�{�=�B�         #��[~�����2�8��4s��':�      ��k��뮻n���+���e+..������d29�         &����XX�0&�ј�5��}��/޾��Q�-	      ���׿�U�V������Eb3�L�7�|�}�~N(        �Igz��x�o�
      `r������\.7"�WTTĻ����������M7���                &��n�)���Fl�O~��f�XA.���b                ��~�ӟ���˖-'��               `�y��c�ƍ#6�������DV(               �	g���#:��0��                0���׏���f�
O�b                �p���Ft���Ҁ�D(        �I���>��☬66n      ��r�\�T"        ��������       LB1                 �P                �8'            0J>y�'����>"s�dK�]~��W�%'\#�Go��n�,   ��!            0JT-��V��>���oT��v��    F�P       ;�d2         �/B1     쵼��Q�_~~~ 0u���?w         ��@(    ����f'�� _��         �"�     ��h�@_P��m��l���         ��h    `�������JKK��k4d2�Q�9         ��     �Z6�MO�ooo�}0u���G~~~������M�yyy     0\x��X�Ъ��~���   ��     �Eee娄b�� @EEE444��~��\.     �ȸ�ޫ�   0XB1     ��3g��͛G���d? 0k֬����GMMM ���i�QY<��eee�����~�E=E       �     0L��l����֭[Gl���QRR ��̟�D���4b�H�dS�-�L& �S�-L��l���|O�P_�_z�{       �    `͞=;��룧�g��NNX�;wn ���O477G.�����g͚  L\3�gĖOo��jɕKb��u      ��!    ��),,�}��7�|��a�{��Q\\ �CIII̛7/6n�8��&q����/���         `��    `XUVV��ٳcӦM�6gmmm: ��fΜmmmQWW7ls&���� �k��Ɩ�-1�lh����ܱ9j|h���{�            ��g�}"???�����+	 ̟?? `w-Zyyy�u�ֽ�k��1cƌ `����WbR���}��/��2�~��   Lv���(*(�eyWoW�v�   �G.�K�H���M�x�<����0R_���w��<&�     F��ٳ#���ƍ���g��O�LH�3I( �$	����!�qZP.����      I�|�?ǅG_����1V~ce   0~l۶-�l�2��ihhH�5����eee#�����t�G�LfP��     0bjjj���2=i���^�����c޼yQXX 0P�f�J�$������'y�uƌ1w��Q{#         `(�b     Q�p�3gN���ESSSZ���r�&9I���$��$q���� ��H"c�/N���\a%���;�����K�:�De����         ��    ��HN�Ob1�HtuuEoooz�~6� NItl����H"1����ϝ���t$�2  ��/���x��a��c.�UvY�?O�Oܾ��!�[SVs��       $�b     �0 ��$
��  ���������a�����7s��wŕ?�r��.�Y,      ��    �M˟۷o��v������#���'  0��-;::����[�����~JJJ��wٓڢ�h��         �>�    ��Es���u�ە��G^^ވ>����hii	  Iq QDF^[[[���#���s�Fii��[Z�4ַ� �������û]___S�UW]�\sM��z{{^��[o���k��7o�Sե�^���f�~     �H�         &�$v8������!0PI( ���h*Gr     ��'                0�	�                 �sB1                 �P                �8'                0�	�                 �sB1                 �P                �8'                0�	�        0`5y5��M6�3ۣ�����Ly�Λ����\ol�m	       ��b        �w�+�rU1�l,���c������첼;����|       �T'            0��= .9ᒘ���Hܴ��    F�P         0!UVVƒ%K}���ژ�-Z�\n��+**
��9s�鿧����2�̐�.ӧO ��:pցq�[����[��%  ���������3`<�         &�+V��]}�#	��+W�����?��     `|������l�0��        0`�Օ1+;+&�m۶0����b֬]��t�vF<       ��?�������[���B(       �+,*����l
[Q\�����       �עE��Rl޼yD�_�zu�r��d2�@N(               �	��o~s\w�u#6����c�����/�b                �������-�����#2������W�0�z{{?%               ��TVV����\�;�O<1`}��ϾK(            `���ȍ��+  ��;��Scݺui�e$|�k_�ŋǢE���=���%��                0�}����������Gd�O}�Sq饗Ʋe�FK.��qIIɻO>�����B1         ��mY����,���       FG�������={v|�{ߋ�۷���\.���1�>��x����l6`��=����ҧ?����b         `/����?"���z�����u=��       v��d��|g{����~7��a��x�q��7ǻ���8�裣��2�o2`/u��{��}ϧo�y晻�a,        �����W�{u��n����O���{z       �3{�����������7��M<��3�aÆhmm��hii����]����;����t$���c�ܹC���#���9��5��[^^ްϛ��ҿ�+���D~~���+��)�<����e��|�3�'��}�[N?��=��-        �����~��       �����8���w�����јm۶��IF���uMMM;�\:::b����u�g�#               ����f���:�5��LCCC�r����               �A��L]]]�H`���9�����M(                F�P#3;3��d^+2��������'                ��P3��Ff����C(                &������ECCÀ3ɲ�~/�                �_C������y��LSSS�����                ��P3��Ff���7&+�                `���LCCC�r�τb                �Ia8"3uuui8f ��dYr��                 LyC�̴����I�1��477��I>&c��b         �t2�LTW�d���=�=      ��+))IGmm����ޞ9����         &�ڲ����-1Y-�rI�ۺ.       �:�b                 �9�            �Qr��wF&��e�C/<    �E(            `�|��o�   `��b        ��la�d��f[����~���       @(    ��~s}ln߼��jjj"//oDKkkk���K�6_rB΢E�  �'�|2z{������a�]w��ڢ��x��M�P9�2*�+b�)--`lEEŮ�_�z�       �   �!�޹=��n��v%%%#�ٶm[����|N� ��K~7�PLggg���HK"1]]]{ܮ��0         B1         L:�:�ť7_:b���������<�������m?�;�s���5   ���]�,:f��\����]_   `d�         0�u�ŕ?�r��?�u'���m�m��{�:l���i���   ��U�*.<��]���ȍ��+c"8r��q��svY���qW    #D(       ��������1�tn�`lݾ����C_�eyOoO    �����l�.�?���ƭ��   ��&       ��m���RG c�i{Slض!   ��[4}Q�����<   ��O(                `��                �b                 �9�                �qN(         )/�       0��b         `��
�       F�P         RUIU��K��ö�������w][W[       0��         � ž���w]eq���z��:�      ��E(         aٜe�����nִYö�Y���՛����       `j�aB+������ƥ�E���촾��+�z{�Ϸ�tD.�   ��R1�"�+���]UUUd^���p+//����a����K�  0T,����a����=��l��Y�fEII��{���  "ޱ��]�bފa��a��wyKgK� `�)��Gq~a�yq^6�y�;�ߞ�Ξ����ѝ�	    ��r��Br���ly�.��ŕQ�-�i%Q�-�����c���oYyAq��y_=�������m���������m�Ե-�ƦΆ��ј��   П���(�+��vI�%//oDKQQ��  �555�6W[[[l�>��Y���Fii�OS[ �TW^T�;�}�]�|��t���ֽ�����w���M ��K�c�]\3
+�����Ƿ��ǸO����q��?�}o�v�GK�h�j��Ǹ����dy�������;�?    S�3G5I}^IM,(�s��cVQU�J>W��g�F�队�{���{� ^���ѐ������x�����M�:        `����bNŜݮ/�/���޸Ɜ�j?ӊ��9���w݃�?  �䂧���ba٬�ST�K��ܫ�e�q�{s���z96Ss���q۶�Η/��٘뾩�1^쨏g�6�ǻ    ��P#"y�za��8�|n,(���>/��y٘h��e�x��y��K��϶o�'[_�g�m�g�^����+        ���������?���.>����o��ݝC��EtQ��Ϛ��  �SZP�׼|l{r�{ɌX\>'*
Jc�I�.�̎��f�.��<�Qڶ��q�m[�m/FsW[     �P{-�W�+�o�XK+���O�*SA�Y:mA:v����/�?��l�m���qCl�Te       ��,����Y��Lf��.��$>{�g��?�sT�?�:0.?��ݮ�� ����������ba8m~z�����
��L�IƉ3��a�����yC�m�k��M/���    �P�V�-}9��Da*���$���3yi�=g�92]V����l�G�6�ھ�Om����         Ʒ9s�+o�J�<h����o��h�l�����G.7�p��Y���-Q�-�w}GwGܷ�  ��e������x��I0��5�dz:N�up��־�+M�1-���gc]�󱽷+    ��M݃=����/��T-���+�Mc(\MQE���xS�A�[��������񩸯��4$        �y�>�;�sQUR���~��O�M��)
�wZ��d�ӧ|:�^xt|��O���V���ʋ��c�~,.9ᒨ(���v���-�;o 0��:=���鯏C�Ga���Q^P�O]:I$�����ǹ?��B     �WB�WE�4�Wp~������i��VP��.MGbC�ָ����E��5=ݹ�         F_xy����gO�l�~��_s۞ޞ��M���O�<�^zv�ۼ��o�S^wJ�����O��l~$��EGwGԔ����ih��'�f f���*  ����lX� ����5o��%���)����|q��}:9^�hH�1�X��d�uw    0��b����iql��xӌ���i�#�wct,(���s���mq�K��/_z8lz:zs�SYr@��N��^����MM/���x��xtˣ�ló���      �w�#*3�1�l�n���n��9����@�vY��w�f�7G|�I &��\v�eq�>��>����c��k�x��B1;�^>wy:�F�����  SEI~Q=���ڃbE����s
�h�S\sf��������և㾆u�ѳ=    ���U�)���4��y]W�4�> �3y��J�MN��"-�������Η��4<=�1LA�E�q�Q���[Z��ϟ�y�����G~۶o      `�f�͊�\UL6]}7`l���f��^�;�=�����������~������������؏�'�8q�fz���o��q �I�0/�V����Լ!����U�)�?���HF�Y��T�Y�H����h�   �Q%3���E�f�1�X�(��aƭi%q����h�j�_��H�d��x�����3���禣��9������?�K�^
       `�J1+����N�lP���w�|7������>����}�/*�+b$$�3���� 0%<=|�����㈾�Ey�`|J�1GN}:�b�3��u�?[������c    `d�L!�ύ�f'�X%�E��R�-�3���m[�[�oZ��m��@�KN�$>t����q���       0�$���������b��僺oGwG�͏�&����\.�ӺǶ<��?��C��y�=t]|��O �dS[X<sy�1爘YTL,�El���,u�[�-�-��M    ���I���(��]��9<�/�LJg���]xB�W�.}1�����|��������8f�c��/����       ^VXX%y%1��������()�����������G ��S.�7�y���ȦG�=�~O�����v���9�����_����5��Kw~)>���GOoO  L��8�z�8q��qL�"/�L|5����y��9�קǸ�S�Xt��    �I(f�گlv��{t�y�AQ��&��LAW�4ڶ�M/�:n߲&:z���>t䇢��"��Wo�7    ���l6��l��藗��.����ttww�����{+y.&'�'#�|���y��ӓ>';;;�?�TR9�2fΌɦ��9��UVV3g������#�i��&'�m��ⲓ/R ���9���+�w~1ڻ������q����_W�k�����u[��_����|  �AMQE�=��8e֡Q�-&�L�퐪��h�j��6=?|���    ����d�V,�s�GT�n��3�-(�-~k���'[�Ī�����;����Gkk7���v��Ҩ.�������GIv`W8|���Ƿ>��vY    �gIp���4=�o��=Ib۶m���6a-	�$�����a�3y�':::���5���  ?��ޱ�i fٜe��WOW\}���|&��n�}�x�8��;-N<�������б
I����o�kW_����va `RH.�zƜ#�Y��d�Ζǻ�)�9���ևc��g�m    `��:	d��������J'���҂�8{�Q��ه��b�sw�3m[&���^|g�wu����x��7���]�/9}�a�O���������    v/	qTWW{ f�d�iӦ���$ʑDc`O��󣲲2���FlI|&���Q `��-��U����8˪�V��]붮۫�p�w�#��,��<��اb��*��l~6��Ե�ņ����G����=� `2pTvH�y8q��t<Ҳ!Vm�3�kx<r�\ ;;pցq�[�ث9����sޡ�Ŋy+b�<��    F�P��AΜ}d�=�Ș^8-��v����3������U���� "=��'��$�/>>�s�wbNŜ�n��ɋ9�_�;.    �_iii�I0���"466Fo���ӿ�9�ċF������f�Q__  �ē��z�7�e�]k�_3�s�w�ǽ�ޛ ��,?�����y.�J��N[K</�o�������ߥ�F�e���pɈ�}�ҳ�   LlB1Pq~a�:kE�k�qQ]X�Z����> I}��g���W��S?�C��и���;����n�;v�c��Q����   �Β�hEb^���ӧ�Q�^���$���F}�;�{hjj
  `b�@ �T��[{`��b����=ٯlv|�u���q\�ܝ����    � �L ��8e�!��'���i����?��������3?��[� bS˦8��g�}�����n��C�+   Џ�����f�XL]]]zb$���X>/KKK���#:;;  �vb.���x�� ��K.jyd�����'��������ϊ�s��om���U�Z��    �k�� vbΛ|�U�C��!/N�1_{��xrۋS�Û����������6g-=+.��   ��UVV���c��(Hyyy���$'%TUU��R�� ��I  `x$�$p�Sb��9{kA��Ԓw�3�6Ƿ7�\0    vC(fK`~S����SbfQU�pKޜ��p�����ן�Il�l
������������Olڧr�XP� 64n    ^VRR�A�hkk����`j+--�������0�(yN ����'~��|i�~nu  04o�6?.��X2m^�p[T6+Ƭm�W��5o}>    ��5�G�ү����ŧ�AFR$:a�㘚7�/�����h��0mnٜvĂ#v�Ͳ9��:STP��;,�ZxTP{@,�^�Q\P�^����1��n��u�������;}l��}����{L,��4����&�K��u�����6<�my,�~��x����w���<�?>��c���d撨.�������F][]�w���קG  ��$�/f��/��ʢ��9�ڒh�x��b���  {�{�{�����  ����"Λ|�6{Ed�n0��X_Z~A��nm���?�-.�
    )��q�"[�-8>Μ}D�e�FKa^6Νw\�8cy|c�O�-��
�j�|����,�z���O���Xy��(/��*���<{O\���q�o������[7��5m�.˓��I_=i��N��������MM�>��{̛�9�p��]w��W�c8$A��x����k��}7�l���.���/�/=�)��&_�����s����wZ��NqƁg�ǎ�X��������ۻڅb   �$3��LqI�(/o���2��?{wUy�}���d��6�$a'움���REVAl�V�^�*Z�k-�����V�
EѪXq��\pc�!�=d��I^���Uf�/'3�o>�#�3s�0���<��    T}����֭Z��V   �c��%m�iz���E
h*�{Q�&��Pww�q`�^����*���1'<�8G�������    @`�b,�fӄԡ��a���x��c���~�&�����\����BIV^V��I1I�����֟&�I�:��}2���i��=p��ݲ��/���§�2b-�z��;�+����Z�}O�5A��Wy��)�����F9Ʈ�]�/#��ŏh��i����Km�ژa����lF~�|�N-8���%�K���3����7�����V���'���    �.�Ŧm6��v��^&�*��!+�$�   4;�=��O�����ۛ�V��L   ��a����x�D%h.�����H�m3X���(*��/����     �������'�]T��@c��N�S�h�^������BAvQv��?�pT%���&<f�B��f��ֱ�����u���5��iu��,۱L�Ϙ�wlt���
ŌN]�uN�>��@�(񖘫�ՕH������؇��`��!�hb��L-ٺDM��7��O���6��    ��	��f���!��P��0I   h~���c�ǘ��R����3_=�uY�  ���:ݺ��dH�,�*��^uT�z2�.�      j�5[6��آ4��(MJ=Ka��$z���rB�PO꥿�z_+�o���U�h�����~�	Z<{���z�Ð�C�򶕺l�e�l�g��}FfF�1#���O��~��m�������q�'W<Y�c$E'i@�~Ǿ��ˋ�߸�8-��@���D���ֻ?~W��}{����������m�w	    �6�(KDD���� tY��'Z   XK�3Q���ܶ٢�腕/�x�q  ��laᚘz�fw�(�C�J���\/��D���PEe���      ��PL3�w�h��s;�to�+�͉����w�]�/ X%�$W9^T^T�>��������:�U�c�*|����D#���K4��q����>�[��w�KR���.�z�y?��S[#����
�F@ǈ�x+j���n#���Y�c���xΖ�t��w^����C����K�0ߐ�k��&�=��:Gb�_     ��iX���ń4�=�>_�_c   �4z��֣�Ճ=�w6���ּ�%ۖ��r  �`�9&E��_���X�#<B?��#�ߪ���|[�=Y      B��&���v�H�[�Ҝ��g�;��=j�5���l:�;W9~�s��q#����Fb����v|�׿}]+���a�a+8��h�%�)=9]zOЌA3p?1��}��:�3�y<S��,s��PL�3A��k徕����kt=W�KC���{�n�cddf�z�C���j#1F��>0�����u �U�+Sld��ĵшN#4��xM�;��o �O~\�ٙ�׶���;O_�t���q�?���y��Ϲ��b���Jo�n�#�S��     �x�^EFF�*��	��2+=��k�V)   8]�=RSL5���,���e���ig�N  �
#�qE�9���y��Y+�T�kL�O����ᕚ��c���      3B1Mhd������ڣ�T����&iDro�i�[�.�&F$�*{s�V9~��;��KUV�_��޼Ik�9m���Hۏm7�����{�ޣ��>��ξ)`���,��HC�jFKj*cG��;�:�c���n�P̩�6d(&�$O�������2�/:��Ǎ�ʳ_=�?~�G�>���u
J�Y�i�z����fph�6p�����mzi�K��߽�XKC2"4��i������/�Vnqn��O�N2W�  @��<���j����,��q'Tz<=z����t:ճgO@u�/_��K��*�v��ӧ����L��r������7
@hZ�~}�ŢJKK�����v�����R"R @�j�j�9#����W{�҂��p�B�
   X��K�=��]T�����ɩ�48����Mm/�      ��4�h{�~��"�k3D@�0^Dv�-�s����F���c�h�#ั�uǻ%w���_�1^]��f�cv��.'�N��ެ�W�a#0�π�t��;��Ǐ��223̿�� �c��1W����I]���vy��DQ~"iF��6���!��ғ���}��S3�R���T?�����j����ٮ�j�_#(s��W��4�O
;}%��d�q�5��YjH���ϝi/M3�.5�]���w.   �\MN�4���P'�Vu?��}��p�\�zk�;yc���B�M���b\\� �����yC�[���	S�  v�{�#:�0�����z{��f4fY�2^7  A��r�a�i�ek�E/����L���N���T���**�u5      ���idFa}N�˕�lb�Q���T=�]O�|W�5_ Vu�{��vt����q�����d�]�kT�+��}33q�qzf�3~�.�_������y���>�����?��ic#:��3©�����Q�F������hJ�)rE��w��N����#}T�1#|S���z������٫�^���?O|���ʊ�������4C�-L�oRcX�c�&ϛ��v    �F�v[�����|!4����J   �y����|�0,�{�Չ�����3�m��͚�j�^^�r�ߛ  ��֑.��}���:	6��p]�a�'v�c�-ҡ�      ��PL#1^\��n�fuEaAot���A�mS[��	h�&���i�Uyc��@���K�]p<�x��.�Z�H�)�}��z���m���w܈���_h��sj�O#��/co��������^��w()&I��L����H3H����j~�n������15>��X^I�ƿ0�^��S����tn�s�I�?d�B��~���������]2�"1    �Fg�0l6�|>�����Xeeer8Bh�Z$�P   ��<�s��	���g�9[���������~��|�r�}�ś�k.   @S;7��n�6I�v��`�+����3=��=e]/       X�i�Q���c�zƥ	mN~�?��Z-؛�7�V���R@KqV���ʌW�hG ���j~����P��o{�6������>]1���������:����ψ��׹��w���4�b��6�ۨ�.77cr\J\�i��SǨi(�8F��a�am>�Y5�p�Q�@�Yz��\C�u����Xi����f�i��=��E7���@     4���p�\.�8qBVaC�������xd%�b    �ؗ�OO|���������!ר��S��g�iL�s;QtB�6,�_������S  `]N[�n�6Q�Z�*�푺��ru�ӻ�S��L      @KG(������9=.����d��ǝ~����z�7U�-`e��zέ�ݸ��a�z��n���;�]��\9�ʀ�]�u��5���|�z�5o�<��I�I�k�yk�ӝ��[�=�����?��O��>j���7ڠcǔ����v�9F�ֽr���&P5�����~Ƕ�n��֐r�s��W��Αw�6��{^�|��;޲�e�p��    ����nB1hv��n%�b    k21��>zH�;7��ꌫ�S��#����v���9�F/�y�܌�  �U�s&龞��1���P4&e�zƧ顭�j_�1      -������ѵ��(��ʆ&vדn�C�^՞�#��X�k@� ]��"�l�ϔ�J��6E�E��;��0L�b[��gՐ�����I����M&��X�P��ԣ��V���~hp�`%:�S�S�~F���,۱���#[t(��i��Ai��Is5� �����g�8f� W�+WC{�����b��cC�b^��    Д�P��X-���O(   @-TTVh���v�{w�����c�c���0�g7�G�?�w7�k.Rb,�Q��O����x�w�^����DG��{�`ll��?�|��aI=uG��c��Ҝ�zb���㎷���      -��m�ԯ�/��^�om�n=9�z�y�{���:����w�ڡ�V{�G�=i�j��ȸZ��ެ='��}L���ǵt�R5�o�^_���Ym�?�~C1FT炮�MoU��@��w|l�ט�fgƠ�Z���5��H����:�`L��)cB��.�;fL�id��vߡ����>��ic�:k����k��    �)������*�v����vb)   ��W�-ջ[�5���f�b���I9#�u�_�=ʌ�ۮ�]��z�毚o�g4�M�6i�ܹ��f��������b �1��]��|�h��(* �i��==�����w�9o      hi��S{g�~�k�:D���s�G�闪W\{�e���V�4��m��[cy裇��ZU9��YǌId�r5�EŤ��� NV^V���l�2�;�^�cF���P�=ܮ�>ɣ�W��w}��oDc~�1��mt��#Z�����;���Ј�#�Iy��ܷR�=��X���x�i�wo�݌���k�1cB     4���DY	���d��n��'^    -SNq����y�v�o���O]��衋�>���~����5/���H   �%���zNՠ���}���W����qi�ݶו[^���      @S"S�&�1#Q6� 6��3����(��$��
��x�=����^�_j��cF��1T�����k�1&�Т#N_���TgH�!���?���~���IƎ����1�V�3��XF���2�ݠ�coTc:�{�����-�ܝ����z��>�     ���햕�	=^�WEE�y�9!!A    �S��T���Z��x_xD�����G���W����6k���d��/�1TVV����v�$V�5����=C�#]XWg=1�=�u�v      �R�L]��l��e���j�@M�su���o6����Xٷ�Ս�n�7�����1���op|]�:5�E'�7g�:&v�;޽Uw-ݶ�F�2&��ؽBv�𴱞�{���]�љ@��e;�}�����ӎ�;���~�}m��^�s�>F��1��:U�}�ݦ�t��h��v��$�ر     �ILL4W_4N�B1����X���@(   ^W�|�
J4k�,M�?��,�It&��7�ۖ#[�`��[5������jݺ�fϞ-�1�߿_�/6����, �opB7��s����BQJT����:����V�l      ���%ce��u�	�C�vR�����顭�jc�V�z�j��?�����W��m����	]�e��MC1�ݯ�ؑ�7c0B0Ƥ�@E\�\��~�9u����>F��q�OFf�j#�cf���kuqϋ�?��"���V�����f����l    �ԌՂ���,h�'r���d%�b  ���r��l��6�$>>^ �����}���_�����B����ny�M�;Y3�4�;7"���;������>��C-X�@om|K�
�   j㢔A���D��lPsN�C��JٵD�Z)      ���Ԃ���=�����P7qv�~�g���c��� �9/<�U�W�]�i���vt[���:�u�1crX^I㝠r��D�����Z�kY沀c�d�@�g�Sgw:���=�����eF(�Ƴo�{�@��({�Ft�wlá:VpL���J8ַM_sk�c��K8    �<���,h)**Ryy�"""����xd%�b  ��f�)<<\��.� ��:����&k��l�	0�O7�	4���n�u�Ե��r���{���?�76���y^m  @U�C�h���0R ��XP��]'�}t��ٹT�'?       �"SCI�8=��ju�I�������S�Ι���-P/�|A+�U_�/�)�8O�%�����u`ğhGt�1#�RY�xoU���|��Y��N9�9Jt&�66:}t�۝��3��C���T���._����o���ƛ��/#�����Ֆ��9��OcƉ     �Jbb�v��-�0�5F���*��S��    �e_�>�~���mp�`]?�z]9�J�G��z_����[�ḿ5z�����W�y   �ɘ����KuA�~P�S�))"^�mSe�      ��PLt�n�G��RRd�ߴ���0V.pG���;ߣ��:�ؑ�Wֽ�lǏ�G�/iܓS�ڿ3�Y�}�*|�d�'��不��s�S��^�zd�ic����e;���<�([��V������$��)��������T%Pt����aV��Vx    @sp�ݲB1��j��˚�b    MÈ�ܰ�ݶ�6M�3Q���؞ce��t=#:������ɏ�-�јe��u�  �2�ڝz�����  ���Jt���-U�-      `5�b��-&U��{��#���K=S�Q��w����'���j�UxXx��.R���]��1�������+3p��8�C1���/��r}��3�V]&�   ���ƨC��'^���+<�qG(..n� Bc�_ ��j���U�C���o�á��m={�l�����:tH�-55UNg�!��7����J�HT�9|� 4�]����N���W����[�7ֿan�"-3�0�1}������c��jnۏm׼U����O���H   �$DĘsܻĴ���'��~�������+��P      ��p�t�Ƕ�#}g)�^�d8 uwAr?9�zd�k*��
hIJ��'��G�7�]Q�W%../�����K c����/���e��D���Þ��txS�ǹ�;���+���ˌ�㐴!~��j�*yJk�1/��w�Xy-�8G�a]�:  ��	����D����F�'���� ���B1yyyB����r� 5�=�6����،�]�*�0�σ�����
@3[��F��zF�(+/K�-�܌P���35{�l�ĥ�z_�[u��qs��Ʒ�ݱ�  BKbD�����Nѭ��t�i�?�����8_���      X�� ��:��3�E
@�;��C����.T��L@KQXx��XG����UQY�(ǎ����~���6sb����]����m�U�N��223�\%��]����H��ƞ��|����V��	恎a�*lS���"�E��{i�KZ�{�     @�Y-���>0��+?�:�    U�|x��z�.ݳ���:R���Ҕ�SQ}�  ��֑	z��l�uZ�5y X�w&����6�ס�      ��P�g���7=��! Mg@Bg���L�f��*�
h	{�;ڭ���حb[;��N�4"/ƪe?��L���Z�o��]6:}��}Tp)*/��{�6�0���Ґ�C̱�a'�n��C�CWd���L(    �:r8���Qaa���!//OF����@V���     �	c���w|ln�.�U��L2߳�m�9�   �?�9�5��5j������?������w�-<*      �����s��hN��e�	@����\���M���:#�b��h�V��~Z���Q�m�;����:�ӈ�����h���mT�}T{��e��b�c���Q(�Tl�.���������     Pwn��2���#��6^��
���4    �^nq��^`n=Z���3����wI�"  �N1)���%:b��qz��l3����      ��D(�?���I$�����h�k5g�<��ŕxK�'gO���$i�PLJ\��Ʒ8����:��X�,#�27c��g�ؽRz�v��w�!��1��.z��ct�G>~����w����c>���J����-G�hr��~���r�     @�������
����`��:!!A    �-Z  BK��$��{�#�� ��5���lݱ�E�+:&      ����_g$t�ݽ� XDט6z���������W&��6�03���F9��ϬrܸOu�����Ƕ�{���<B���ˋ�h�?F �&V�[)O�Gq�q߻|x�኎�VQy�Ƥ�	8�-#3Cue;��g�'�    ��3B1VQTT$��+���B�]~~��$11Q    P[	�]1�
�2K�;'  L�#]�ۏH`����s�~��*�      ��}R�����t9�x8 +��^���ڼ�B�UzX՗{�Ԥ>�����5^Q�(�xK���L8f�^���؋�P���0B.�x}C1�
�>���&����#�f���<Fm��ϊ�+���~z�as�iцE     �g�@Fee�<��v?�y���%    �	�}�]G�q���_n.�  pJRd�~���j�  �q�k�W^���\      M-��(=���H����9�z�H�_��B������>V�����\f�!�#1�]�����Fd�>223t�����@����
}��Z燡�S�0�����{���\}{�[Օ��|�纠�~�猜�77�i�L     j��v�J���ń���|Y���PLL�    �*}�����35{�l�ĥ  ��\1����F�7`E�#]����j��)/      ДB:�9&E��3SN[� Xװ�����T����`5k��jω=����w܈�4d(��C���؀�7-����g.7�����O�m�z��4W�ic�֙��
�1����������_E��Q�.��~�.�y��l]"     P;III���#?+�b\.�    ����T�4C��F}���׾�9
�W�ׁ�  �'��G��R��V`]�4��5�s�<�{�      4��Ŵu�5��l�ٝ`}�$��Ͻ�d�;�������3��㣺��e�.�?7����J�I�>p|�~3�R�E�����n�ic��kJ�)~o�lǲZg��M:�9r��h��iꀩoW���c<_��{����r�ǉԊ�+�_b���     h	�N���
�A���˓U$&��/   ��/���_���g꒾�(�Q�}�xK���w�Қ��dےz/�  �)���#}f�[L� X_��=��j��8O��      �BH�b���z���J����c\�!:R���|.�j����1�9l��Fx���;<�71�yşUQY��2b,�B1�p�~y�/ަ6�����~���]�u9�?�����O�[s���;޳uO-�j�&ϛ� �'     ��e�AS�x<����   ��ˬ!�4c�%E'�k_k�1�0/�y�\�  ���wv��qi�r�<�5{O�iz`�+�9     @��P�=̦{zNS�3Y Z����XY�2��`%�h��y�����wrw�;׾����،��Žc��5C�	8~���iF����;�/TS�-Պ�+�t��bÐ����}����g���a׫�����	�'��i/�7o��sV#�c�7��X]���     X��n<xPV`���#��   `���3��O���ғ�뵯E'�h�"��˿�ۃ�
  ���^��I�����]�u�H��Z*      ���T(&,,L�H�D:@�t��8�,_�sw���>�OSL99���Z4k��/������fmE挜���>\���z�.yJ�#�R�+����������ʋj}�e��jw���~UJ�%����ʸ1C�p���a�mh�KӴ���9n|T��x�~y�/սUw�?H�
    \eyyyBp+,,���U�   B�3�i.Bb,R2��hs^K]�*|Z�s����9-޴X�r ��1.�LMN& -ץm�����}�k      �)�B1�;�֨��e���tO�i����u��� �8ZpT��s��~��^g\�qZ{�Z��_��-�+W�WJ/=w�s:��9U^����U/�����_�.�������bω=ڙ�S]�������T�]�����o��6�u���wl�?��C�}�6�X��$:5��$]��r����i�     ���v�*��k�E�d����   ��f,�b��?s�L]u�U�������ݦ���k���:�9"  z�&v�ϻ����Ʈ�XY����*      ���L(梔A��V���X_�=Z�����?���BV�`�sB�ug]�:F��k�6'{-ڰH���ҡ�C��v�v��G�NӰ�կr ZxU�љ�Z�cY�C1�u�s���b2vd��=��#j�j�ξ!�u��v]=�js���wf`f��ڟ�_م�:QtB�p��	�ޢԳuO���s��͜,    @(�R(���@>�O6�MN�GV���(    ������>�J���J歚�o�}#  ��c���=�`~$�N~���rݹq��y�      h!����[�M�����{{]��6Η��'�*n���j�J������!�{��[�c-8���c���223��EV{=O�G�����q�v}��3-F�1��ϛ̉xw������h��ܪ�    ʬ�1ºFH$!!AN����
�á��h   nu��TTV諽_��,\�P�e,� @�Kr����3es@�p�G�^W�o�Qv����      A�q;�tw�����Z(���w�O;_�gv-`�rM{i����y�<�ю�y<S_��mG�5���U�
J[���g.���[���㤭���*��l�25��sޟ�=9{�ǉ���o     ����X3�QVV&+ ܬ���   �p�.�q�b1���9{5�|�_=_{N�  ����~w�+̹� �����^W�W^dAT      4���/����@л����YpH�V�U���4��YZ�o��h�M ;eцE����S���bo>�����W��>��q��s����Z��mVy��Ŝ��/��Ow~��N����r^��S���}      ���MLLԑ#Gdyyyj߾����U�   Z��i�5k�,M0M)q)��W��T�l~G/�yIK�-���C ����e��X"���3���?������      hHA��Y�q���@H���D�.<���C��/�һ[��#?�i��+������u���{[�SSX����PLC\2vdT�����';?QS�rd�������g��y�FtѠ��Vx���aN|k�[*,+     ���v[&���//#d�b  ������N~�[�v�� �|ڄ���3N��w�c�wC��WJ/3sՠ����^���9��|/��5/+�([   ��j�_S���7���zf�A}xd�      �����ѭh\���M����g��-�GAi�������ٙ���9{u�+W���5C���P��=k|���\36�p�B}��CUVV�����]�h�#�x��D[�n��q^��U�F�?�9�E'Ԕ�����h;�|�&����m�����F���|��8���t���o�돶�������    �)++��ÇUPP��"^?�!�ݮ��h%&&*99�ֿ����P�Ux<��=�f��P��
�h��s���D�>��a��IIIQ\\� �%i�����ٷ?|?���u曆m�v�7��`����m5u�Tsk��C��h�X�����_���o  P��1)�-}� ����;

      hA���F�u�$ �%%*A��~���*�t!4.c��ݠ`�+{����~sK�OհÔ�*]:(�� ��a^/�$���_��VmTEeE����w4��z�js���כ�=K�+ʥ!퇨{�����v+љh^��[�����)�0[��3�@���f,�!=��3   ��(..����a�3SQ�<�_�4N�S]�v�g��.]���+�b�������/� �o'N��ڵk�e��Ϩ��W�^�Ϟ֭[   �x�wr�ɚ����+{x����*|Z�s�����M��=a  �b�N��k�"�# t8���M�+�scA�r�      @�](&�����./�!�,w]�v�^;� +;�HomzKhY�̲��    ����i���Z�l���ʄ�1;�6m2���d]t�EJOOj.11QV��x��TTT��r뜌�r�ʌ~�����UVs����\}��W�fD�.��b�j�J   ���h-��@�{�W�=����rd�歚��׼�Þ�  �)#J���)5�:�u M�ud�~�~���
��     �ނ.��n�&�:�4�YGi}�.m�     @�����+���Ç9Y�!?~\.ԙg���c��f�	�s��3�=//ONV� Y)�����ݫ�^{͌���v�ڥg�}V&L���  �����є�S굏��|���m-X�@�2�qR'  ��	m�j��� �.�{��6g�C+      �GP�bF�ꯑ'7 ���9=.����UžR     ����\�����'�U�V)''GӧO'S.��|�|>_s��'���"�a,�p8���V(������[��=�x�^-^���<?�� V�n�VjD��MII� 4���8�k���K+J�=M{_�X��~N�.TaY�   �Ct+����뻌զ���SxD      @]M(�U�K?�:^ `H�r��c�x��     eeeZ�p!��F������_�&M�fDY�����wE��E||�\���d��{(:r��|�M"1�h�����W��,��Z�(��4SN�QH����������6�����ڗ�������;  P_�v��~�"�# �0���1U��{Fe�M�{      �OP��	;�qG��kw
 N�f�����g�7	      حX�Bǎ�ڵkկ_?u��Y����D(Ɛ��O(&Y)�����P�t�R3T��SYYi>����r:y/  �1�zK���w�Қ��d��*! ��sM����* 8�Stk��8Z���@      @]E(fz����Ť| ����Dm����R�,     ��������_M�/� SF(�*�P����W�˥P�w�^�ٳGh|���Z�f��9�  ��l9�EV/�+_����  hh�\�4%m� ����kr3�.w�      ��j���4�� b�N�"�Rݽ��檛      �h���*++��G�z���[�K��J���<B���J�������[�
M'33�P  @�)�����3_=�uY�  �X���wu�\a'? ������~�n\��<�b      �Ѣg����u[�I� ��	]tQ� ���     ���,�锗�����jӦ�Xbb�������J�+}�7~�4�C�	   uSQY���=��sz{��*��  ���))2^ H�#N?=���v,      P-:3��y��* ���۪��.�Ή      �ĉB�2sB1UKJJ�UX)(�����'�p�\
5��iZ���***Rtt�   Psy�yj�P;�  @S���[�! �����c�6w�      ��j���v�$]��<@M�آtc��ȶ�     lrrr���c^������������
�� TRR���2YEbb�B����4-#�C(  �v�|eDb  @�r�G迺M6_���+n;�=�uO��g��=      `m-2v����K�k�w@397���'�җ�[     L��Ѵx̫g���r������w�PL�x<�
��!�өPbĲ��
5�㞖�&      X׬�#��� �TJT�f��@/��P      @M������3�7�� ��~�u�6��Q��X      ����TEEEB�2N�G��n�%B1FTĈZ��k�R�'11Q��XV��q     ��.1mtI۳ �uY�����&�(8(      �:-.����c u�>�=��'��<��]     No<�5c�����SAA�����`�PLBB�B���2      벅����Kd�	 j����Ku˷��[�      P�����8�ڣ uuq�!���:m�     @K����#//ό��lL�����Ux<B1A�PL��gO��q     ����g)=�� ��:Ǥ��^2To�J �+�2\EEE    �������6-*�'���I�- ����03:u������R      -YNN���וrss���$f�P��iۖI����X���R��gO�      `Mqv���p� ��ft�e��+��`U��g    hP��嵾M�	ń�����83�  ��3.M#[�W���     hɘ��|�ǞPLլ�����������D�~�4��������p   Թ��zm�k�����Z�P��LԜQs���6�_5_  �y��4F��h@}�ڣ4��(=��=      ���P�ؔAJ�e�O �'�/����W&     ��*''Gh<��3B1F ������<�<��IHHP(�����c��III   �1�c���VkцE�k�]ڕ�K��as��7���7c1?���  �G��V�2X �PƵ������#      �i��-R�:� 4���x]��-ؗ!     ���ĉB�౯^DD�bcc-i!l\�	�4���\3��A(  ���8��S5��$�훿���A{s�*XEGD��C�;Gީ�	�  ��].�-,\ �P�O~O1��ܵq�       ZD(��(1"V ��.O���Ց�\     �4^�W�/��q�>��v�-�����Cyy����e�CN�S��HV���  �/������~6�gzsÛz����f���833g��Ƨ
  X��^��M ������c���*      ��,�i�tkr�a����Џ;^��߽.     ��&77W���B��d��1B1{�6�j�D��������D�"Y͋�  �j�a�:`������ۖ�ٯ�ՒmK��%�ۦ��v�f�9ی�   밇���N	 �u�/����l���      ��X>3��h�t h,�%�ћY� K      -	���e��o�z����P�x<�� a�PLBB�B?{��?  ��UTVT�;���k���;�W���yA�r���#�u��+�@��Ϯ�m�>�  @��f�� * 4��(����C+      �'K�b:ƴ����
 �1ihF�t���     hI�P	����UAA���Xѻ*������***RLL�в�i^�J�?�  �-�8WC���/}ZC;��i�4�����mˑ-zc�ze�+�~l����Ԙ�1�:`�.�{��"k�Z��8<����j�  @�q��ue�� ������#�TVQ.      �K�bfu�0��'��w���zƵ�6�~     �������PLլ�1�B1-���E��y�������f�	   ԭ޿Zß�ϾQ�}X������[�_x���9�Fn�P�d~�/�|�²B5��p�K�]Gjt�h��>FQ��߾��B�W��]K�ұ�c  MkBۡJv� ����m�譃_	      8Ų��N1)��K �Tfv�{6-     @K������t��Q,))IVaFRSS������*\.�BIee�*A󩨨0��Y)�  М|>=���zc�f,��3�U�-�F��6���u��}��f�7���Fm8�A[�lQ���A�g'w'�O�on������*9&�N�2�6�|��}  M/����v� �ʕ��ӿ��Q��L      �����k;�Q�� h*������6��     @K`DJмx�%�ө����+f\-_^^��"�b*+c"zs3Bq��b   ��h�Qݰ���?���Դ��^��q�s:�cn�x+��}b���?w��߃��xL~I�|�>��(��H{��"�d��M\��o�v�vj��ތĸ���\��N���^-ٺD  ��LJ=K��X@SqE�hB�P�q`�       �%C1=��t����S|��.�/�-+�xʋ�T�(��=�e�U�T�|�^Q^�<|�6�p��",9�����w�m��0{�3��6&���e�Nt;b������fv�;7�     ��UVV*77Wh^�������VVVVs�y<���󘐐�PB���K�.  ��vߡ�^�G3�Cc���k��OF�%=9�ܚӖ#[����o�� ��m���i#���2��DyA��[�]�-�*��.�,?R��ey}���u��+�l��
��>[xxDEX;��v���=,�m����fK��;��G8���1��8���5��9z��*�J      X23��(!ty+}�_t�s�8w��[���[���2����.m��^g=>��#��8��c�N��������f;���������T�ӧ��V�@A���c�i�o��>�Ev�&����V� 	K��"�Yd�d�$��m�~�3��*$�����s������dH8w���;��~�:'�k^6+�>���b���wJt���//&w
     ���PB�\��h��X%�L&��*����K('!�e�{   �mk�V��΋eA���W�eg^&a_X�Ov�D���^{�@  �igI��X�)0ujc���P�/?�k��y1].��(���\�q�˻��h�'����,��ϛJ\�9R�(2�����ϒ���"      ��b��dE��sTkUٓ;��;z�C�콅b��w}a��S!���G��ݨ��ޟ�xከ���3�h~S炸�yr�BC��s�      �c��5M���Tʐ94�T*2::*V���i��X�  ���1�C����7��\����U����\��L!#��t�\��k�  `~��i���凋�3/,��KW�w�sw�Z��W>�
�7�}�����	�n�G~wns�i��_�jt����X-	      ��r��O�8[`�jY�H���=���R��w]��M��o����؍�Jww�����O��cW��2���D@`k�Gȼ�Nٕ      �b��5�r��5
	��P�J:��Z�&V���i��X����a	��8`8 `6�����c��������z���3W�%g\"�:�S�n���l=��i������?�v=  �����$�k؛:��st �+3��p9}��k7>!r���������W�̵矓D�0�����M����fX���mц��      �f�PL�?"�/ؓ:p�=�;�c���C��?�]9��������w߾�e߸��]��_,��Y�5���r���ϖ����     ���$n��Äb��*��d2)hlVZ�NŨ�̧������ `��p�4�7A2
 s��~ijz���[��an/��P�~��/��.���a�Ȓ����l�%[��#o>"m{Hx�ٟl�aT  8��o||�{��[*��޿q�8�w�y�a*w\�ȓc7�*���+;��>1:�C�վ>1��䡾�&ֈ�     ��
�\<�,�<{�Tr���=��d��Wm�(~��!��l�����]�Y�<�����r^��r��Gd���    �51Y�:Ժ�>}��Ȭ�)�˒���4�t:-V���i��YC�T�l6+���  ��˕rr�+�կ�Ү�r���e嬕��¶�S������<��9yrד���'�P.  hg�.���6���ky9�{מу�v��7H�{;p�1���7�����/.�̞�s[j��ӌP���X,Om      8�e���<����}($K���@-uŷ��x@l����G�n�R]/���f���uyl��~�O��T��c�Δ;vo      +b��u�.�M�^��X,�}W$�L�i`j�YE4')
���AE��   L�W�_�_���|�r���'ssen|��k�'a_X"���Ai4K�R�L!#�B�ٟ�/��vׯ��v�+�����  ���8[`�J��5�{�|���W��[�<x��͍���4-�z����s[�aΊj��y6�      ��L(��]+��4���p��#;n}i ���ݛ�� ��ݨj"�}���6/�q���R_o|�Z)�����@H      �FM�5��D"!���f�I�R���%hL�tZ�"�������>f͚% `�Z�& �SM�ow���lޱ�~  ε�y�,��4�ty��BrǏe����?: p�U��:vsޟ�ta�O���&���6�Ė��-�#      p&K�,<.�\<�,Ac;TL�6��]��k�w�g�iaMp�6�8vsڟ]��Ýw�[�D=�јT������O     ���r9���k �3>V	�X)4��S���F��$�b����lW�x��Ć��� �}��{�wO��;�oF(  @�Č��-_-�~:���ʡ?������߷��x`�����M��������<�b�j��O۾+      p&K�bV�IG &hL�JI�~}˛����_�0�R�ܹv�c7']zÇ.Z�<��%��킆��i�����x     �R�n-���Q�+�Rhg��$
��Ų� ���Omm��4�}�֪  `q��ݶDИ�{���v����{w�ѭ������৯�`���+�OusRԆ�[�K���"�EN�      �D��\ԵBИ^J���Fn�ŷ_����p���4vӱ�Ə��{ZO��V�#h(3B��,2G~��-      V��pkI��R.����!wˊ��b)B1�*��*�g��bY�     �xt,�����h���Co~���=�m�;�u��7�nN��u������	w4	����ǶQ��yB      �<��Zo�Gde|���3է���u���K�1]����ޒ������j=�,���Ý+�      KX�:#�������,�H�$�IAcR��L&#V�F�i�X�8      c�\.�P���R����m�葋�w?\�
��]��i�;�i[�����4u��{z~,��      ���Ṗ:O��兑�o�����ݫ�/��\�����{���#W�Vb�u큨�?��9�K�Ɲ$S�	     �09�z��UB1�TJИ��T�U��x<.NC(�Z�٬
	     ��wJt���
ǎl�š7w�U���ms���f�?�>���؂�4M�´`\N�͓Gv
      ���P�K(�7��J����+7���?\+���Vo�9}K凋}���/\"�<��+�8U~���      X����url�HD�^���eS����e�u���I��V�z`-*R���%      �z�:C�*��<;��������4*����n|bG�y�+��󾎥��uy�wQ�
B1      dj(��	�p�@�F�+۟~6���Z��s�����?�7vs��7~�t�rE��Xۇ;W�     ��&��ZX'��r�$����M��bQ����AAc�R(&������H�VX�      cD�a9;�� �p1]�r��+o^��:�q�ܽ��Y�������e7��-�b,Nm�"���J4�      ���P������m��[�~��`J]���Wf����e?����5��SNl�)��=     `�R�$���fhhHpl�D��P���#�bO2��P�#'agM�      c��y��ܦ��8���%�=�ƹw�ѭ�)��;����hY����̄��Զ��������      8�iG�[�!Y�X$��r�"��z�]��s�՛6Ԯ�,:%�����3Z����     f�Z�&�&돏U�*8���!h,�tZ�"����}���     `�v�&��g��غ��s�ݟߜ��ᾳ2cdh��3�NX�      �1-sv�I�uy֔�j��^���>��	w����|�����p��U��K��޶�r��R�U     �,L
�&Q��%8�D�'��Rp�J��
����B!qbX�488(      �Z3Cm���K`M곘������������!�S�������;�����X���m��p��=(      p�B1�-X�`1Uy��/>q�ڇ(������ϺO>򾶓?(����IN�Γ���      �0Yߚ��r=b�FG���
���Xe��b1q"e��z     �z�3�ݪ�ղ<r��_�ƕ���V�z��>^�����;���6m

�✶���      �`�Q��/,�F�	��P1U~��/.�c�ÏL��?_~�����<�]�ه�F} H(     ��P�u�uC(��Z[[�
R�bR�P�i��XS2���ʼ^&f      L������B�$���7�~�_�P��������-���;� w�y�)�b      ĔQ��V�q���[*lz��o�����T�v���vK-w~�i�q�Z���[����r�"      fX�Z7��I?��x<R��{|-�NK�V�L&#V���I�c?22"��nT,�*.     �F7;�.s�:�2Z��xi�-k�Q`���n���F)^�qڍaO�X���
�շ_{�      �gJ(�Һ��GJO��r�7���E�%����}i�)_ر��.�8�UD�a9-6_�~S      �044$�&�ͱ��n�F��?VD/��訔�e��H$"N�J�,���T��P     ��x_��k)TJ������e�"1q��7�n�/�8���;� w9�m�|+��      ����b�f99:G`��Teˁ��������_�ߗ�oqG/�8�����     f��j�L&�4D(f\���U:�4+m��s�I�ضY�     `꼷u��:�Ւ<|��knZ�����|�Cw�nt�?�q�MA�_`�S��=�b      �@{(�춓��r�a���>z��q�#O
,��.������$��v�K�����=R�U     @����T�?&�r���sϭ����p8,�@@<�1��T�V��ǡP(H.��r�|Կ��+�����_L��D"!;v�0�>��y)���3x�QX)����IԾG�U�V��+G�^����|��~H��Q���P�������۷~����      �on�Cf���P�Uec�����5�.���Vo��{�g�E]+����K�j�yM��+;       �7�U�EkP��͇�^qǚ�X�W�|�����X�X�L`�foH�Df�/��     @']����y���577������k	�0Y|Z[[�
�ɤ��3�Q�R)�
��btF�N8���ZZZ���THFG(�H     ��X�X,�������<�-���V��w���s/�\~��V��     p ����+'G�
�W�lx�_o^��:ACغ��"�ٻwitv��tg�O      ��5|��F��7:
�f����$8�x<.V�N�	�4��� ֯N�k����,��]�B1      Sce|���:��3���{�@�����i�m��Ӻd��tg�m˾��c     ��iŜ�+!�}x6�'��������a��^_����B��D@`�3���ݏ     �N�b&GW(F&s�DB� �L
��ȈXA,�a�39�PH�r�~�V����      LN��%�Y��;�����
ʖ�������'������li�%[�      �Kk(��u+x%��?��E"���?/�/xm��=c�!O��&��V��q[     �j2�v��Ũ��̙3G���A60S*�4�t��b�Ѩ8��}��B1����r����D" :}:�i���j��^�g��<gzϔ�>����.7n   #,�.��#0סb��ux�{7wo.�Zg�����oy�#�	L�q���|���      �����1[~��rvߪ;�o�
�mWo��1|�G�����4j"ˊ�	�q��     �����`���:]A�F��z�����P�U�#��E�>*t�$�\N�y=g�[������b�h��Ծ�P �®��k�����. ����ma�������  �8��|�jI6���w]��MAC���6�
]���G�����c&�M#     `o�B1����
�	�S�U噑mWܹf�>AC���^�yG��|2e"�"     t�!�[(&�7��P��$	��)��G0>VY_�hT�DW�L�[(FQ?��P�ZOs��      LΊ�	sm9��wo[��{��v��~�>vk��>�~��L�2��~R�Z�&      �'m����Es���+o��;����w��B��@�/0���q��&`���Γ����7~&����j�v�eChÄ��2�2Y=g�<��3R(&�o�=��%�eB���������'^zBj2��z�=��O&�o>�����"����w��y>�����%�K��)�ܶ�&��W}��/��    8�L&�e��b�P����߯���
��޽����L&�!��I�T+����$:�Wv��(*��1$R     0ys��pV �j^K�;��w��|_��½������ޓZfw
L��ȜP��=       �'m��Ӣ��ّ�K����Ʒ��x t�w���W�s�����!9�y����`�x�.�GZ�.��m��W_^��bub��Ү��l��E-/Z�N�LCՉ��X-���I�:���2��\���Z^�    8]�������v�	��ZB1###�c�Bl#�J	���U,'��1�ɲc(&
iY��� ����qG�n����h��D"�ܾ�.�  �)wZl��<�R��ud����^�Ym����z��?+��R�/� w�,۶�     �/m���"��(U���?^߽Q�醡ͭk7�6m]�����x��K#�	�      -tMW�<�؍��#��d�A��/8�D"a�]�\.'�RI|>���ŘGg�D��FWl�P 34�4I�o~�o�
 s��w���y��  0��8P��'ï�t�U��*��ۯ��r�-�uu��\`��ƶm?�}Z      `OZB1ӂ	I�[�xj�M���x���ި�~hAaZoG �l��2[�/O	     ��tMoi���P(�e9�ZM������Spd���b*@b���#K&�bj;�&�:�ڞ��v�m���3�     ���Z8�Y^K�;���p��������n�����|hf�e�9      ���9)�t�����/��w.�|(~C�?���U��F9�     �C�d���f�#�?��c{��Û�PLcH��b�hT�FW����I\.�؍�PL>��\.�-�     `����"�
��l��w�{%����4m����Pu���eZ0.}y=�1     @/-���j�f��������Q��ݸ恿_�ͮ5K"��Zq     �s���<�k]5�@ P�e�YS�
�������8ҥT*I&�Ѳ,��{t�b��1c�      `��n�g�_�r������k7>1��O�i]z�@�%�ٌq     �)=�����^I��a���,p���{�paˌG�.�@���9D     ��s�����u�\��U�K$��b�ɤ�����F��$j[V�մ,���Y�Hg(F�/B1      �4�w3ӕ}��%p�����g���#r�Lm�;�      �~�4{�2��]�W�V�W��>-p���nzt��/��X|�@���g�#/
     �Q
���������А�����۷����N��g�PL,'���k�,���J�b����      Lܒ�Y�~:���ߺr��#|��͇�����F�'|    `�2���w�}�T�V'|V?�C1� �k��^ٹ��5�H�(;������R���sRt�      I�d}B1�O��jd�D��`� 	��*�Iō�DgxĮ���U���R��     ��&OP�;z�凋�
���R*V�G��3�����Q?�s��     0>�`�T�M�c|(fa��^�ZEve�.8�ݟt���;���ĉ+��	�K��|�(      F`������x��mdd���<�B1�dR`m�bQ
��XA4'ѹ�k�L��ѹ�      �`A�4q���^J�顫��A_hs��:�����/�vƕm�	�ն]      {1<Ci]��w���M[��w��%+����@u}v�]���      #������tM֯V��J�$���
��+�|b��8���e�=����     `�:z��
/���$p���:5>|�`ܾFZмp�      2<3��K�O�V���_8�]_ڸm��/�L,Z&�F}`H(     E��簾&�3]�E�3B1Gg�P��訔�e�z���d��O(�`0(N�+R�r�l����Q��g      �7/L(F��S��ks����Ժ_qK�ӂ�?hC�zOxJv�v���z�]q   0�*��Zt����v�ev|�,�X$'v�(Mc��y\	{��$�	H����C��7�'�������y�UsՎ�Wj���;�����]�v�ԕ���D���#�n�L�?��I^������8������6����At     ` ]�������t��:�?���T<A�7���i�A��S��%�5xw�dR� ����׆��^m<�ؕ�}�Zg*R���.      86�	z%K�ա�N��p���ڑR�S1_��5�� S+UNI*�X{   !�wqc��/k]V�.m]*K�K$�3�e�JE2�L�$e�T�~��h-*��q��|�o�YEc^u�\?�}�T*=��/~�_p���m�BzmO������]�i��o��[�3M�     #���:���A�It��it*����k�}Pp��.�x<.N�"1�C`��	�BږE(     `|\c�9��z1�s�]_�<"p����Ԝ[[��۾��-ԶNm�jR     `>�91~�,I,��m[����V�U��r����@�A'z��j/�\��Ǿ~�T*=�v��A��343/L8A���H���ʯ�<(������E���@���.q��]��2+2������ߜ�A�5�:v�T+R�U�������x���z����7�SV������]B���y��ӟ����k��c���>3��(d׮]������ۂ���^^8�/o2�#�ˬڬ	����&ٳgϤ&��:YN��0��%��'�3��t���k'����/;]���>Y&��J�U#�L̔�`�/�<���ͫ���73���c������������b���   �Jj�����Css�ؙ����O�S��C1�^_���bb��8��ؕ�C1:����|�     0�C		z�=*��(}I�1���k*m՟{8!�j[7=���y�    �[{��ׂ0��0j^����0L6���aԭ��T�Us�[�=�=����^���Δn��hL����&B1:��ڻ�k��ㅃ���_}O"�������s�%�K��"CŴ8էN���w�{�ԛ�N����M�m�������\���7bp��~�2�;w���m۶I$1t����`P�n~��q�ݻ��M(   eddd����C1�	{N���B#kmm5�.X&D�w�N[�+���}�3�h�d)     Ƹ��Zz_��W>�s����M/�r����Zf�B�d^s'�     ���� ��&�	×[.���_UF�N���j�*Keq��z�'?v-��`�]�7����Ѐ��0��t)�*ҟJ�� o�ܽ�|���'�۶�<��ƶyN�؉zd�]�`o�b����!    Ǧs�~SS�ؙ�P�����r	�,��},"���JȇP�q���Q�Ǆ��     �c��ڙ�E�_�3;p�I-��J����=)�
     8~j,،��(�H�׃0*ctF�?+
��QW5�t*�VG�1�����0c��B�kS�?CC13B�	�)�����K�	�+��#�0vs�@�i��������L&#�թ7�R��e��$    s�����,v�3�~_�f��L��B1V	���%�I���b����-���I��-�`�����t�7     �F6�1�ڤK��h8�/����s�m�+-�0g\Ѐm     ���k�b'ԯ�b�~�u�k�xd5�9����9�(���?W��)]N���݅ݲ;��U�a�ˌAk��b�.���[z���o~�k~���Z4:;ܮo��u�5Q      �kҷ��m۶�K��@@�R�ԃ���S���]3���J$�=��xX%D�wR[��D�Qq�����^��/v����b1:��Q��Ծ      G�`��.�e�m��3��q��qk���sn���"q�"��:�    �Qy�^��2KD����zF�No��e�j|�:9��
�Lu�X+����zfW~W�:X4.�B1큨�]z=:]�Z�d9�O�����ͳ���3`�ُ    ��蚬�&�X�R*�Ď�^��A��rZ���ݬY�G���R��̒J�֤֍���фB����ItE������]�=jߪl�|��(��_�b�   ��СC��A
ٲe� FPg3Qg����n�]��X!'|M`�.Ƹ    P��0���zf^d�,��u;?:_='�T��TF�'S���T��+T�S�=�=�[蕾b_=S���aX(��>۳}��\�q� ��@~�ڱB1t��!     0�����'�؝�P�N�!T�������!��+%�:��qZtC�&tśT�����'TG��!F(   p<���|����x[�n �[�.�$���e*�����x�P��l%��&O�%0T��\���    p�X &3�g����̼�zF}���7^M}F�Q��TGaF+����O����0{�{�@�������X��b&�t�	����6m<��?�����rz ���"     `j�j5B1SL�ϩk�5�D"aj(F����4aR�ڬ w�g^:#W�{��Z���      ���`L\B�B���}���R����g��K��{rt���ԉԶ�'wH     ���?"3�g�um�!b~�i���0���d2R.Om�5W�Io����Ga
{���Gơ�tP��H9}� G�{t`[G v��PoX�ހ���D��v     SK�+��C�#q�d�P(�mY:c�L�b̖J��X��ZA4'��
��:N"e    �ŋ˶m��_��a�?� Fs�14.��P����F���0���2�O��$    h�GZC��l����׷��w�C0ӛ����7�>
�z�pF�N�x��Ҡ�/엞BO=���{�aƅb��:��Y����n�$�Q�'8vC(F��@\v��ŉ:��l2�����R���\w�u�3Z������I�l�rܯ��˗;�L�   �/����~�>0�Ig����c���T(�c��ⴈ��ȕS"e:C1D�    (+W��_ ��w}��7p��z���@�q    ��.�w�|��OJ���? ~�u�3�y�*���������멜��A�z���˯s՜ Gc`(�Y�f�ғ�+�1d�;k��_�\.��:1ٙuf(&�
ϱ����)��T��zA�x81,   �b����9Y_�~�����v�Z[[;B(ƚR�bL�3r��:v��l�b��e�     8:5��;P)���M/
pw�y��󿻼��6�o�"�    ��E�E�k3�>�j��x��Q��a���U�����_����/���`}��Dv@-�k�P!�� �p��y�w���qm�x�m�x�8�����d   �[�L=��#>�OJ�����BWW������wA���zŘ�}�1B���P���     @#J������P1N�F���#s�����    ��*�1\�|�����j�:%�PA�����[蕾b��ߺU��jmj�(��b"���x�������Ю��ĉCE�l� �x�P   ���k������%N�~���Q�P��E��z��R��vFFF�c�P�z�:	�c��Yՙm��l��      ��Z|7�a��~F�q,��se��PQ�}     )���qT�"0�+�K�x=s�*����A�C�C2P��aTf�̉���!���#a�sv��X-Ir���a��ya�P��"^�a*�xh�b   �_7<���'M�W���tZ˲t���b14�>�z>`�T8(�͚}7$
9�x�:[���]��^��ia9:�Gj�C(��\��$    {!��G�4�#�!]�o���Cq2T    �ݨ��v8��VA����M�BFb�ظ���ZI��d=�W쫇`TF�y�4$ձ`&CF_F|aG�}�,}������E�![��x��SC�1��9��b   �_�+�>ٹs�̚5K�:�,�+?ذa��r9m�Ե]<75�J�֢�=V8.���N�3n�֯��,Y�D�-[��   �cIDAT&v���'O>���J%m�T�q�̙ FjK�I[�M������\*x�����K�Z�.   �-B(�p�ZU�J��è��`MjDi�6	     �BE`�x+}Q����χC0���B-�0�JRR唌�G޺�����åa�V�?�p4Ƅb�kq(��/�8e���j���D��ř&�^�H�(�b   ���b&��&�?8Y�t�L�>]�R���Ȉ��:�����U�o7oƟ����n����F��$:�V�5���H$l���x<ڣaD�      �,�	�_)���a> ��|�ʍ��βRg0��H    �����=���H���d>)�BF*�ʔ/g��v9X>(��Q���PL��H�G�	0N�y��}��)�V�!�{��� B1   ��0c��݃j�~KK�� ���'���|�d2�D�`�P���M�̈[�b1�33�CD�  @#R���3�+  �Q�.�4y�d��|� p���ƺ�i��3���&w�u     ����s�+��1$%��E�VxM�	.f2��{��6ۿ���� �G(   �L�7��u(��d}���K��h���w����X�UB1vh�&3�Vv����~	�B���-�P  hD.�K|>�̛7OJ���޽��  `ʵxC���X�rn� 0����!c �;�����     ��g���P��J�%& Y=8vc��>&ja�7��8K � �k   0g��SB1{��ն<���
����
��
���I���'l����:�@�
�Ř�����s�D��ۆ�
 s555����eƂr�����#)UJR�  �xE�!����n& S.��Y.0T�&     `��b���x�j�& [����,&��o�U�U�n��~��B�    ��鞬����vgF�AM�'stj��M����� c�p8,>�O�.�K���e2)���l `��<.�tH XDG�C.=�R9�����O|]ny�  8^!o@`�|�� P�^����P!�@      �0$�s�ů(VK��m�%�䫥}Cy\nq�]�5�& 0Y�`�P    �'�B!GL(�D"ڗiF���x��z�hddĴ��J��a���NQ�T$�Lj]�SB<fE�:;;  ��͉ϑ����5�F�}˿׃1�r^   &�'��JR$�	)Vʯ�u�     �cB1n -]�U������Sы�b���g�`��=)	   �"�q����9�d}["�05���b��ᔀ�a����x�SB1fD��   ���]�|�/�W�����M�'   ��0�]�bMv0�jy��p��     �CB1����-�LP�Z�'0�O�b�$���G�b    �+�˒�d�.�)����9uG�
��ܹӴ�R)�5�c������)����V9e�c�s�}  ��r�,�lc,  ��ː������M&�]�����<      � Ӡ��b^�	*��{��{��� `��    "����'<E"q�h4*.�K���d��1;�A(�:��T�U��F}{�$jߣ�Sc3�8f�O   #���ox���_�l1+   ��u��*V˲����`r���ؽg��M��H<�      �aȑ��P��ʵjI�	rWj�t��#|�8�8�<�b    s�"fLb7��땦�&�d2ږy8��582�C1*N�z��D{�~N�fFX�)�3�8D�  ����)��s�lޱY `���yٲe���}���ŋ k#�`�R�ĠOLJ�V���ˇ4��      �aL(�H��V�e&�䩎
��SˌP��������իWp�-Zd��53�-�b    s&�;)���:C1�r�!�D"�#kmm5u��j���hii�K�^��������8�1�B�P(h[��%   ��/���u����(�������޽{��bV�ZE(h �q7^�Z%�I)�*���qBh      �0�f�%�`����$�<�]osDo|*�a��3�8C��e�	��b    &�M�bzzz�.SM؏�9*u<F�1#|X*�"cj=X��Z���=v
��h[��ȈT*�x��  4�]C���{.�Ƿ?.   S���N�U�B(�R���1'C     �C�����0XM8�	�U�%���.�`�91�9�    oEEtsR(ƌ�U�̙#82��/MMM�ɘw��d2)3f���*�'EL�qX���P($�@@�B�{t�b��j����  h|�ZU�����_�l1+   S�%�q׀A����0`�hn��      �aH(�R���r�H�c�j~W��p�jY0u�`v ΢&��n^�   p4�IM�W�����F�H$LŤ�i���觞���c�N
�)f<���	B1  ��l?�].��Ryb�  `�r�1�Fs��&���p�N���     ؆!��R�H��<�2d���<.O��p%bYS��� �
�2::*   ��߇GFF�.�I1Ō8���O�R���{���|�J��
��p8\��:��(��{�
�,X�@   ��Z��uO^'_��-�!  0��y]B1���Ȑ�8*     �}�!�`8��C(��H��p|� ǏP   �,�LJ������3��q��$3>*c&�������1־L3��f2c_k�z  ����;������   �1��x>�L��Ȑ��     `��F8�d���`���.0����Π��T(   p*3�"N"�1Y�P����I��s�c�VXN�.����D"�$D�   ~]�V�o<���%�%N @��U�NV�Z ���w��~�'�?�_߽�(�8}��w��O`,bY      �aH(����y̞Ƅ��;K`8bYS�P�\�b   �d���ڗ� ���P($�\N�2��|}yj�82�C1�dR`���Q)�͏q;m�Ⱦ�xfD��X�   �sp�\zϥ�y�f �>�O�%�\2����}M�z�)И�D���چ�}�� �T��O���6     �>	�p �x;�!���u{fGm}����P   �lhhH�2͘�n�x<�5��u;c����PL:���b0�yR��X��"&f�{��755�CeŢ�)���6  X�zo���ur�}�H��   �8����!�	py\�+���     `j!�`�&O�����	��}�� ��z��R��*R ��!   '־L�M�W����۫u�j��9:��`(��9�R����h=� s�1�=T�����ږW*�$��Jss�   �m��N��=��-;�  �YJU"	:�|�yL�W<s���      �aL(�Ұ�\c�Z"�r�KFO`��� ���*���c	8�   8��А�e:u��nf�Q"��������d2I(�D�b������L~���r����QԾ�P  0���ݳ�����l1+   f*��" ޥL@���9�A�y>      �aH(&]���.�b0���4��Res�tlW�b �"   '���z���ï@�jD�x��PL:���*���B1���ڗs`�L1#R��=�f�   3��!��s�l���&  `i�xj�
0aw`��p��     �CB1�2�t�'01_�3G^k�� ��"8�   8U6��b��u�jҺ���1#R0<<,8���VS��L&����Y~�_�m�SC1D� ��*�*i��Mқ���] �Y���=(7>x���ny������,�]~\��   �$c<�h�(cB�� ��     ؇!�j�z4yK����"̺7X�P֔"8�����+�rY    '1c2w<'R�ݘ�?>f?'���<Vx��11c�d�6�
����3<gH�f�}�>�>B1�qR�/��^ٽ{�,��{j��e�  p��ՒƮ�O`�x��K�	�{�Ck���      �`H(&Y�
��7/`�Nh�?�q�P͒��>�� �
���y   p3&s;-�p�?��G1UG�H$L]~*��'�L�}�]dߣ�2  `g����^6l� �bQ   �J��l83d�KW0���v�]��z�L���b�;     ��2=U�	����;Z%�^ 0ѧ��ق� �   8���#��8���C]����e�c*����.82�C1V�8����qq3�=1"eژ  Σ�S�{ｲ{�n  �:B1�k�]=O����a_�S��9�%0T�1�      �bH(&W)H�Z����)�o�|���u��78�_p��p�2�, �*j�&   �4fL�v�d}%�j�(j����knn��o��S����\δ���Զ�I���8�1>Lm߼^���em��f�R($ L%����7�ˎ?`$D}���eÆR*�x ���*K�!$��B1�����pi�}      �bX�%U�I��E`�fo�Sc7�Cg0�L`8j�SK*�\�b   �D*"�[<�R������4c7�D"!����,[�b�q)&8�g�H��Z*X�N��/ש��]Q����A��U1���.�����&����n���z��e����iӦ��|5/�]   �[�X�Q_��n�F�cHZ> 0\�ȶ     �N�ŔF	�h�7_(�bp����v�-!0\��LB1���  ��Q֝ʌ����cS	�B1*����$�2#X�n�1Q�$��a�^��__f�b��B1  `����۶m���~��� ���w'pr������VU]���{ $��5��uT�GQpA�g��ܙ�;�2	$( ��@e�fS�%l!���tWU�յ��4����T��T�߷?��,Os��9�O��w T�47t�غľF`L�y�Pq"Y      5�b��̓ݚ�8F��1u	&F�S�����"����S ��   x��s}o���@ �hԻ�o�1�j�L��^��i�q^*��U/�lī������+�2�=  �\���G}T�7o  @���:OGLn�|�¹M�/h���YpzlR}kL��M��     @�X(��$gLihm>�y�o��\���c'8b� w�.��b�}�   �kl,��b�^��H$�F���xm�̈́bƎ+8+������بp8,��q�Jq���{  ��*
Z�l��.]�|>/  �j���<���T��JO	؎x��Ű�bKZ�.�X�     PK*�a"�!P�B�����.`;&4�+T\��Wg��B�Za.4�m�b   �56q{}��	�8���{8���@�H���X߄b�T���|�񸼄s��l��� ��a>3>��ڼ�{X ���5��i�4�]��v�
����"Y      ��b�&��3���"��8�y��5�����#6v�X� �G$^8iP   ^`c7�����7w^71�o��I&�V�'cG&c?ĝH$�%�������㟍��   �~��.˖-�ҥK��  ��+q���ч؁�u�	���     P[*�a"�1�������/=
�J\��������.�e��C 0��p8���A   ^`c����n���8�sG6�ut\j&�C�XL�`P�\����b�p�v��{�s��l�c&Pf���
  0�sb{{�:::  Pk�C}���>*kR����/�7�'�?�T�_9��yGN�o�*�?�>�     �vT�j@�	�i�ă����Y��?�W&ֵ|Fp��Y�D(�Q__O(   �a�!Nk&V2,pz�y��O�.l�����s˖-V�O�����K3k"N���Ǆ������cc��Z���  `G
���-[��K�:�y  �i�S��0Z�,3�?�����O�+�#�6�*o� k{      jM�B1=�~��� ��qu��E(��+�6��0Ep�&B1eE(�QW�gI   x��P����c#c�̎�K&��B16�^��f500`���T����\��q�=�1�Ѩ����0ߜ{�  �1����� ���k��{���~���P�̍	�8cZc�)�azØ�Gp3T     ��S�P����K3��	�73:�ж�6�Q��H��R��8�$: ��   x��K��0����D��1mD���͠A&���N��6�	�؈V��H�י�ӡ�=  `{
���-[��K��O @�{��� �m� s%N��86��E����zJ�_|��y'L�om��k�     jNEC1��6�qHK8|���o��^!�/�5�����U����)� B1   �
�X�韅}>�b���.�;>��8C5���f����W}}����bll�1�s��:�6�=  `[�g���vutt  �KV����)f>�5����ӓ��غ�0W��q     �=A��W�����$8grc�E"�����ysf5M#8"W�km�P>�b �b   �6oG�Qy����6��(�LZ߄K�8�����F��ay��s��c�q�  �
-[�LK�.U>�  �׼��5�N: 6�s�=7t�W�<oιsB��&+8�c     pHQmbq�C��M��Կ|%J��/:y��>y��>�\����~�_pƚ�-ñ�� �   x����,�����f���;���%	��g2�C��)n�x�h����;ہP  x��\�裏���C   ^��o���/_���G��������?�;�q�4*�n1�c���,      �n	���V(�Bs�+��8)�jB�ea�驂�������cS�
�y�w�P^�b �b   �]]]���L(f��h�y�	��	�����;�ېJ���q�2{lls�1��>��  �*�ղe˴t�R���  x[>��]W��1�a��D(%3��/�q��t�     ���pPPeU�k�;�J�)j�qpb�Ig_9���o�w��4�?�%Li�I+{	c�� �   x���ijjR0T.�st\�O�8Q�>�1!!%#���!��n���̹g���`�s���  ����裏���C   x���P�sfE'�~���>������Y�.���}�&��5�     �1>B1N
*W����`&�j�&8#j��'~Pz���fŧ|Fpԛ}L��� F(R ஆ   �y6B1,�����tvv::��׼%	k��T*%8�P��z{{500����x��������<�9�r� �[
���-[�%K�?  �;��ݨcZf�0�a��\VzJ(�æԏ���p�J�q     N)*+8&X�2ϛ��b�v@|�g�l;��m�y3y��}��'׏��$: TN$Q__�   �Ze��a� �B(ƽZZZ��oX��/�d2��O�bl����wĄ��Ѩ��s�2e�  �7�s{{��l�" �N:Ip�c�7N �7tށ��3��蔣~t�CO	����wP|��Qo�r�     ��h��TAY*7�=g��K�'�y����sOikk�w~[pTz�O��,)'��
�����	�   ���8B.�s|\��ƶ�i�66�F�b�c��n���K�E�*s��X,&���oNg8�  ��BA˖-Ӓ%K���W������o�r���B���ԍ���t_�sf���8���l�:     ��'RV�&����y�&�>�̅s������3:G?w�Q�5�z��\���nuuu   j���`���^�ZZZ���J�g�X�����F0$�*`��̹g��Վ�ɹ ����٩�����  ��m�R�P��C��si�>��N=���|T��/^}��ǧ�en��~�ya     �����c����� k��(��S,H��I�±��`�G��+x��7έ;�n�E��^I;{!7 x�   �:��
���؈C���*��*ۗH$��m^���AE"��2����jD=�~��.��e��C( ��U(�l�2-Y�d�9   v�ī�Q�N���4#:���i�g�l�xC����rz��y'     pLQ=�c�j�Vedf|�`x=�FG&��ut�>������ߛ���kB�k����IV,X�bj�P^�R���  @�c��}�����3Fؾd2)��gm�(�N���U��T*e�[��q�s�}6��  j�9Ƿ��k˖-  ��y)��P�ŧM������Y$Լ���cS'�{���     '��!8&�6�t��K�+v[NS"&㼦@�ojc�/JOj��/;i�-{}\p�P!��z��E(���  @�3���X����M��Y�G(fǂ�����p��B1ΰ����׎��{쳱=��߯��z ��W(�l�2-Y�d�9   v��"
6�@����ߟ�6������P�J�q���W����     ��M���v�����([sXr�Ͻ�g^���5k�Q��A�`E�e������ x7B1   �u&�4뿗	���yGǵj�F&�c3���d2��O����������XLx��}�|�0a�  @u3����vm��uv   {��(��00�
Κ���0g\���焚5gl��)��q3T     `���{�۳�檁�*5�����
����6�����3������Y��w��i�1K���*��� x7B1   �u6b!�x\x������tww;:��HP5J&�Z���<�g�a;{)c�=6�`M�	�0�bs�q��0�;�  P�:;;u�]w�P(   {Ƅ����~�ɂ�m���[�����,j��W�z�1�f��`�9��c     �c|�N'z;�Y�A��!��Y�Y�I��L�{ڸ��KO?&Ԕ�,8=vĨ����a�K��B���n�b   P�������^
"���&�b�ɄblI�qD*���-x*bb#Pfp�y�`0���F���8:.�  �_GG�  �2z9��P�%�:��Uz:Q�9�'&����V��5�     �y�b�v(�����*B1�2����?�c7~��_	5c�����G���b����@(����~��ae�Y   ���܆x<.������XC���qC��2���o�S�E���s�ys�q:ù     �^H��3''�q@|�o\�����+��P��X��E�ǧ��1�6      Gd��x�z+�+m�
��_ڵ�It�"���5�����ы/hw��ST�W�>��j��P��W3��ʏP���D�   �&�Z�m#��v6�Iww�������}6C1n�ԺB��x(c[�1�q�ihhP0�˜{֮]��6BA jSSC���Tk����](RSS��v&���$  ��e�75T�)���-'��w~z~��7|��'�����'s|�~�	֘c��c     ���b��֌vA���@/�W�??��@D�crCk��񏔞!T��/�7����k��	{�t�& �3̅�,�  @-��X�|�61F���H���R)�!�j`s���i�������э��
����N��H$���)��P{���UWW�Z���^&6Z�￝��F  T�@>�ҫth����@�oN�޿ɴ%Z�-�nbU�����uoc����0�v��     pؐ�	�y+�ӛ�(W��O��::9K����>�_��#�_p��/T��ms����x"���ZҵB��C ��/v  �7�X�m#�Rl,�7L,�P̎���	y���:>v���,�+�1�EL8�����b�L�\N� w�     x��q ��f4��m���X��QB՚\�،Ʊ1�*n�
     ,ȩYkǼu`Q+�@�y����X���tҘ/X�m���#T�&�}|Vt�(��L�_�{�U
� �P   j������(ngk�����	y��&����"T�B1^:.
+ۼ�s�6��.f�ݜ{Z[[     ����¹�>(�utb֑-��\p����s�5�/sS[�:B1     ���jSNp�[���V*P���e����ߑ�f�1p�Ќ�����*��k>z��-�)��Ү* 8�P   j�֭[�����ņC�Nlm��ȄZ֮�s��T*E(���8���[�|��q���~��=s�!`Ouv�_��5]YB�p��|�6l��  P)��:�y�[�#ޙ+t����=�}Wg�х��J��.���F���.s,3�4      ��)8�P��[�REg�ߞt������M�o����B��������w��g����/f��t��$�dp?B1   �E�\N�L��q�	�lS P4u<ZA(fd�����2�enؾ^��tu�Y�ιg�l�{�{ �ÿ���I�jU��-O����   �k���tƸ���QOn=������7]���}���r�b��	�qsg     `EQ+G�������J���5B1.�w��D*ۻt����j_^p�}�Mu��`���,�Z!TF�P �5B1   �Ef���Xj,�̈́��V؊6T��A'/qC(����4[�B1����Р��>G���     �~&�@(��h�����5�i�|��͂k�s��GG�z�%
�`�W      �qػ'�ސ��';_�'&#��aɽg�ˏ����~���W���|౭�?5�Wx�g���=Be�X ���   ��Z�� ®2!�իW;:��� ���,�H2��6v*�*���x<.��!�}f�8���     �͞�~]�����;Lm��_Ⱦ4�p���sѮ��pn�A�I/Onhm\��̱     �q>�)8�ݡG*=/gVk�`J�#޹���k������{��ˋO\��<n�q�f?=�.\㱎 p����Y4IL
   ���"m�o��X��Аzzz�F���qCȤ��޾f��K�E�����l�9��_���1m�      �l�0���^��Q�0;:iT�PX�x���tN����/8=rX��WfE'�\��̱     �qEgZ%x�;��^��n���';_�ߌ?Zp�G������;>)��YW͛v\r�����(�����P9D  l�Y�UWW���~   ���"m�P�,�ǶيE�}�P̎566�\80��u�iB1c�M(ɦ���B�i��8�؈pU��������s     �;̍	Ÿ���)�r��W�l;s��m���u��"<'���A�iW�f�     ���Bb���	��̩A���9e�A�_x�{���$��s����-��L�Ū�y!��:��r� �B1   �5[�nu|L�P��&O�,�X"�І�PL�HL>���=���Kl�b���w��s�yߥR)k�=      �Z��5�����qp���!ߪU����Ӌ�e�ޢ3�m:�)�ʁ��Db\�??�%]+     `�*]���wB1�,��ո�J�瞵�<��������?����w���+�^x��'$|b\]",��c[��-&   ���Y�c����}�%�I+����>�r9�A��2�Qn/M�'�u���͜{v�湇�     ིŜ��zU'�(��~�)c�>ߊ�N���[�;7����<::��}��F�󇭯*[     �/�{��+կok���]�A�Ţ�xQ��x��>Ǎ������s��Z�u�umw�	�9wѼ���r��p�.T(�d��Be�s l�   ���oww��� |���|>���[�r=�H�P�-�t����*��	/mkb���}��c���M�&      ��c[^$�R�c�[��UMN>�Ƌ�^}���f1z����S�K=��z,     `�����(jY��f�P�{�i�kf��s�;��X#T���|�Ni=�@�Op��S+Օ�*�P��!  �Zb��|��q�	��P0Tcc�zz��"32�bj�ٮ�5���D"!l������%      �ߒ���'ׯ�`��>��65����������o������>pBr����%+���\��     ��'
����M(�;1�k�뵾���sa�[���l
�/\�����*��?��sG����/ �W;�u ��P   j�����87��� �N6C-&���d2��Om�A����P$��pt\�=      ۖ+��d�+:m̡�;���C���sOdQ���	s��������3l�F�.�d��*�     `E�P��ŘZOљ��Ţ�ߴT�L=Up�	�-uw���"W,8�����+�6όO~���^{	�֟��-/	�W( �B(   ����l���Fk׮ut�����@ ?��X"��6��&�(�N����WN#R�^�ܳq�FG�$     �}�oz�P�˙pɇ�����>�غ�Ƿ��S�(���6��ė�9!���~�_p��6.     �%�Z�������998����?�)')��U��N{ط��t�+NY|A���ӭQ�.���#�g�fb<��oyA��A��LH ���   �%]]]V�%�s��f�7n��}�hT�`P����z�!hR�R����}>��"&6�=�pX������P     �{��^�U��5�q��^f���Q��iZ;���ܛ�����=v���f�F�m?*z���̱��     X�+/8�+�NkU��'���3[�똖ق�O�'g9�tG|A�g~t�}w
���{�=���[��l$�ý�� `{�   ���X�m���ي�}�P̎�y�D"����Ƕ4�U�L����
yg��ƹ�@����N�lV���|6      ؎�6-�W��.�߾��c&ԍz)�(�ݫο�߄�v�5����~/n�N�U��ұ
     ���+������C�����"�[�>2��;��5�r�z��^ܶ8+���r\sb�/���"T������g�  v�E���   �[WW��c�����v�V���>Q��ɤ�P��I-2��t:m�{�R�dppP}}}���L(fDl�{�      l�C���s����/(�_<��?c�a��zC�+7�v�W���]�kN��wx�}�%�ޟ�'V�l1�G6?/      �~/X���뢞�O�q�XڵB��5:��"�փ>����;q�i_��k��Lء�ms���K�xܨ}?S�0{^e�ݸDp�Y  �SWW���   ��V(;gk��֭[��ki���N�RBy�h����"&�bT̈́bF��9ڜ{&N�(      �_&ׯ�oyEs[��	���g���V7/j������{a��_��;69�_Z�Q�HU���9�#�      �??�[�?��דrp�~��u���t֔���2���~|}��o�x���O���GV	���E��!�闚�%T�laH�t,�A$���  @-��������Xdl-ַq�6�D�ʸoGM�A��.�L&c�[��q�V��H����9�      ��o7.!S��&�����F���՟��>,�����}�&�t�ؔqBU�o�R     X������￢�I/*#skLǮܼ�s���s�����t��Y�f��������;#]_���A_��q��'�v`l*�b�b�oyY=�~��b �	�    ���b�fB1#����0q�����$�I+�y+.�}T>�t��� B1���{fDlE�8�      ���7���S�[��|��Y��M�ѨgVv~��X#蜅�&M�kY|x��G���պ�N=�^)      ���y��^�
�����>��7�%���/i�(���*���:�O�^�3G]��}Ն��-�ʃ�^x�����^H��L�W����^  �   �Z�b}�3���P��f�r9��)P��J�x��B1�c�L�����ʸ�gF���~8T��:��5B1      ;f"�w���.��a�:��e��WM�>��������`�Y��=���aɽ>5p��*��uOq�N     `�OO�l���B�E�9�1�\�{B15`T8<e�!�]�z��k?�����_��#��SO��8f�!��$S��zC+z7�� v�P   j����^
"�)��֯_��f^���[�F���D'������cg2�|��I$�
"e�g�=��i�3	���/}�|>՚���B�p3_�+��k��ͼ? �n��>7�$łB���G|ǌ���t���1��Z7�:=�Rp�U�M��xhb�)���@L(��zp�     `UQO
�l�f��C��N~#�{��ԛ: >U�~�뒑��ܮl�3�k��`��Z�L?�ӿ0�~l���)��>��k�k9?9�P��	�B   �����ֶ2���3���������ةTJ(ۡ�/y)�e�����♑2�"�C1===�f�
���]u^�yj.���k�ktK�p���;���kr��.�L   N,�7�է'�(T?J��z���B���~ܺl���o�p���S����N�T7j������õW{�0sL�g     `�]�?�l;Ӥg���ҳ�N~3w�{�PL�I������1TȽq�O&�}�o�U�7vy[[[U��眅�&��7�i�''7��5���jI�
�Y�b ��   Ԃ��.������F����
���7�Q2����6�5��gSS�g�r����mB<&ȃ��.2�1c�      ����O��U�j�	����#4�9��H�����U�}__������L�\8�i���;�G��t�Dn�Z{�
9�z��     ��^��m�V�����`��g��f�޺\k��hR=wL�5!PƦN,=.ݜ������o�l��ݷXU����5���	u���':q|��/{jٝ�$Zb���   �n�V�/��bñ���P��}�%	+�f2�|l�bl��mH�RV�^m�W���H�     ����#�����j���5�ql���l&����n�����wt4,Xܶ8�*pfۙ��־���'�0+:aV4�@���=��yu�     �*����Q��T|�K_w���.��B�i�G��}���fW�m|�c ��w��ڛ���-�ҢS�jD/I��WӸ�u��P��f3�]���� ؙ`�P   �[6�U__�����qa�lm/�X;g+>ab(ۡ/mE���)"e      �v����1����Q�L`��^������־K���o�v�f����[���J��YW͛��]4:���^M�f�C�1��u��X     `ِ��`��W�f���*��9:i������)'�9�(Ծ1��p�a��s�C�r�>���^L�ޛ
�n��+�op����է�4�m2?n|Cr��H2"xί�?��BN  �	�B   ��Y�m#��b�]�b}wkii�2��I-g�d+8d��cK,F�H�j�E�$Uk��D"%����ۙl�K�^E  �^��:�L�r��G�}&�2'1c���o��os��=���o�y8����o<����������|�%=eL8�ϔ��&��6��<]:�c     �eO�*qQ�e��\�]�%�gG�A��}B_�v��-�@H�4Mh)=N,���b�y��7�y ��=��zfh६�����OO�t��mmm����+�6��c���a����x�ဖpt⸺D�!PG���ҹ>ݽ�i�� T�@     ���Z�O(f����?L��I�����#܍t�l>zzz����ٴ����q�V��s�.!R���5�)���444p;sc�h���;3Pp�gt  �m�ٚG	�x�	�Lk�TzZ�S���3~qXa�`wWg6�F&���`n���г���37�Ӿ[^Ͼqn]�7|D�:<6�5MiN$�MTa<���g��     ��
�w�W}���l(Ƹg�3��c�{���,�i��Kjǿ�׆F�t���!ߛ�/d��������|������B�;P�������Hc0j
Գ���?k�T_nP��P��	�   ������f7ntt�\.�L&�X,&l�	Ř�c���x&�ǅ=�J�l�zm�@lE��Ucc��ܗ98�P     �Ƚ�Y��������x^s��_z������o���bA���Bo~`�??8П��T��|���3O�l��}�|��@��>�k�GB�P���L��t�س�g�      �+�q���b~���M,��k�Wg�!`[B��ᦀy������jc��P�����`� ;c��X   �����q���l3�C1��G�����l#��t:���Lp�6/ELlE�x��3�e�Ygg���ci>�W       v�U���L��}+�~~�_�P�����<�(�3�K޲�     ��J]��v������z��lo9췛��S�Uk��Q θ}�c����FF��?L��Ĉ�������[��/�o�}i�   T�������®����>2u�Taǒɤ�P�������rx��x�ƹ�DG�Ѩ�k̹��PL�P~O��*      v���Mzr�+:nԾ '<���^�u�      ��s����;�;|�E��g9l���mk�E3>" ���ٌ~��YyY����ޏ[�̢۲٬�l�R���ܙ���C7�|��ϟ/`g��'��Y�a5�)��ټy�6��̙3]���,4ړṖz?���m����ڵ<�\   @�lݺ��1���XL�5�B16��jd�+W�t|\B1��d�����4����s�����N9殼&�HX�Ą�      ��-kѱ�f�'�� TV����5�     p�p(.��`���|(�x`�s:s�qWg�H �qۚ�4X��� ��	��!����"����Wye!   j���ڈLx)�PN�b��VL!�J	{��v������1�K۸�l���~2c�     `dV�n֣/jn��Jj�xA+{7	     �������
;_p�^��z��l_9,W�׏/��o ��y�[�mZ*��H��D4n�8=����� �����>��n����#'N�ׄB!   �Ȅ
����X��\���kii�2n&��������]]]V��ܳ{lm7[�	     @5�e�#:~�~
��{�/ ��/t���	     �|���#��lQ�(�pm��M�G����	�J��h���6��'�M��O���[KN   ��� ����H$���b�������ia��ގ��8�T[�&�2     �]���S�lxF� ������     ��b�dd���n/�pm��X����{u�_d�>��{%�F�myI�ϫ� �.�GX   �ml-�nnnv]CC��ᰲ٬�����_�����%����8=��J��=c�Sf��K�=��־I�     `�ܲ�w�@끊� �ԓ��OW�     �%��+ł|�*��������ӡ����j=������ �\L���K��%x �T(   P�X�_}̂�����5�ʄ	��3���F���8:n&���"l���6�-�H�+l@��)�h4�@ �|>���ñ     `י�í���g|H PN?Y��ҹ>     �BQ�
�2�P��ӏK��1�[y��H�T���` ����?jy�: �K08�   ���X���Ȏ�P��W�윉}8�1!:��b��I�R��O�l�{��)'j1�m��rCCC���USS�      �k�����{��6� �����tl     p����Ip����ꧥ��ҳFY�1�ҝ�~�OO:Q �����ɪ��0�l `$�]�  �j����y)�Pn����}�ڴ��h͚5���N�	����lz;��������m�F��c#c���     �]W(�Õ���� �õ�cJ�tl     p���J�\e䡘K����E��9���5����kt�����JǓ�ٌ��b �T(   Pm�Ͻ���V��J�lm;B1#�H$����0��'lo?�G��jf�6�H���g3R6i�$     `����=��U��G �'�����v�     �ku��:�v%���"�bC�����}>% �]�:u��?�B(�Hye1   jKOO�������Q�pX�=��ۊ;T�d2ie�T*%�t:mu|[�klE����+�f(      ��7��!�
���	���s����     �"k�F�
��k3ї��Xϗ�$K~ױL'���(��&FrՊ�5T�	�B(�HqGj   T#[�����X��n�B1�C'�.M(�1��S�DB�}���D�      �����m��秜, �?]ծ����     ��Z���:��,��^̢�ˢE�ߣ���T�N� v�}��ӟ��܇P��
�B   ����ׄb������ӣ��!~��	B1�����R��Vt*�	���>J�     `��b��:�e_�h' �+{7�uO
     �E
2��Ү�b��EC�^�Y�,�<��ͫ�W��. ����x��;�0R���   l����KA�Jhjj�$��9:��'���Vkk��}���Ï��~G�M��#����"&�"e�����)#     ���ł������/��� F�X�ZP:v�ܜ     �ʽ�B�W��U���K��&�~��)?j?��, ���ߣ����F  �   T[��m-6�>�oxvvv:>��g�윉!��&����g�{�R@�ֹ�P̞11#�߯B����900���:     `�-�Y7|��'&# �;��^�d�     �U|�\p�]�>]������|W�_�[W|��>ر����'��,���S6 �D(   PmX�_�l�b�s�dR�ׯwt�L&3<�eBB�5oo;��r\4Q��mh�ܳGL$��b���ی9v�X     `��d��:�e���y'\`�l�֭�'      �Y���.���^.�J}[w��3eћ���x���� �ӛЂ�ܭH(���Z�   �n���2���`�$v.�&32&�|>���^555	�&�JY��}�r\4�s�^�ƕdb;6B1��C(     `��t������N �=f�k�V>+      W)������*۷^\��㧫�5'��f6M l����ά�;�bd�� ��@@   @5P����Bs�[��V\����&xB(f�e2v�i�k� ���Tcc����9[�"e      峴{�~��Y}h���m1�s�      p�7�������W�Y}K�˧�eQ�������U���?$ x�Ƿ��G6?/ @�`�   ���EבHDuuu��bV�e����
���T�t:mu|/ųlŦ�	���2     ��p�����4M�% x��}�~��     p��T�r����*[��P�n(�x{��� ��c0��+~-�_�X ����S P>�   PX�_����q���U(���������T+�����b�������     ��`aH���X�:WA_@ `r�t��#      \�K}�Ap�=�4�ne�R��~�����tT�,@�����w�'�/��Y� �"
�  @�`�~u���|��j�:�X4U8V6�ut�4��ݒ�d������"e^�ƕdk;��o      j��=��U�S�	 ��J�sl      p���"���g��6tq��b��V�R?�^�d8* �v��G�,�R ��p�   TB1�̈́H�� 6b�f��uܹD"�M�69:&���c{�y��Ĺ���ڎ�TJ�\N����
      ��?k�Ԝ�tp�t�Ro��u�     �u+�+����W�]�;t��Xzv�,K���w���%��' ޴<�N?[�P=�Ţ `W�X   դ���ʸ�x\�sf���b����־SmZZZŘ�v��P��
y��o�q�28���َ����ܹ���q v��k1����������M>��7 ��Q,}}��;u�!�+l o�����w      \���u��x�J�c�����W�t�\`i�
ݱ�I}j�q�=f��^��rE�����G(��
�B   ��֭[�����,���K؈.��w����G&�v����ݼ11��|���Wb<�f~755YyϘH� #��'����㾉Dn�D<��k�0(  �j�9��^���m֧�!*�A����w�c��      Wڢ�U����G�ҳ��7����5�՜��;�����ІbeՆP�]�Ż$  �:�r9ka��`k[���عd2����tzxN���G�m����+�E���8瞲1�7�!��     T�S���kӧ'�( ��5��魯
     ����T���(V��b���r�B��K��?����4����^q���٭� �}�`9?�   �cB��f�9��ֶd���$	��4���>566
#�JٽCf4��|���T}}���P&��f���%R��&M����ڭ��hI������<E�8����   x�ͫ�^M�uxbo���_�OW�     ��6*�EBU)��W�A]��J�N��s}��MW�%��!�m��nJ�N6�$�:�B|�  @u����|fnhh��f(�̛�|>a��ɤ�q3���]�N���o�^a+2E���lD����N��555iΜ9������?J�F��N:d�>��	   ��ͭy_}놨����p���n]����!     ��O��6�	U�ܷN�V��L���޳A?|�^]��G�vm�������� �*   �6�)[��l6���>b$;a^�`0�\.�踩TJcǎFƄul�ݰ�V��PLy�ڞ�� ���ת!D���V����e�e�����5�B^   ��'ׯ�x�6]yЗᆨ@��s����J��
     ���ԵB�)o(�
-�ź����r��n\��M����w�' �-��,�c ��,    ���k�������1E2����NG�M������^��O6؊�yi;!�Y�|v1qw�s v��`���z��i  ���ѻQ�_���a�O	@m�z��z�g�      \˧o�*
U��+ls�N���7�gv�^܆E��F�Z�ol� �s���ݥ���f^K ��w�  @u`�~m�F���m�a���&Mv�����PL&�F�v(�K-"e��V�,���l�j      �䑎e�'6Qw� Ԗ���Al��      \�a]����T�P�|m�ź���?��bNm/�LW�eM�k��pӪ��hǋB�+
�]��c,   P	�B1,�/�@ 0�����U�d2����TJ9���Vt�i����ss�=�e���H�      g���{��똖�P��Z��W�/      ˩�o
U�2+l��\�]z��\"��ӿ�x����/+j��v����� �Mf�&   �vfa��0����lS��X;g#bc�f�L���^9.ڌK5s�)+Jnhh��8��GS�L      *�X������e��Y�IP�^�Y����*��&     p���J� T�ʄbڔ���?�gw�E6l��{�v]����W�?@�-�Z�+~-�wCP�B��    �3��\.ge�x<.��	��^���qmF�I2�t|LB1#g� m�b|>�b�����1�sO�����P���ޝ��Q�����t�}�!	9!܇ x���/tWD��*�?wQ�x�G�@ �,����E.E��k�oP��}O��L�Ꞟ����WOc4H��1]OU��W�t�g议ꩩ�SD�      ܕ)du������U��d��;���ܠt>#      P�~ �Z�j)�u�.�έ��!K7h�������*��_6o�OV�Ny*��P��a��   x��I�L��"�bv�o3��|>om�����K���F����Ɨ	�l޼��q��      �o ;��,�^��5Vs��ܨ�����k     �ӊ�H?Q��k�=+6�s�+έy�c��hJ]�>3�T���LR�]z��ri�r��7��    ��5�ڼ_6Q�/3Y��UMM��s��1qx7�5e�Y�R)��!�HX����[��X,&�?[�.�      ;:Fzt��蒣>�HU0��@%������j�p�      <�5�����O�^�u���\󛍏*m�'�U �/�K��%�i��	  o�D"   �n``�ʸ---�`Ɨ��Y�&M�$�	$�u?��:��� ��ݐL&������}Ɵ�ǕP     �=/'�k����7=SU�*�B���+o��5     𸌳|^sT|����Z����s�y����T[�D�}k �3��E�\Ge�B�y�g ����+�   ��lM�nmmƟ��Y�Ō����J(f�ĉ®��ɦ EL��T[�k:�V*�"�     `�#=/+
��C�Y!qq ���9�?[�G=��      |�ǚ��BE(��[��l}NE=�܋�Ć�+W�AuUQ�<��L!��/�Q+�6��P��a�   x����A
"��<��P�ʱ���al&�v�ZW�L$��l�b�1�d2�2v+��������1S�L      �닪��˳�/ ���������     �,WF�	���c���wn}KS(4o�m�G�����;rż~��f��X/T.B1 �FUUUi)
   �*�[����Q]]����>6���cB1nK&���l?NA�.�����D����k�=�b      �s˳j���gf�* �r�t��'     �U��R�B�p'c�g��s�Py��Q�h�o��#�֛c��}&�tي����+��F(��2�4͕�   /V:��26����Lط�1���F(fppP["��:~�B1��)+�h4���:�R)��&R     �����j�}l�?�7ܶ�)�v�c     ���~���x[a��,TJ�l�����ǘX̏�߬�)�<C �1���+o��K��G(�ފD"�b   �Y6'W�b1�<LaӦM��K(f��X�mP��fP'
���YA`s�C(�|�ck#þ     �;�{��G���o ����^w�      |!�ejҷ���^(Ƙ�E�@?pn�P��gt�+��{G~\'�, �3Ѧ�V��HL������    ��9����E([!#����4����R���M�dR��PLSS�����u�-��=�񭯯���{�l����6�C      x��Zs���i�=�d��MO�W�     �O���Oh�F������M�DI���)��BV�_r�.<��:��pO���OVܢ���	 ��e�   ����j�0Q����	���q���;�D����j��D|�k�TJ�\����O6�������P��=6�w      ر�:R����f�[ ���M��W��      _�H�P�ܟ];G}C�V^/9���A�b^?^~��?�u���
@����`�o�||�,n^�@e1    ��5����Y�pX(��	�N��y���d2��i���
;f;�����=A���`��5�Ry"�     �-&V��g���G�p�9�������O	     �G�W�
�Ι}�k�.��[�ȣ�ł���R4���@�������t�CB1 ��_  �eL֯L6߁�al&
�~�zW�41B1;788hu���A�P��X��)/[��9vo�=&L      ��[�U��׹����� �Rt����;uO�"     �Ȁ���� T,{�����k��sV�Oˣ
ł~��e
Y�1��0��a]��:��"� {��  ��lE=��_^6���C~cB1nK$�v��tl��N���K������o7��o      �tw�s-du�!���P� �/s��y+o��=�     �3��m*��ٵ_v���hy�	�皻�9կ/����8ڒ�w�\�M�^�>S�OT% ~�D����T�*���q�    �*��jxx���6C&A�FU__����Ƕ򛶶6�ǴB���A��e�h3&��-D�      �3n}I�̰.:�c������g���ӟV
     �g�;n*��P�<����
��s�ӗ����i�e����T4d������F�Yz��Y;���zy���7���e��=�wL� �V8ޫﶆ۔�f   ��L���3ok���V���0Y���$ėw�v(&(�E�1�V�=eUWW���Z��i��H     ��-���/�R?8�P�p6PN}�������"      _)�I��B �/���*��O)�;�{U��{��wtPs�<[-��;O�.��+oU����P( �Vu����   ���z0Y��ZZZ������f��	�B!a����]�v��l�t��żf���'(��M�1��!R     �놻����.�bf5N����y-}o��:�E     ��lQAg�j1y? �1�v���������<nYr����5��Q�Ҕ:�O8��-��5�8/w;W� T�H$"   ��L��&뗟�O.�S2�Tss��s555�����Ȉkc��;g��ijjR8V�
z���<�(/�����v}\��i      �g�2I�~��ׅ�}Ton;T ����5����j$7*      �1q����"�7B1F��hH'����㶤�u�K��{G~\G7�����|����?	��\ �Vu�w��   ۳5Y?
�q��P�a�-B1ckkks5�HpU�]����b1��}��������=�����     �C*�ќe7�˳ޯ�Oz� ����ו���\1/      ����	!P�3�v�
:O�R�LEb�<n07�o��k��A��{&�  ;7�ѥ+n)�ց���/�rEp   �����]`3300��3g
�fB1�6mrm���Aa���2�����2�YM�Æe�������ؓ�}      �L�X(/�m)c�C�c�y��zÃ�ݦ�     �S����Jo�X�~]�8��t�6y\���OWߡW���Yg(Z��Z=�E?\�u�휤o#`_D"��  �7���L�v��(���ߘP����P�Ѩ�Z�d����XLA044�l6kel�=�)�y     🻻�ӆ�]t�G�m����$���7k�`�      |�1e��@�V(Ƙ�����I��ܫ�<����u�G|\k9Q����/��w*S�s�: ��UW{�,   P(488hel&q��fx�V��o���u��~�	�ek{�MP��6#R6�YAbs]���Ӂ(      �ϒ�:�ūt��ӑ���U����S�n�     `,WD���ɛ�k��q���(��8�B���[t�KW�ۇ��7��d�BN?_s���^$`W�Ţ `o��a   ^�Ǖ�筌�d}w��Ԩ��V�t���m� ��ḞP̎��e�h3"�J��6�e"e      �֗I��/�J��q�>:�$Aww�s���sE;��     �*�]*N�
0o�b��Y��P����`vD�Yr��eƻu�
��q���t\?Z�[��0B1 �E$   �5L��Xwuu�>.��wO[[��c��x���%(�E��V�=�hhhP4U&�q}l"e      ��/�����#գsg���*λB��]��=��      |,��>��Z-�wC1��P� �֗��@�/�ߧE�՚}��m��.����P.%  ʭ���oe  L6'S����0���PL*�*-uuu�Ι�BMM�FGG]3�H��L&��mb�A�.�	�>����>.�2     ���@��Z1�I�<�,�0Y@P�Ln�e+�ͩ>     �X�Y>�yzZ<�ϮM�+j���{�#/����/�\��!���p�l$7Z
$�����=Q( {����4�X,
   �
���c����a3a�P�����͘����z6:MMM
��
[!s\�<�p��P���6      S��ꋿ�ǧ�K��~�B��R�s��zV׬�O�b^      ��W5O�	�B1W+��t��t�s�d�H";�9�n�i�ӿ�Ն�*͊�Ra�3ŉ��s� ���je�Y   ^as2��@w��p�®�����I&����贵�)(l�{���[��L&���a544      �!_,膎����z}��3�_�Y@��M�����z     �^Hj�~&�/��1*������׹�N���/j��&}밳4�q��J`~It��'u݆�(�c����"��   x��x�PWW�h�P�[l�b������b1WǳD�2��KP�Y�tZ�T���n�΂�v��P     @�y)�N_\�3�{�:y�1*��Ku��;���9~     0�j�~"`;���4�o���!�t�|fc�W_[|�>1�d}d�;T�
���[�p�Z��(  l�����Y   T>D���Vƶ9y<�l(lň����������Z&�j+`be����om�V�=���x��l�ԩ     @�Χu�[�h`��������N�_fGt�ڻ�P�b     T���|�/���kf�eJ�\�GQ=��;R>�-�t��H��:���&N����yݶ�)]��pi}���< �*&�   �R&��26���e{�>��v(�QL%���:~P��6�Q6�YAD�      �t����U:��������7��.����Q��      *įդ���b�+գ��ңνY������K�轓N(L�Gx����t���0� L�  ��0Y?8����F������{��&����.��P�;lƣZ����H      �-��ܕ��.�z�3�������?�ޥ���	     ��ܬ}^�� `��1j���w:���ν��CE���]�����{�:��`^4Z��ƎG���O�Pd_ ��j��  @eb�~��8OO��Q�d2�\.��Cchjj*=F�r���2�M��bʮ�}��]߮mC(      X�ܿR���C��~�>2��
U	�3㞮E�f�}J�G     P1��I���nQ^�N��L���l����9���Ou�t�+�鴉��s3ޭ�h� �x�w�~���f�^���X,
 �U8   ���f����cn#c���um	�΅B!�b1W�#�a�I$��6�ss��������^�Ǽ�����m�g      ��\h�W��׳}+��?�Y�x�ʡ���5wiEr�      *JH�P���9*���b�yڪ���u�s����_��KK���N;Iѐ���ۚ�.]��n��X/�\� �HD   �W���[�P��l>�bvO[[����x<.���p���%.kk߳-Zw�
�)��(�
      ��$١�t��c����X�Q�-���n�xX�v?�B��R     ����<}���l���5��*��z������;M>��gJ.��~^��q�N��Xn̍覎Gu�g9x��#`<TW���,   *��P���g�1�����	Ÿ�fŋ����c��� ��Y[�8.c��H�ĉ     ��):��(�Ǧ��H��\1�����_oxP#�Q     T��.�}K�n��#��4���A�u��"x�|�g4��+o-c�x�{5�a��r�v����i8��B1 �CP�   ��F�����e{�>��v(fppP��ᜠĳ���6��Af�q7�s�      ۶��>���eƻu�~G	(�g�W誵wkK�ߏ    ��d:ͳ����������!��y1|Q`qb��}�*�{����'k�N���2{�G{_�����t� 7�0�r5   �bttT�T���Lַ��d}�-��:���J$���v�涠�}�D�      ���~�x��zc�,}fƩ:�i���t�C�nx�4�     �BeT��@7�C�5�v�r��/�-�I�H!�\�X�}�����/�'�Q��v��k���k�����5C[���PL6���͛����:Ngg�.\��}�s���1Ƈy�<��#��{���}��cmذAӧOWs�w�{D"   ^�d��!�}mmm��G(�o̱���k�e�h3��1M;l>��{      ��̹�f1���q�m�"`_���M��K     P�҇5_�����f�����t^�9�jUrż��zN���B)��駨-�$`O�_�����2�Y ^���W�6m*{$�0���zH��u�9��SN012��+V�2���V�ZU�Xg�1�pX^S]]�og  �?�b������3I.�s}�D"Q:�
���^V�a~�u�X�a�(f}�gU)�LZEe�Ⱦ'x��     ����|a�?jV�d{j��V����[�ًQ     ��u������	�K�{��ݢ�Y!����Ob[0桞�:c�[��)�PK�A�X�W��kyr� /��/q:;;�e���5�f,X��K��_�"��S˗/��C+W'7�@���4k�,����K��  @0X���Ep����Ǿ�����M���b5�ZUUU�9r+n`�w�c=�XLAg�O�������������� ��l�o      ������?�w�>9�M���S�QF��ꆍb     @`�I9}PW�[�>��������PXw9�TI�3�e�����k���蔓4�~����?�_��l|T˓�x�W~�c�����[���ޫ��}�;�QSS���=��S�7o��٬��!��hŊ:��=5(�   ��?W�2Y�����f�>������\}}�@J�PL)�c��8�������ǎm�w<w}l�}3���      �s��/��Wt\�A��ަ��&��-Iv���O�ɾe*     �xE����I�ш�}T١�Z���&U�&���0�BNt���_�[�Շx���:K�T>�����n�������0�;�������f�ҥ�袋t�%����Q��j�*-X��j$f�B���kזb1^��V]]�og  �&�a����؛���3�	Ÿ�f �K��������9�j����v�}��P�96h�9���      �'�y!����0Y�<�D�<��CUBp��"��iyr�      ��\ͺPsD1�"3k� ޫ����"�Ĺ]qG����������5��][���;��P.% ���۫��.yɺu�t���?�����`���)�����
3	ɬ�f�Uss��oG\�   ^���gmlB1��|�mƉ����p����%`bb<�\����e4창�!     �=�zx�殼U�u<��Oz��?��j�
�a.��p�bݺ�ImN���*     ��
�Ӛ�;��`�b^U�<]���y1]�ܯ���L?}��u����^c"7��D��ֽ݋�L�
�y~`b6e�YmڴI^�|�r]y���7�!���s+W�y��]�VGq�jjj�~/�HD   �mf���(Buu����;l4������b1WǳH�����s[ln��{��P�Y�f͚%      `ot��������M���L8V�t�j�$T�5C[tO�"=�u���i     �K*��Z���Y�B1�Z�?��z��͹w�*�9�~]�C���a�z��7�Mz{������$���uw�s�Js�`�K�P��-h�ƍ��Vz���u�����O���'��s�='�2��9���
��}�p�4���   ��m�'mii���<�l��잶�6W��>6#n��{��<�^e����\�      P9�riݹ���rH�:m�q:u±j���o$7�Gz_փ[_Ғ�     �դ��(���b��Z�/���/�٪pE���5��=ڤ�x|i�\��&_,�O+uϖ��\|�
E����̕��pB��W_�c�9Fp�,�\N��կ�u###���Ԕ)S�~����f�   l��`��]6�&���q30�H$���7���477����)     �x[5�YZ�]���5��g�	:�i��?K;to�"=ֻD�|F      �RQh��K@3c�\C��O�|ݮ�~��D5�/��o6>ZZf4쯓ڏҩ�G4��L�gir��Y�G{_�@fH��ٺ��6����L&�k��V^x�,O?���n�*?0��	&(�Z��   �6��B1v555)+�ϻ>���h)�Y__/����<On�KL�8�̱��!{Ǳ��]d�\D�      P�R����ZTZ��iՉ�G�	G騦�wu����W�p�bmN�	      ��(��5_��YpC1�,�-�@RQ�;/�� ����:�!�贉���G�=�$���8L����Ae��1��l^�xO�`�ҥKu�G
�q�w�/�빳�S3gδ�=�I   �M�����f��]�PH����&Λu�P�����];d)&dBAeb9�B����X0��6�=Ay����w����qv�ޙq��      @�l���ΧKˤژ��vx�<��&�m�Øs�7�z      ����Q����p�j��ڠ�t�fh��2���f�Pgi�j�=:�e�Nl?\o��)u�;2��'��O�+�d�R�e��,*��P̶��䦛nҏ~�#!Lte�����<y�jjj��O(   �ي�---�]&�ck0�N�:U�5�X�n�+c��N&�䈓�H��W45#�Ͼ'�L�ʬ�6^k�lV���jll      �����_�13���;�;Jo��C��($��n(Z1�YX�'z��B1      ���
�s�����Y��ܢ���2��c*�z��,P���8���\�{J��[g��rB�����3�RmI�������j��P^�DB~�x�buuuiҤIB�[�h���L�����P   l3�m	r��+l>6�=?ikksu<B1�B1&`b"�.�J)�N[�P�}fc�f�=�b      `����Z߱U7t<���z�z`������h0"�nId�K@5�?ݷ\�!     �u���>�+EY�cV�ߛ��u��QH�w���W*���]0����+-��j�<C'��1-35�a�¡*a�ų�Z:ء��k�h`U)��Jؐ��522"�1��C=���>[�|�?�������32W�v�   �d~f�����o%c��`�� �w�ۡ*�6m���f�9(���>kc��Ԩ��N�+�������&3}�t      6�F�x��r��t��;Doh�����6v_*����F��X���Wi�H��s}     |�\��ۚ��X¬�Y����[��~��~��>AP��+N�b�TEtp�:�yzi9�Y��99x{&c�0K7hI�C#=4d/344�����O>I(& �-[&?�d2�SCC��c�  �M�����rV���jj�ꈶٌ�،E��ۡ�]�d2iml���(e����lml"e      ��gersi�ɹ_�Ҵ��tT�9�}��v�����^&�UC�ZR:ϽC+���+�     �1�t�F�o�R=,bV��Ջ���)�X�;��3�=l��}5��,����l�_G4O׬�I�퉚Y��µ�t�]���ֺ�n�Jn���FfG�;���j�ƍ��Mcc�P���x����Wf��1�c   [��x[L$&
	v���X������P��P���%bbs��J(�l>6�? �M5Mj��w~�{�յj�oS��e   `G
ł6o--ww=W�ڤ�X風��K�D�"��٬/����9�]Z3�U
�l�      {d��|I�t�  3�92��B��U�j�.a�L,�Jq�����Kᘃ&iz݄����pT~S,՟��T�֏lպ��Rf�s;����)
V�M�R�+��Y�b�N8��r� ��ي�D"   ��u�b1�>�σ	vf2E��;��&�����[?�&	��PNP"&6�=6�X���"e �����Շ�������>���^����   `�����!��ׯ�DJ�X�8�H�\צ��:�����t���w��0k��4��§      ���&�TH��<ٙ@	� ��ݵ@+��'k��PQW8�vKw:^Z��_񚯷F4�6�I���X�|�i-��߹�\]��H���t��ȣ�l� y&���x��{�}���Z���}c�'6��S~�f�B1n�֭�;�P���--   ���w�n&�{CSS�B����f��ĉ�]kkks-388� ��	J(��'(����|`s�      �S";��kJ��µ��N�i-]uR]�纛���R
������s������o��ʏ
      ��a��5��bì�=5O�yz@a}EE]�|�I�+��piY�ܴӿ�\]��H]�sK�ܮ/���T[QuU��i��-��HUu��E��P.]��90n0�H~T�bQ�|��I�K�KK.��_���5q*��w�)���Vhe��z������   ؞�t��d}o0?��X��8���cB17nte� �b�q���!k�e�hs�C����`+Rf�a��i���
      �D����w����ה�mo�4�.����hU�_���{U��ҹ��a�g�*8��_�.�����|�s2��y�۟�n�}     �k֨�ok�n�Q�b��B�����<ݠ*�Ĺ�Ig		�n�t�{D��' �W�BA~�L&����PL>�/MN1�T�T]�[Z   ����oml&�{G,�����	Ÿ��1ǡ���4�؆���y����U�٬�����>s<�����1c5�4i�      ��J�GKKW�^�      �nX!�S�.��x�j��Bmv>~Z��ҋ^z�  c�q�S�P�nttT~gb1n�["��    [�����*x�y.6l�`el�렟��1ǾL�#ђ��H$��m� �y�k���U�H�w����1c)#            �B�+�]�*}Ws�%�Ō�z��x�f�4u�s�� ��I~�(RSS#T�Jx�C���c��   �I�RJ����	�x��p������b1W�d(�f�8(�D�q(s���^���oڴ����{             T��B����-�J>¬��4O8(c
���0/ �g��a�Y'Mcc���Dbl�����  ����Yۼ���D�������vW�3�� J$��J(�f��<�6"��1�=             �W��r���;������rx5�&���ď��o ��X,Z��1���&���=c�*mC$   `��I��g�0�Dϰ9Y?�+�ϳ>�������R)W�j(&�LZ�PL��b1�;ZZZ��ms=            �}����M���|�PL�5O�ݥ!�߹�-�k'
 �f(�����d�}5y�d��M�6M~VSSce\[�   ��$i����z6��B�P��p�y�ŔW"��6vPB16#e��͂w�\�m��             ���
�v�5O�'�Y��6G��J�:���Ug9�Y��+�@2��l�����v�aBe�9s�"���٬�����ʸ�0o�   `��I�A	"��	ńB!k�\-"3���6uvv�}�.� �3�<��������v�f���}���|>L*��p            �eI�ߊh�.S��
��{n��E��O��Xy}Ź����j �HCC���|�S�N*��Xab1�V��ي1����L   ����DA���\b��d���f]�5k��kn�n��|��ӣ�!S^f�2�[Z	�x���ٲm]loo             xL�B���u�.��+�eD(Ɔ�Z�|���ՏT�Ϫ�/8� �͐C]]�jjj4::*�y�ޠ��*���-o�e(ƄZ������KW1   �40`����͂��	��B16�E?ikksm�L&���Z���q�q� l��81�U4-��GFF��o"e�b             xD�YRHרQ�k�2*���������r�Np>������� T(���\9���K~s�i�	�p�I'��o�ߘ	�����Z�  �۲٬������d}�1�ɦM���m&�cln�bL�!���T*ee\�	Bd�v�����}��P             X֥�~����\��b�b�9����m��)��9�r�  ��L�[(Ɯ�����0e�r�!Z�j����Ճ#��FGG   ��LַC%�=6����p3c+�b����M:l�9L����I�����26�             ���^g����G�W�G���2g�^QZ��Q
�,�q����
`s�QWWW:y>�H�/�������]v��y智��K�555֯(�k   n�9Y?
Y�׳�����s1�v���Q�hT�L��c5f��c�#A�g����m��I��>   {+����gv�5���������~�5����g����Ƈ9�k_��&�;mڴ�ޯ��Rmm���^CC��f�����g.hd�5       \SPQO+�[T��5W]��^�PK��f��]4���� >e;cL�4�7�3�C��,'�x�f̘�6�8� ���   �m6'G��חNB��؜���fK�L;g~v5�Swww��"㮠ĳ�e2Ծ
J��ol��6�G   �Oے6E�_T�ºx��;���TJ������9�dG�
��~�6s,"Dts����>��r�Y��X���8�W�l�%;{��}d�0��}m�cG��R���秿������h,��#      �R�t��t�.W� �T�o�oј�5[oSQtn��Y�u~��7��{3i�Ll������	�s��g?�Y]|���:�~ڜ�M5�   ���������b�IB1ckkks%�N�4�x��cA��،�����$�����<�^  �;���z�^��W���ÿo�
��a�Kl�RB=n����}���՞0gA�v��V	       *HZE=�*ݣ�n�e���aF��5OO;���m���*�]
������Lm ���ӧ+�L*��˫=�P�~��B0��Mo�)����~X^eN2�%/�,D(   n�9Y��F��툂Y'�M�&�[�3��f8��Wj�v�f�,(1�����r��1���f            �>X�,���T�{u���K̨��y��|����q�ϤNTH�9�w:_{��4 <�愑�+O��S�ׯ��+��[�"~p�s�/^���>yє)S������V   �6���mI�c�hT����2��x������6ֶXLPd�Ykca�8<<��+I���}�'����C�b             �-��Bz\ݫZ) {���d�r�����Hg)��:\Uz�s�*�]�s� ��]A���]�TJ���򒪪*�w�y�0a�lMMM��w�[���iy���2q�Dy�   �������mO
�Ι��V(�f��O�Ř�GMM���g��KB��v*�	�c�1���֎��rƌ            �]X+���P���PK��ޚp�3j+�-�;��e�����t�Bz�����g�c��@@@M�2E�������3��+_����0f͚���?_�^zii2���Wt���P   �d"1�|���---�7�禳���ض#~�f(&����SP<��V�5�)�1�Jg�5ξǻL�������D�             l'�,��������T�E���`\1�6hj���,���k�T�r:FEg	�h�pLH3��& S+ 'Ţ��P��X�v��X��^���/��SO��������7��y��&�����T�ט��K�   �M�'E�	��X,fm�~B1���.�ϐn�|m�0?G��1�`�u�&��qs(H�ߘ횭P�             �̉C��z�F&
Sp�a-���
@�1��eJ8����Z_�dU��1:���)�W�sn��|n/�~�s� `^��b1����=��������[��V;�w�C��K�J��|���O��H�A(   n�=)�L�7�|nFFF�N�U[K�{W�ϴ�y��+��)���$���V�J<�f����Y�pX�&"e             �I�Y�	�=
�>���|~5c�u�8�_m ���ص�j���,O���}Y��S��SAag�o֭m��lp�u>W9_gP�"U���O��;^�f�Ќ3���X
�
�ƞ6m�.��BM�:U��w�q��+4w�\�Z�ʵq��ì�&L�W�I(&V�jr4�  �8��c�,��csRt]]!�����4i��kmmm��bL�'Hl�m�ϲ��iH�ǯl>?�b��ЦC�|�_ ��������AC��������W�OG
 0�jj�H�Z*       ؑ�rz5 c�J������R
;�S�ӕ _ ���s�K��e� R���+T�#�����Рe˖�=�Dt�Yg�#�H�6�;&O���/�\�^z�+�+FO�>]555�=	ż�o/\��  0�n��!plN�J��l�̺I(fl&� �b�q4[��րDL��;����;[��t)eBv���������W��w��"�}T�M�-��TX}�� @Y���zO����        �P �5�&��)se�P(T�1L�Ƅ>L��S&�b�-�6u�TM�8Q~�'�   `_1Y;��P��V(&�˕*UUU�t�l��ح�d2[�5 1���bV�7��              �f� \�P��������z��b   �&��ۓ��k555� m:��2��u�O�|�XL4U�K�R���v�v�P���z Rv�              ���  ��P.�b   ����!e2k�2Y���s���eel�1	�hoowm,
B(�lm��jnnV���b��muuu�팭�'D�              p3j �!�\�   �-�'C!��w---�B1L��-&z
�\9V�J���2�yl�sY�lG��v�f�k[�n�2v?�2              \ŌZ �k� (sq   ��'C����6��Q"�P.�#�9�3�	_���e*'NT����2nP��6#P&�C(��l�b��             �.� ��P�r���*M����   ʉP�b�92�^L,���]ص��6WB1A	(��X�HP��6�=���ħ|�f���{#              ��3;  P̤%B1   (7�чh4���z��lN�7̄}B1c��b��344� ���I(��loӰ{l��ɤr�A!              \�{  ט�Z@���a   ��d}��v���:�'mmm��322� �d2V�m@(�Dq����[��;�ϓ9�oBz&L              (?B1  ��PN�HD   @�ٌp0Y�b�����d}�ͭP���*�	����V<�z\�}�?�~-��G�b              p�   T��j��  ��FGG522bm|&��C]]��Ѩ2����mƌ�ĭPL:�V��f��ƶfr���SK b<���k�}              �a6- �6�z �   �ܘ���e����+c�^O�bB�PُY��~.���Ym��ᰚ��U�l8���C}}�"���p�              �S�g& <�P�r�&  �2c�>vW,��1�aL;g�
���J&�ektt��fu�1��	�zξ�üL��������b              pO垙 �B� ?���Q>�/�����/J�YW˥��J~RM(   e�d}�.3Yߖ\.W
w��v���͕����`�g�J���ieܠlm8lnϰg�k�V(��{$              ��ٴ  ��GQ����G-`_�y��k�  @�1Y��v��L�'36�ٰaC��I$�<y�*U<�2nk@B16uuu�F��?�|�`��bQ�PH              ���M p�9I ʉP   ���d}�~���Q��Q5�9s��k&���aU2[�AŘc�6#e�XL����|>_�b�$�             �M̦ ��P�r#  �r�9Y���Y�PH���mF��ĭ��Ȉ*�9�g��/�d2�\.gm�V��b�5a�=�3              ��i  P� ��k��c��Ď���?���ۄ@s1�k'ΏK���t(��DT�?Z�R�*jz��q�����J�;��rIU��Q@>(��,���@�c��C�������L�;���@�=3��x���3�̰_�3�<3�|�@#�A�K�.���������fԨ�4+����:U�ĔJ�T��f��ӥ}ꆟq'ɵ@�lǎ         h,Ӵ 4E��� �$ @#�HL��m뷗����g�JC�q�v111єuC�J��[�ZiG��{�Kڏ׬H         4�iZ �B(h4�  )��F7:I�$Ձ��/����P̆���������u�bꯧ�'����N��k9������X��Q,SYƹ         ��4- M!4�P  �4cX���>i�bVVV��A��&&&¹s�����z�҉�[RY7��b�����Φ�~�9�>�D��zϒ��         �E��W�  t����   �277��������v�'��\[|���;2�����ʺ�.	��)�
Ŵ�)K�y���         ��P MQ*�@#���  h��/��~�������[�l	\]�Ph�:��YXXHe�n9&��SZĦ�P�Ǚ����ndd$          �#@S��� �H���� �8i�g2�ԣ#\��Ci>g�I�B1�����F�I+���P���JX^^Nm�\N���Z��#         �e� ��  @���i�э����K���333�kkV(��Q_�|>t��"<W�b�R��=[�n         @㘦���@@����$I  ����|X__Om�l6h?i�7j'�
�P_�p\L�5��iK9�         �xB1 4�P�,}}}  �mff&��s������X���	�b1���~޶�������VWW�#�χN��k8+R֖�~�f�{         ��b h8��Yz{�� ��fggS]_(�=%I���S{���χ��5A�(
�����L1���{���dB�TJe}�         h<��  t�8,  ���гa����b1�;776m��:�����f�!�N��Í�������4��         @�	� �pq0	����  �[�C�1�@{J;���B1�C1��\�LҊL]��Ӿ�c�V(fqq1�������          4�P '4Ko���  �_����E�Di��~|>h�pL\__����2<<hO�5r�̙�֏瞷���         h�� 4�P�,B1  4B���$I���x�=�����	\[�P��\�b�y'�ߩ�xR<�Оr-p��        ��1I@�	� �" @�-//W/i�>���=��f䨝Ŵ�l6:]ڑ�\�x:Yι         :�	 N(h�  ԛa}nFڏ_���v1>>^�<���h}�|>t��_����di?~3�=         �P&ih8��Y�b  �����T���okccc!I��~7277W];�xs���#�����/����=9����)        ��f� ��! @��=�3���zzz���x�t�R*����ڞG�V(�b�@|M� S�s��f��\����CG         ��L��pW��� �!��2�L���ۯ�' @���f��0�PL�ÞGז����J �ӥڈ?g�ו�ҫ������Ce��         ԟIZ �j�������� j�� �P  ������G����3gR[?�bv����B�h}�pL��KM3.�{�^����)�J���*         4�IZ  :�P  �#i��޴��ôcG�"��Z_7Lb`c}}=��c�wtt4���k��ٳ���=B1         �&ih��Wp�!�bs  ��8������!+���[�;j�֗�PL�q�x�I�$��r-p�ٹsg          �O(��*�J�Yb(fmm-  @=�a�4C���á��?����O;:�.�������b�u� �vܩ~�� ��         K(��Js��>}}}B1  ԍa}�!�ͦ�~���v��d����Wk���ӥ�H��E}d�{         �c	�  �1�_ �z���Ku�B�hqX?~V)������������P���kNܠ�e� b���gbb"���~�~        @'��=��S�7��\.�f���� ��I�3�;��@���S�m�N�>�ڿ!�b�b�-��ZW.����N��C=��Y.�K-ز��         ��0I�M۳g�?�l��v�F�a�h�84�$I  �zMm����p��:�{����B1�3���@��&&&�+��v�g�4�=�6m
[�l	t�;�3|�{�Ke��>         h� n�׾��-I����|�4���t3=���[\  �c�Ν�a�Xl����sO	t�ݻw��{.�?��ko޼9�-��ZW.��`׮]�?�a*k:t(�v�{�7<���aaa��k�z�         hS� ܔ���?-��qJ��o��Z��8���� j��P�P  �244�����6u��۷���?�9�g��}�c�_�B���6f˖-�ֵm۶�b(&F6N�>��u����w�+�9�O<���/������#{         @c����MMM}�\.�j��V(&���7� �U<���ᥗ^
�Νk�z1�я~�:dMg��r��ѣ��_�rx��W������>��066
�B���	��P��w"G�	_����ڳgO��>�<1�Ce�<�LXYYiʚ�
         hS� ܐo}�[ٕ��?������7�  ꩿ�?|���X���['�T�����{O��n����O�cǎ�S�N5l��طo_�Ї>�>1���|'�Z�򖷄�[��n#���'�W��p��ņ�300P=��߿?йv��>��O��~����ٳ['F�z�p���          4�� n�����l�\��ҥK�I���������������˕����os�L& j$IR�p���?�������R�~�̙Ϯ���/^�_^ݼy���]�o�PX
  p����ѣG���?������ٺ}��y������j��7::�x���/�g�}6�>}���ݷ��m��Î;�/3�㲼�h>�`5��M6m�>��O��~��azz����x^۽{w�����$:_�}�?����s�=Ν;W��_��s�С�y��          4�P �mjj������~�ӟ>�裏n8� �(�c�L͗�sss~�ǎ  �	qz�޽aϞ=���E��/~��_����I����^����Q��[��]�vU��>�|�;��������<���K��ŋaqq1Fx7�=2�L��4>>����W�ߖ-[7.�F�9�y智|�q1�/�(��b�)��N�:U=�\�p!,,,�˗/o�{V��1s�-��m۶��;wV�7�%����;��W^y%���1�\���2=����T�=�\.l߾=�v�mհ         ��+P ���O?��>_���'|���@��.��ͽ�u�$��رc��c�  p��u����C�P���^h�y�{�=��~������G���n����z��!�����         @{����ʦv���f{{{K��600�7�/_~}z*I�?y������_   p������·���@:b���ѣ��?           ��P 655���������~��d~�T*�@����|���r��ym�����?�l�e   ����B.����7���b�yv��y��          x� 6��ɓ�Q��we_�$����w��� �*��b��t{���?������ϧ���9r���   �w�qGرcG��X��O~�����y������]�v          �7	� �!�������[��P(�MeS�0��R hI��b�jtt�,--�T�O��n�T.�yzzz����>   6dxx8<��ᡇ��b^x�p��Yј:)
��[ow�ygu          �9� ��رc�(�˟���������=5_�@�����
�\�/^|����y���ue��   ����P8p�@�R,���\�+W/���������/          ��� pU�r99~���U�������+۞��	� -!I��CR�}}}}����n���3���;|���   pzzz���D�          �,B1 \����'�$9T�ott��L&so�R�$��r�\�g�{&&&VΟ?�Q�k�*�����z��ş|             �-� �����R*��}�$IGGGw��_���9 ��r��*Ǫ��ձ�u���###�-..�]s�{��}���|              �6 ��*�J��l�����t�$��e������T h�c҉���{+W�*��q����������qm��t�ĉ�<�ȹ               -N(�����㏖��߫����{f``��׾\���O����� �b&''�zzz�@�$_���Uvm�f�5;;�`��Ƌ���+��              Z�P ��ĉW�	����+������J�҇����� Т&''���ɓ�;>>��r������}}}����n��ۣSSS�w�ȑ�              ��	� ����U6[k���L&��r��+�#���g@�;x��J�\~bzz��$I�o����W^y��7��sǏ���Çg              �(� ������͓���$Y�f�o�\����{�� �D�V�l��я~�ROO��^YY����-�r����              �(� ^w�ĉ�R����r9S�?��=[�wjaa�<xp= ��}��}qzz�T6�����qm����?~��_>|��              Z�P �+����yO�L&s~pppjrr�@��˾����}vii��ܔ���?��7��;��              �� j�8I��߰����C�ݻ��'O�|�r��/o�muu5W��     ��rE          B1 ��ȑ#_ ]�������y&  �$�  @�)�J�        �T�    �J�D(  �6�         @*�b    ��+            4�P    ܸb            �&�   �T.��b            h
�    �q�            �@(    nP�"            @�                 �8�                �'                ��b                 Z�P                @��                hqB1                 -N(                ��	�                 �8�                �'                ��b                 Z�P                @��                hqB1                 -N(                ��	�                 �8�                �'                �����3��>    IEND�B`�PK
     8p�[����  �  /   images/b53b2c7c-bb6b-4047-8ddd-b279832d777a.png�PNG

   IHDR   d   B   �s   	pHYs  �  ���R/   �eXIfII*            (           V       ^   1 
   f   i�    p       �     �     ezgif.com  �       �    �  �    �      �w��  �iTXtXML:com.adobe.xmp     <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="XMP Core 6.0.0">
   <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#">
      <rdf:Description rdf:about=""
            xmlns:tiff="http://ns.adobe.com/tiff/1.0/"
            xmlns:xmp="http://ns.adobe.com/xap/1.0/">
         <tiff:Orientation>1</tiff:Orientation>
         <xmp:CreatorTool>ezgif.com</xmp:CreatorTool>
      </rdf:Description>
   </rdf:RDF>
</x:xmpmeta>
�[n  IDATx��]	�U���{�����F7�Ѐ���*h���$I�$��8T��c�ʤ�d�d��JU&��*Sٜ$f☩%JD�
���4Mw����}_�s޻�nO׭��������g������oy1|����߹���hT�.>����v#iK"�f���!�#���8/�`�9-���UaK�q�aN�aIZv�`��)m�rP�U�9��:a��\v�'�w]!74CQge!�,b�\A7���]w#mM!mNɻI{Yc�0��<�c�,
��a��G��u
�!OIsRڲ�|!.�,D:���}��n����:~�_T�w}�i�O�<�8U�<�ن��۾��˞W��.2���p j`�ۋ�� #����]7�F�9]���n����b��jőA?�m8T3z����`6�7@���5�1���L#�a4�*O�0��|w%B���8Z<��"�OQ�##a$�,�{�	�r�c�8�8*���p�ì��-�� +�#Tv[	G�	wc�~|�u6�_	�ǰ��J�W����{g�)Mt����CX2�6�9��g��4$T���;��;��� Ӯ��Q�U�$1N&��O�c*,�
��13�f��b�F=�^,;M�py��[�٤��r�
M����R�Rw�`	Y`�6"�5��J���E�6��z����
Q]�".��Q�����8�`6�-�h�z�l��v� pu��Ը�%#��eWT]6���I�P/��c�~=�fŘ�h�<�������ճd3�""߫A��|�z�ë��|/���@$q���ɀl.W*'R�w�IR��S��NJ9N"L@��?ǸO���XL�0R���ap+UU!�	�7�~�7�A��zy�လ����C5��C>�O�K%\�^q�g�d�R�W�p��n0L�HB�*XC�e�i�o�1�Buh9g��~�%�V��f�����Nt��겫a%��)�'��z\FQ����K��\����h����x�?B>���Յ�����\�%�b��PSmCo_v���V��rZ�v�I5E����C1TU؉��p��s����%�PW�T:�?������}Ǎ@(�h4��f��cH&�C#Qd2�z00��
8���=S��XE8�u�݌r�E�q�Y�v�1NH�BX]��-��:y
�Ch�)��:�FR��[#U�D�jcƸm�?v����l3�usF�e��q2����ߡ{0ؠ��`����Tfc�7h�2�,HO���20i�h���<�0��dΩȐc@���S�@=�ޑr� >��
_W���yאe)��1#x1��n�Mǋ��sT��u�ڐ#��B��[��b\����qS����+II��\��?�&�A�{��%�ep!E�nfB�:��ݻ�p:�t:�*s��r��U�2g�B�U8]�}��`~��26�|�T��>�0C����W�n��f;�C>�ZB����,�K#�����hA����p=q�����Hw'�,���e�%cApI ���<y\!t��eDx^���q�#�at�w4�&^V7yS9GqG]�e5��G{Y��l��� -I�1K8���0F�H�~�?���,����Ŗ<A����`NY� /�6���g��`C^nQL�aZĳI<��"z�c33��s�Y+�=fv��arYT�V����"���G���Ov���H�6m��l6��3��'؀_�]$���`���ǉ��F��R9RF���cu�jx^8MN$������*W.&&g0�2�2��~��w��RC�D�r��X�gj�>������K�c�X�]f"���.��o�\��
eG�T��x���k�rw����%�"�3b��n�%k9��Ʉ��r��ԉ�iR�Ia���COOrd�X���4!~04����Kh�^����X�X2&��,0j�N�+�_9_Ž�S�~
���Y�U�a$8�zo=�c�r�����D$U�O|��1�yꤧ��qy��Bv&�B8���D:��g]��^x�^�3q�n��>dHO���kE�������
�'�b:�:��WͿ
ۻ�#j�N�m4100�w�yG~3�-�v;���p饗J�����:U���3��1���R��'��	p�-�-XZ���c�zہ�Hf����BrG��i`È���R1D�Q!�4�t���ف֊Va �J�D���jTQ�G�5���ar�33wU�@�܁XJ�i�{�|��֭�33�I�^�3�TJ�Sq�	��$(�F�.fÖ�[P��Қ��ӻ/xQ\B�نFw#C��uբ?�/�r#���t��v!~�X.��@�"���W,C�x�0��l"3l42�D&1{f�"���N� aJL��gF��b��o>g�gg"��L�h�֒�%����o�i�&<��9|��Ϣ�]���0�8ʬeⷳ$������p�/���1 z(2��+�a溭n!<�5�������%fp;=6V6�D�x���ܹ���.�"�UY�0�9T�bC���Ð ���PSV�M+6�C�����U"ꨨ�G"#bK����?/b��a�j��K	��C���Рq(<$��sl_�^���ƌ�;�U�'f��-�S�t̛7O���>L�b��0����rfB�94~[۷bm�Z,�Z�n_7�D �ԃ�!z�R�����Xd���L��}gO"�}��>�c�R�I�W{,[�L~��bO��ߝ;wb׮]%�rf&"�;�ueuBtڏ���;�{3�������v4�[G�B.�C�*0�6����q�ݻW<)6�2`$�����Du��3��`,<�߼�X�A������g X��� {�6�#xy\�R�6���IT��mVLf��I�`,h	�������R))��a��!��F�>:���Ư{-���uk�e5���m�iarAB����r���<�~�h����&T<�^L�*Y��w6�z]<
_C�,{~0����Dg�S��>�]�pGBGND���=��@����#抦+Ļa���o7"�Ȝ�����h�9P�^M6&�ug'w���N�������-�>�.2�rX�m,2�*op7`�W�A5.]��˰�gϩ�TH x"���@ޜǜ��Z9âAS�*�}֓w@jN�*�tm��L�afn��������!f��?e�(����h<#���9�4s��+�H�ϐ!��C����x�`l�����	����L����g�!�\R���Ig�8��y΂N�+��M[]��B/�p��ڊ�����6�s�=������|��1���G��f��b�N��#���;wZEBlZjZ��(vD���с�a�@veY�2ll�(㐅��b�;�0��i�x�8ĻԶ�WO���*O"-kZ��6���\��Z�@RQg��u��	Cd��hjIXp��p!�[����f����`����3��C��,�c���D��0K`� ��MN�ӅK�"֚)�����NHp������_�fM�f�)�9=�u���XGi?�� +"�7�t��ȒADZ�S�}�7��o�4.?s�aWT�(��?���ق9x��XV�~��er������)��DB�B��õk�ʴ.K͉��u��ˬ��CNX*l^T9�$z�JN�a�p���S]]��(�!֒������p|�9�Ygsn�#�T�1�a줃Y��9[w܎��v�,�gY
jjj���(L���uR����O�����(�/�Bm�[�H[�3~~jJQ��k[����#5y��
�d>]�GWUU�1�L�ϛ�k��Μ�T�-K�T"��uM�pB�Ф{Lt�ۡ'��Y���hmm�ē�rY�X���.�gƪ�;�;�t[WY����Kj�8'<p��믿�����^��h4����YԴ���?� �R�P���s��(��wvj�	ӑ�6g/������԰*[�`�̭�'�N��5 &d�3�~|�RE�z�8׃��4*�k��Zθ�:��A_{?���%#��y�p�9�t8eĞL'U�'��X:x�'�8�w���H�R8-Pp���Z�p��b�M�J��^/L�Vf���"����'��P�j֭�;h�r��N�ө�/r�礄���9�� R�3����+�wC���ց������؍�7�x���,G�B�i�HR�$��A93q������l-\4fd��:^�x���Dw_7~�����M��G� ��b@�H{�s���%R�ϕܯ�:Cv8uHd��6��k���j�*(�nչШ�����<r�#b@9��#���,��TA���»6�qo�^��z����X�-�[���H����.}���bD��"!��Hޱ,E��s�I�K�R��O6�;�d���i���u�oP"7����r�L�����|�|!cD��w��f���5�U_2�}�1����G�rT�����C烺bpU�*D�D��=����6����Z�x5�*���g��[֣�V~J���TX+িH*b�a��k�5]�����b�W�^H��o��-����?�_<���h�"49��q����4�{ٽXQ����i(�,W���<<F�Kz��<�%'|�po������� >������ JK�Kp�^�VX����tUK��dCq1a"p��N!��n\8�BNF���T�j�"R~��'�2�����U�i�|�����<�s�rO]7��9 �3��]����W�%���G^�;cߚ+�%��K��b�yr���~�_�Jl+���a���*yy�Ǯ��u���tY3�����W�BK�emQ,����?������/�><2��e�Y_��ax��>Z�L���X����zdÁ���.�x�+�U�?b�v�`��y�fܵ�.ɗҁ����?~����6�͞f�}�m�84Œ�3�8��u�2A]{��
�>��o��
&V���$1�d �d�(S&o��j5Ye�ˣ�+�D"�8&���~\U�l<0�ph���sj�\	���l�d��pV�]-�B��;���ϣ��(�����P�W��xu�[�o���W%?�cU=���i(�D�tV�s��1Z=�2�Y���ό���ے�󹔜O�r��b8{�Q��������/���0GGFq��<nϴ��^�Ep˂[D��e������薱��,&����Z=/��\���0#&��d͹�)�+��}4^�ۡ:$$#s���S[W{�tV����sެI1�''��h����9� 
�<L���x�^�=n t��$��:C �:��*���cccbG�˺�(C���;�~o�	����e"���eG�˨��*�P��L-����o�k�����$� ���H�Ux�&�͜-ȹP|��esΑ��d���ק�=�;����"!����Aڢ(���*�K�`U�j�����x��^B������!��Hޯ����!�I#K�n�)={O�'*.�g�C�E���{�K�o�'��oO��x.[��7��M�j(�*fo�ĉk%���\[�+����zo��6sc�*��,�ņp[XR��=�N�S�b�z��|�����w���I6���j,�\ ��m���]�n�t`�{#��Ll�!�SbXd9��$�����K/���.�Hz4�N&c�r�G;�ʸr6���
K���_Jrf����K���>�h#6Ԯ,П~�~�O~	�ӻC$���⭡�^IXдi��ɀ�"	��9Yz�^�rO��t-74�f��	�b����WV���α�׿�W��`Z�f]w����6���ͺ�l�";�0��ڄ9zV�+�-��ό�t�[o�����a��h(���t9��#
��"�ب�wE�aZj�u���ɺ��=N�5���j5u��4�z˻�C�s�}��v��Ų��Y\K����/�Iy��'I]}O���<��z���}7|?��?�QB�zŤ�Q����]xz�ӳ
��HL|���\r�H�T2#$%��[�װ(oܸ���B@q7'���4^��F���֪�}��f��7�w����.�t<dP��Jb����-w]�nA7ｨ�FD?n�1�F{A�f)$,�U�*xN$	�����`j8�f��<�ؼ �y �Oe����n��이��L��S��0�����%K�H*%�f��J��ҥKe�H�'��80Umlߵ�=�%Ǟ�sv��ŋe�Fuu��É�ŬVr����r�U�wl�HG��	�ۻ���y�������3��[�T��2�l�� 1���÷͍\:���x�����)�Q�l���Ɲ����{>�0^3�q&���EOJf�74xN�YGʦ���=���'�.�=9��Ib��c˳�:�߇��~�÷IK�3*L���@:
V����K��C�O=�����'����Zn4�������Dy��c�s��l�}~��L XJFͳ���S�,�ng��b�0�a�>�TUWU�*J�ܭ�[Q���϶���Y��E_Cw���bX]�M�cB'��s��� ~ֳ��s���}&*��:�\���j�Z�y�oO�+6��e��y,�l�::�EԈ1������R���l*��țb&�/�f�y�����%�����6�U��R�4f3���[3�&��6ILVF�Zs}�eq��F�G�F�#��t\ֈiYʹ�/��-�VQ�:	�A�o�!b��!��W���~�wdW���ށ��L1���G�xQ��&)r���/�~Q�\��<'�D�t�u���:����uAk����Be�Z����_'�r�K���x�՗�!�����B�1�y��;v�J����3��y��+����}�髷������W��?F�w��]A�y��f����󹛖�/?���8>�i}���x�!���K���Z�8�;��솽���
^d+U8O9mq�"�󖓷/�!���r8�	�\�M~�;o�5�k�;�;�#w/KPt��:�����r.�+΄O��Ϸ��<�R�223x�A�~\q�B >n��Fa@}}=�7�:c�����o>���#��$��ƫ�'�~q������\�kw�1{��4J]���{����mYӂ�5=	���ţgeϖN�U 52��    IEND�B`�PK
     8p�[�ة� � /   images/8f771a2d-db90-4bfd-8b3e-8d66edcda07a.png�PNG

   IHDR   �  w   `�3�   sRGB ���    IDATx^�}xT���{��T���DE,�"��

XP)ҋ��.ދ���k�^D�B�bQA@��zKoSO�����0�7���y9��>{�{�w��῟��@	3��wV�;%����_\�8���Q����O?� �9r���[P);3���qڣ���%�mݢ�!����f�Gnnn���|��펳Z����Yv�=�cǎ�����Q��l��wϙ3����|�^U�ӄԩS3`�Zm�+WFFFrrr�Ç�q���~���o�fV���f<�ࣻ���fK�,��p�¾?�����BzO��yN�uH�EQ��<,�^�@o۶�;]�t����O�,�wD�����:u��g���5j��F����F||<� �n74M��b 9y�$֬Y��3?�(����^0dy�'%R�>|x��S����`�k }����~o���G��5~���Wi��#5����z���Z��xM��U����"Pa�[�v{��4o����p����X,6x�n�]�z�@3���������Ҽ��q̈́	:���K|>�ǒu8�1��e��4M���Oo��$���͛�ְ��iU�&���>n����� a@@�KC��os��8�i��c���x������C�L�4���c�/�w�qǏ�7onZ�H��$IN����ݻ�;w�"���=�c��m���bذ!|�>����C~^!lvt]��a�8�s�<�g�hÖ-���#����8��O���֓V��ׯ_�j֬Y��RB�e�����E������}����|�g����}�-��g� #�4�~?H�(x�l�,�2��!>.���ߩ�y�ũS���ZNڅ�ްaCԝwޙ�q-$�g$?!#��Isйs�W?�䓱�����*۪�a?����C�ݷ�w���2�� &&��DE![�
��w�4(��4	A#��o�y��'NG���Y��ʂ��4y��^��0ܫ���J��� ��n�?����z�(���&L�wԨQ?_��/s�5Ɓ,u�xRS��?@��MS�ωlW�N��H��K����&JQT�\��f��x��^~�^�	��իW�G�������(i�d���Fk�O?�dmٲ%��~�	0�m�|-ǡ�����1P��PT?{9r?�v;��5�Y�W�!�y<X-vH��S'O���׍=�����q	O�5jI�8�[BFgq�_�G]�.��l�	n��_v���<��(QRG��6l�w�]w����u�Z�2�>7,	���@"�dZ����oUNgR�����fs���3�����e_WoժՉ�zn)n�Z�j ���q�8"噄@@�A(V܆Y�vm�{��P)�\�K".1jԬ��e�{n�4i
��A�UU�� [H�+,Aa`sB�)�40B*�|����i�rv�$�M�a�;1|�h=z������R�F.3f̰q��M*~Kq�"R��燤=�~��$$5j׮���={�/��xiD��q��w��8��߿GժU�q���7�X�/i|(M�n�����
�=hذ��g��.P9����������عs���o�7�+���ѣ���Nӧ�D���4}Up"C�� 0B;'�H� B�t���>��#FM��:��,Z��Y�N�~�����ҳ���>��È��8��-�/4iҘ�L#��wd�Z���!�!�Y�7�c,�d�]��6��Ė���Z�Z��?<R��a��U��sy�/1`l۶�r�[ۺ�7�岳!��p�~�v��&�$�V��K���=L�\�&���b��~�?��2Lw�/� �[ψ=h֜�&�9~�o��GNN&����Gr�%F(d�g�Ġ��iԊ�S������no׮��H,�o��fkҤ��������Y�hQ���~��p��7b��޽�7�ȵ~��B9�j���)���(�Bh�L����p9���3]��f�^�����Y�f�ٯ_��ɨ&uY>!���C�N��V$�1`�~{��Ov|�A��]���I#���C_q�A�P��^7ȥ3�᰻0c�l��������#������6m�4RY��s��w��/�D�m�08�E���4���9Z,
}_K�<�1����� D����^�W_}m��u"���?���/���?3���ǉ��]���8�g$%%:y�d�+�S��Gڏ?~�רY��@�$��敮��8��(6B��c�;��O���q��K�n���Z�DJ�hů)��A�UD����k��U�AF�(�0��0p& ���n���.ɦ*�bԭ[�����7$IU$�c�X@��s3Q`lܸ�OH�g�`F o��j��U08��OCӵ� #111-##���H������.kD��s���$��^�;\�(�%C�xԪUO�`Ȳ|6qV$����aG;3�OĀA����xR!`��k��4'|PRQjZB��u�͛6��q�� ��J�YQ��R��C(��o�q�n��]��pqĀA6Fz���G�O��BU�,���Q�Z]}��b��΂p'����<��<.�GO�^��|�@�7��D�l��{%g���Aң�u��_ׯInڴuF�� ��y�ru!��R?��䢟W�\�ܦM�ӥ~�%.��� U����')! ��VWR%l�ѐ�p�s!�J�6v�J��ur��|���ڵ;Sn�A�����<1���awX���آ�///111����Lbs��!F��*f�~6�A�gO�R��dfr��)�|A)ϞEn�M76P���?�!-�	EQUU5"��p�R��K�,I�ر��p�1���������M#�@�Ofv��J����$U��p�٪,������M՟U�^[�LZqJC�Ob��@�.A�qK�����[ظM�6�Ý0ATM��-0>����~��7@Ā���C�x�UfR���e���366��<t�FLBQD"򒔠�UU��(Gt�b0(��Y�F��#Ӈ}/Gd��w��w�;}Z���<60x��t]�˃)	��qݮ]��wDD�J?����@��*��?����@���K+�� ����l6dg�2U2�(m��/y�kT-r7�SR�s�\��H͚�����F�N��1�	���r��>��N�n��� I����<1�i7��3gƏ����A�XHPp��8��g8��7�STT�QEݣ��T@���Sy>ǒ��)q$&U�ȑ��=
zA��C���#:t��}E��Q^���ϬY�����gO��1`��������TQ�YK�w�yk׮Ug������nI�
�T��oѢ�Gg22�����n����'�|jr˖͹|��s�l�H�ጢ��8��^�38M��' F��m�-[6cݺ��{�v���$�R�<����}�W�疄;a!�Q�As����7z�6���I��G��P?۩�Mݵs��l�j�q�$IH��U�=/�����s_?nB������J��0 k8��p�4�j�"UU;�����O�����g�.���0;�x��<����ڥ����p',����
�㭷�j4hР��1����S��jI�+�3{�n��X�tI%�q��F�
{�zv����1�m�'���z���G"ٖ*�o�s ��ahX��c>۶��"w�Ac�Y���i<��S/0�����(�z�:uj�!C��]�Q�q��>��G8�}��4l߾˗-��{K 9����f��N�}���?|�_��'�fø�Z �E�>A��A�k���i�9���';>9x��ԷK��+\Ì�<'��I���z��������x�,0�n�+��&���.T�{o��Y3gM�R�R%��C��<x����_�J/gF "�V):�(<��3���cC�84|�r	���3y��&Æ+���������-_��2�q�T���skv��s��e_}���UwO�>�:Wf\��`#��g���f֊�����g��v��:h�ЩW[)~_.�R''Nl:r���J�����I� 0v�ޗ��˓�Ԋ�E��_�<}���U��^_����2f�k���{��� �w��NZ^v'�v�zdL��ao�;a!�3Ϲ&�7n\�1cƄݰ�cǎ]ǖ/[U�r��f횪m����oV}튣�4�^��x`ەf�0�E��̢ş 5u�1��	J�E>{t�V�=���!#�]�y��}���q�;��رc���=��c۶��Ƹ�($��Æ��vΜ>��ҥ_v��}gi^��� �WK�ʻ���<�n��Ç�~�4���h|��<f̘�ƍ+��z%۶m߳��k�]j��ΝyO�^}�=x`�QQWbb�/]��i��(�"��8�/Y��c>u�K�WB�7��ѿ� 4iz���^~�4������G�~�7�X�{F^�\��رk��e��_r�<'�ӽk�_�.]�c��A=E)u��0n��-�ؒ�:�UBÉ��F��zuԈW"�̬\���� �dĈ�O�0�r�����<Ǵi3�׶]�V,_}kIݰ�*w��2��� Y�}���ƍ����RK�b�aT pp��ѩ�C��(�؝�ӻ�i�ⵡCG���Ͻ�udD�����gqp����O���_����>���AΧ	��" `l�sǟ+���Q}z���zFfF�ys�=u�L�[n�m����7k��di�e���E�>��� ������4����CGF�)WR<�9z��r�С�Ǔ�-0�6��������Z��G���Q�R��^ ]-�d>F	q�H����CL��_~��q��}QڍuI���I����].[��D���~\ӽv��N��qƌ���:&�0j,Z�ɾԡ���e㵾>$5ƌS~�����v���pv�ؽm�ҕ%�����{��*�U�~��ϗ|qw��OP$�L�0l�/؟�:�ʶ��+9?�y-$F�x/��I6v��'ǎ[>$F���aڇ3���]�X�u��f�������=~��EE��:uo^r`������2�~Ptѧ֧tg���������[��_���:��w�dc��m�_+V����4y�i����`��M�9|�U�jի:�g����R�h~�=�K	w�l]Iy�}������[�=�2�a}"��� ���wo]�l�m%�����uú~�Q���pK���i�jպ�2�E��9$u��K��=-Ǧ��;��q�D+/��!`��	M�8������0�������t?����.��ֻصk��W�hc �,]����7�K�wc��_�\s�}��wUD֏>�3r��a6o��1�B�b�Յ�={����2|��s%�`�.�y�n�<yr�aÆ��x>�C;rd?O�������y�`��?��\��D`ԯ��':�?���/��E�uz��#G��q5���'�SG�6��A�'}hQW�=(�v��Ç�5�.~��`�6lX�l�������-VʄӉ &O��CiǶ|�տ�(iAޛ���o�1a�/������K��3kN��K�<��y>��:4uȔ�;����0�8��Z��֭Z?�ਡCGN����S�ޗ���C�����1����<eE�k��c0s�ll�c�����X9�^�݀����6�8�`Z���K�X����Ͽ����0�դ!X���ܹ+�<��!/}'��-o�Bxʔ):�8*a}"*1����H$\�X��w�ï�7;~½X�����~�b��<��EQ�2�߉����)o/�ۧo�Z�R��1}v���ռy3���ʈi���LFe.g,�~��wx|�K/�%^ހq�<M�2���C��)��]x}ĀA�۶m�mv	v�����ǫc'�b��i�$��0���z�s�<�X�_~�ن��@cd�Ra��L�d��:B�u5��e�&��塨��U��� 2p�';>?`��iaOX96>i3L�2�Mjjꪰ�3���'c۶M��i9[�XXX��>��3�|�]%�B��t�&՜R-�E����c�[X���73 ��q����b�@�Ջ��nʞI�c���<���ܩs�^tU�����w�ԩ�<��p�5�����U�Āa&u��y�5d���h�i�2�X3@�=�ݏ�\'{'RT�j�������zj��	p$u��%;;��H�(�y��=�g�v�3`���aOX9�4��&M*_���Wټe�b�d���O{�R���_꜏��z�y�ŗ�R�5�Cq�?�>���лG��)o�$�����6��9s�4�իW�) ���-���Z�k�j�$S�0}�=���c�����f�۳}>_\y�|��W�Q\�}��߸ظ�$�t�ڃ�6I}�ǳ}¦���ƦԸ�(�pUT8�Ƽy���ѣ�ԮR�͛��#0Z�h��y���]��\�н			����5�Ks�c̝;�0���}�[j����i���'Llױcװ?����O���>���&���G5|��g�OQ���0�Cc�?d^+��2�ju�����}�f�=���p%F���w=z���s�� ��%>o޼[�u�=�����ʀ�e=K6��(�� ����Ξ5�y۶���Z�jmIOO?K#(O�������t��5�S��� �-�ܒ�`���>��pwRJJʟ�� �Ǘ���.�ܹso�֭[��|E�ܼ�W>&&��0��'s�����f�c;�IV���ڲ����m����M��������7т�7τ�{���������Z>))"ˉ�,�M���tE�x�+#**��հ|���k�Dغ�~����oߞj�^�-�B�,C�r�-[�Ү]��|���>��/LnӶ�����A�ʕ@�hGQ��o�vg
���~�x�W�o֤�'͚5+����2eJ�S�Nݵ`��������~5ϋ�=�B �!�}��լYs~�V���i����~O$TI�(���U�Vag���`	 ��#"��hP����G�k�%�a�;Шѝ8r8�D��޻o=�⋃�o֬Uɱs�	��h���W;����c1�~��փ�j�<l`�l��_Y���&���#��S�Wj�|��q�>nu6 I�}
q?w�֣_�^��-�4o�|��u����Syb���1gΜF�z���xF�� ���u?H�j�`ioE	��f?o�eUM�5�w���q��j&�DA���r�4���=��9-ݬY�U7n|(t�fy�!p�XB��C�={�m�{��j�$l`p<�_~�ILL� "�P�zz�݅p8,������g���i�H����н{�2s"�5k�͆Z��-n��U�D�zqW�Ч�L��80Hb���wR��1)ap:$�`?��:-Ag���:gSp��������Bآ��`
��Cw�o�����<�SUU���`MT�x��~}���ի�Oe]��͛�Y�~�D	�1%O $Y8�lg^b�GzW�.�/�K�����dw����82{�y���OY�`AXnk��X���*��W��P^�Q.'t��M���0�'��h���5�n.1���ϡ���5�Ŋ��|n/��a9tb#G�R�WDH�x��'�u������\�s_�V�|�����0Lmi�/��T�KN�����4jamv�g�Xb��Bw���i�?����u�,@x�st@�yS�P:.��"�Y	�|���7wV�=�\u}I���E����u��uo@~~>4��d������u<x]�fpP8��P6���<	ɠ��A{�7t��59����P���;#��bpyZF�#�Η�e6̦��:u:գ{ϧz���KY%F�ƍ�n��G��v�MEe�PD:-�j���1���j�v� U���<��¤����S�<��L�С�������`H4�d���t
I�i�f��e.�K��������Pc��82���m��Tp^/$��|����`o�g��N,�$�e� �_:��O�""�*&���!(*�6<
��В�^�	DAVt]����]�&Nh=d���-�    IDAT�2���/ؽgwGQ 8�S5�#IGKK6�G�K��j*D���غ� 5:?����)�������N"~/;���(�=��^�Q����A�<$��L�X,���q��7x��wS>��0��&���*z�&��f�To@����D#!�Hz{��Ӑ��H@���;k�p�:���q��t� ��d�0x��^S��t������n��%��э<Y���~��_����Ӡ�.r��A�:�H��,�TU�+J@�9f亲J��^�f������\�5�U7>| ��!)?lZ�W�,�x�s�Y�r�<�{Հ:��!c"�q�J_}��a���`���'�<u�I��+Ȃ�^�=z�8\�g|��MU5Оӵ�Nٹ����{�����w]�y���-��Z�	K��4�W�/������ۇ32��[�4v`������7���~P�����}w޼Gd�RU���:u\_�'~�paM^Ѻ@Ӣ]V׷�;?vaMY���׮[�.aǾ}�d����W�7���6���/[�]��ӧV �LF���{�>�ǔ��H\��J�y��!\�k��n�˖�h�G��ջr��4֯���6:�x�36|�!i��_��،�{���ۧO��J�]_����g2�À��o��ݻ��*��\K�,��
�
<_CPſ8C�ҩ_��ҾȂ��|޶"'9UE�Q����رc�Tڧ\��~�駺���<� ��Ͽ�W�>�.��zŊvY��|(R%v%��սw�!�~���o�W_�hV�{��E�*�
6��c�^����p�����qQ�D��/�ce��K�A�������Оm��ȯ�>��ҳ_�+�Kײ��������5T�iH��=�u�;��"`,��v�����G��������/9k�
:Tj0{J��v�Z��ٰ�3�>>�}�բ�A3`�5����
����4�7��p�Lv�.�8������MR+�$�J���Q8��Y7l��;aŚ������n%�7�vc�|7sٸ^� ɀ_�^�"�͵ Bc��2vrn��Qg燆K.��6�e��8��q����'�`�P!@�����%�]K�0
 �T��*/��ƥ����״w�Nl����Zx�4}����Ϗ�Ӡ�`AqT�ϯR�(���$�ǥ#��̀̖Yԇ�3x�ӫP�3�=` �a�7�0�z�	�^X�BX9�z>�f�����C���z�r9�x���h��6��dCҼ�9+�h�Ek��T`��pR���b��'��(ˮd�q�� ݏ���,t��j����3X�������D��@��d� �;)��FvV��\P��l�~�9�cpp^��<��x]r4��~<M�Y����ռ͵S�����
̟��ݻw�<0ޝ��-S_�v���P��	������,5���ag�G$`���)�dx��\ �7V�Q�Q �QQ�!���O�YRe(�D�dȺ
Q7�S6��048�3hR;����'9pZ�×;�ڪ��)v��%�GY����jX0�p��Bw �.�~��ڶS��`N��؜��">Am5� :�����,B���e�F5QK8
��^�"ÈÊ�~d���t�5Oof[.�fˀ�~�Z�OKu�{T�+c��/�>�:n��/ME�AV�ΉP8X��#����A�q~��5��`#  ���*�$�����܇�MSPݞ�?V]�ۚ��Ȕ� �S�g��u�C'"�}��lF�&5�,d��灂��B%,�\��&��P٠����%�.J֕u&/q��S� ������Ѭ�7X���g��ia+��
��*��ES ��L2�^Ӡ�}H�q"��A<Ҩ:�[OB���W�ě0{}6|Q)�4v�,��K�ZOL�4�P���v�<��ilx�Eϼ�^y�G�g΋_�Jfު�������D����P��`a�AF5��T
tP8�iӿ(�I�<|>�6z�A�i\��i8�L��|>����@!`���kL�@#U"�eAjZsp{e�����9;��qX���ZL�HꄀA�i!����er+e�$�z����&խ��zq|]�i.	k��pFLF�Oa�sp���$��9�p�����[+�����N�#����N��+�m ��䎧���~��%�B���OJ�����������6/����E��={Ƀ��NX�腩���[jU @7ll�%䁇�T�����l�18PF��1�	�(�I4����"��\�unk|�=��$��ieع�"�M�^��@:n��D�	�x1G��ܜ_l-s�P�CXg�I����s�.Us_���
��	~<و5�}�7I�Ѳ�6���CF��DW,D^���s���n���!p>�Π�mUPۻ5��TD�`�"d[��[�4��&�I�h�.CV
�80غ�Ll���;a�#={v>��t0f�Z�p���n:|��1l�0`a*BD�	�� ��*g1�Xp� �1���*��t�ixjș�R�Y�4�K���2�d ��|��^f|��eK I\&�ֲ#Œ9��"!�R37�3`�]5S�����'p�|(f� އ�!rH>Ս(;�7w�p�."Yr#`�8��aͩ֜ �Rͤ�e�e�9� 
rϤ㑆5�,:�齰آq	�<M�i>�)�8�G���)0�MC�B$�$=�z�?��W:�����7P���={q��C'���p�&��mD6��a�TN�a2C�O����~�O�*,P�fãk��t
.-$d���d/�!� g(�y*�l���"U�U�"���Y�XT�A����SBe|��-�6���WMPi����Ptd��	�l�m�5������I~ȆV_��D�f���(��%$�߇x��cػ��{���4���adg�#w���x�@&�D�K�x��L�"4���|�\!D�2ȋKR%�F6�;00cʨ���~���c�O�:~�m/MC��Bfr�&ь�|���Ř����)h�x�ᇖum暴:�I8�<�	�E��I�i������Pfk8uրѼw׍F%.N=���W�6���fv�DImJM��P�4��d(A�a�>�>��n�}�Mc`1����<%�,��qB@&��U�E�P�)��B<�Z���Ƨ{`�T�e�Ík�9.5��!OL��=
2�ds�v�;V�#���w0Hb�?@����Ǟ���N ��9s>}�W��5���I8��B�m�?�	8�.�(��2n�2`W��ʒ+c�N�be�Ĵ�� �����	J�k�)yH�4��*8+� ��I�flV�ť�
/d=@���Z�2��`��xxM���p��OH����X�C�;��r��--����$�L��U4�'�J�D1q%��@�!���:�ȧ��1�.[�h�\��dG� ���ץwX��=q�ރ&|_`АhǙ1K�Ee�4�
��:o�����[�POΆ-��$K���Ґ-U��ӵ"� ��7$��%�V5��hYǅ�ȁ���c�8�%��:ѵ�k^	NO�3D� �L��9Ywu�0���X�O�X�&�}�j:p�%�� ֑�'cE�'�
P��Kୌ�G�Q��e�.75���r6��<�A�#&��]f���	A����c��3&��peU2w�=}�L�����@M���IT��`![�@�ø�^<�Z
adC��,1��8^F���Z���x(��Z���	�[;
��I؍"�u	'��E�u��j���Ef1�X[# S���b&�9�dw�{�`r����uS}Q�-�wMj�q�%��B��dc|y؎z<�������E�I�2j o�Ew�Qt�T5�\��|fwe��h�$_7
(��Td�򈗐��Ft�ߧ�y- /�J�-����	�J�R2�̙�	�;��2������8���r����R@�d�I�|��,.
q>TĲ�dՋ�*��~���B��qH�2`3<̨���ٶ�j  ��R�H�1�y�Q�Ȧ`��d�0(8Dn��CL���hp��@���v1�<����0��Z< 
pY�HT֠��rKdWɰ��H�D��$��{�y���� �f��d�yJIP@0|`̜2�}�^].�̘��Y�ԉ��!�q��ʃ�,<nS�2
P�����]�b�aQ��p��q_��q�5����p�̟��nX9-N#��3h^'1�2�1;$�sa�_��WE����&XX��h��f<�Du$#L/Ō��%�j vUA�����n4��D�vN��z��-�.� '�x��pN�"y'
�ɧNƔ,�ֳp}`?�׉��y�������F���\��Xn���,/�*	L�<�]�ޝ�)�P/�e��I���Y�� �K��^��@⑋$1��D��C�����
��ێ����F�I�
q��k^8�'�N#��E��ʰi�� �x8	[��F�%G�X�qq�	���a�ɞСD�%����xY�J��̸6�t*��H��T�P�fl�hf����9�v�8N*�#�E>�S܅t	Ezu?����I�֎஺� �����]�a�_���%�p��X(���+�;��ݾ�*�O{sD���v>��*�I%��&�t��/X�>��
�+jp'����K�����v�, ��ع� ��$��
N�p�I o�M����A�x��>��^/VC6���9�޳yB"�
�q�KD���,-M:s%�JsC\%,�n+�<%�6�	�Cn�QTP�lT���J���J���a��ȓ�q���l>	�`8�z.�	'���D��׫	���zX(��=;w�P�����l�\]�*X@��cƔ�����z�B�5�=􍵥Q%�n�0H���J�l��jR�tT�N Z�G��
��Ǳ2 Y���8�o?ܖDj⸞�B>T�#�^Dk�P�rqȀ�{P/����B�ს���w?��x�����l�3CN��MPĆ*���5-x� �1�Ӕ�3�gh�	Z&�!��CB�D'Tbӡ�طk7r�
8 �A��*|�Cr1�ȡ�A���͓=��[릀d��|�MSpx�.��8�R�%WEg�*;�+�JJ7�KI��F>ҿO��*�K�-���Si�A♀!�b1�� ��R�ս�P�?�
�Rb�
	0vI��c׶��X+ ]���Z�Hd,���A� �\��SvW�zU�-<�AG>�ٱ�rҬ7�W	�A�������t2�Y�$�wYt��O���JPO���	�q
�, 6>1�Xr�34���i��b�Ǹ���E���C��VO�&lEU�l����]Y�X���0�8u� 
�(��5pqڰ  X!�Ac�ظ0|�'oۿw���y/��E��2����:a�5�Ґ����ֲp=w �����e�*��Ʊ�����b�mIB�X�M�1�`񞢍\��O Vˆ�/D�]��1��,X� �@H@�\��J�墡2�>
�P�8(n)�C#����$`�� �3.p��;����y�KR�& ��"���"଎��M����x&m.%5�������.@��
��g�_!Z8(��Э�qT����y�D]�wF�<:.�)#�����
��2���q�"�\ɔ�<�z*�Q��D��	Y�5��a��ԣ��X�� O;������n J+Dd"^?�R�.��J�j`9���9\s՘���LM�j#{B�$Wp�,	hL[�7���B���r%\B��(-Ս$Y�2�`�=L��aJ�:�h��r2v�7���}�5�O�`��HN2�I���� t�
��"�"B��`3#�(�C�gz��R��_�i���y�O���\KP%���3xⷥ�̖���6����b�\�QT4����C�2CNg�$�yEt1c,���((�bK�C F� Q�De�y����7��O�㑉8G%��l�G�|�o�7(��_P��>~�� 0(�J�ÃX�q�A�����r47
��P9R2���#Q�8��<;�E��9�粑�d#F)��zap*
y�(��y|e�u�c��^�"��3	M��\
�'�x����U�څ����ɔ�P������%�b�T�ID#��P�N��E���#V�i!���@�cF��(Z����z�*�� ��A�%Nd�"2����	.慈z �N�W~�̤���	!�,Ŭ�p��<q �Q�V�d��Di� �?'�,Ց%V�1n8 ��ⳢW�%�r�0�hxPA�GIX��*"��"W�J�C��g�.X5�F~��&�W�J�3��|�_�N���D�a��A"�>2���5DX(�3�6
@|#����>Ί3���E|���B�c)`F�V�l��P�;�h#���xx��=�qG=y#Vv��{a��O��8�$�)._�b�՟���\D09�S(;T8}6G,�8'�C��yP�So"F;�.Y��Q�UA6�\Qf�c�Xx�� ���p#^�K��r!n(�LE@�T��_wBlP8sCR�+L��h曣Z����o�a60B�$��8/��S�iXN�v���w�D�</1�ߓȿ�
7��PԒ�G	&����w�D\�I�p��T��
�*�B6���)n5>�r*�gn+��I�au
:qY��>�8����,��h��3@@4�i<}����PMB�_$;G�fD��)^��+�����L"��^h���[0��Ʈ��ޗ@m�,��%TI��)#�������T	�n�:�k~Uq�!�Ɣ<�f)�[�f����j~'��*�A����J�'��0��M��")��4c�S�M1�����b�Q*��T���O�U7��K���)v�j9H�PS������:���l�I��Kę�!�[�&��O�g���ĩ5`���X�I?"�L ��p�jR�M�Px��4�0
gLu��Ϝ�K�"`̜��}}���]i�ϫFH\� �2�A��ԇ��E�uZ�ц� bfA2���u�x��-�i��]yX���D�&�����G�>ˢ�-Dϗ0T�m~�n�S��<�M��lA��LRP��0���Z(dM�8���������ER���N�J�z&U�E�
�XT���>V�
�(�Kd��P�Sb���d�I�!)Uz���p���=׻�y}a�1�.1.�=�	�ҍ��O�ʙGA�.Q��t�\]&^C��ГMB�nLI�ؙ���3��$�M@�I:���E���EH�9骠B�I2PB��`V�A�l?����`?��9�	��榝����0LC��-:e�%O�ĢQ� :EF���u�L����<��L�G�����GX��3糖�R���ZK�� !~��!���jHE��r�`�`�K#MF`*��L��,1����S_+�5�P<�]0������8R%",:-��efw	�n���f�	$�:Ȟ0�c����]$�B@2�"m '��<|��2�i����I�h���B� �Fz�ٔ�W�q)`�|sx��}��w*R�!���WeE7,��C��eC�QsK���䇹8t�?Ȁ�L�ܽ�f>�/��z�b�,xƧ3%G�z��!	�<#b���vס0��R��l�B��ԓd��,Cv��f�Dd���!����ef��]�%� �jp�wa�$�Qy,}�$4�b,yY�\OX��=�,I����b%���6	3dh��GKOM^h�L����G����Aכ��4f�hSi'kP�B&E8�O�a0�N�3$�qd]�dҘ�& O��Az��S)��RL2���D\�c�71�S�i��)�F�2�`�X�(T'V��\~z7��[K�˜ky>f�8Q
B��C2����Ye`p�׹���f�y�?L���'uB�k�03J)k��):J\��]4���Dxyy$h�H��b2��w��n�p�Z�q��)d����u���<���X�����,j�����=[��$�.�."c����H5���)�,�m5�M����yS�7X�g�q���    IDATY��[$%He�$#�?��x����Q�N%�f��2�fRހKD`eQ�57������I�DX�S�fr����\��h����H���o(��D�Y�{��{�0J���O�\�����4v`�����2���Dp����� ��F�IƧPX[I�����x�dl�lA�,��U�(«i����A���̳,+5��9dW
�E�P�EP�U�WĈ;D)��l,��nS�EX}��aJ�ZJ��Tc�����\K`�3>HD�@��E����Ɂ�^)D����x!Zm���q�𞝈r8 �����B�nP�Z����,�I"��� I���U��<���N!KqB���SY�������� @��6<���E�� ��^�����VxM@�G�jq��9�āW}�{���,Yf�Vd{4X]ь;"
T�\�(*E���?-�@�s~�,V�����,9mGAn&��(�UEIY�����Y�vfԒ4
�|��oƅ����eIb8H��¢	�p�0����`�ZqKEoiƴ(#�[�P��ϗ��e��A���.� dʲz�����፞�3�%G����r�gǬ��bh�yt8�R���F�V<�
�@���En���Hĳ0�����Ywb�b��GMn5p�RC��dd4�Y��$B��rq.|n�K�/�2�
�� �8Y5��"�lV��d��{�s�B�0x>�� C�,a��K���1����
�����E��IEH_Nzg���.����b7�5f|�?m�^��n�d��b����W��q�v�(�Ω���1�V(�^;Y;bccQ%�@�u�fW�T;�v~O!��*^�lD1���!�TJ�~�� ��摗uN9 �+
^)�-��B8�S��T�0�����8��6SU�;y芟5!�a؝.x��@S�QV��L�-"
�

Ir	؜�,E�\N�șR�^r���Q,֤�JJ%,Ui`�8���
fX=�.� VMi�Ç���w�m1h�aܰ����1���84QB�Chz�c��Ŵ���K�GBl|~�%�� wUv��7�_v`���3U� �a@��E�
��,4���)UY��[�%������%���w۟�S�F4��d�1��w/~>�°&!ʯ�)�y/��T�W$��!�;��l�����=����x#*D;p��l�{
�WLA��V<��N<vo\9*�������n'���m�j\)�D3�-�J�r�0fLu�C�euWM	q�D�B��Îe���t�M⾐s ���()B��_Ʌ�����`��u�~@v�p�F�8?���	����F��Jl��u_������ϻ�骓X�t�
7�M�iYb�?������a�kϠq2��$D�!��� �}�dWn���t���7�Ѩ�y����E;�y��EeK�"F����|&�N��'�2��0C��fY��B �P�����X�����jX��wtz�.8�砟���Q�6%(C�H�F�M��1"�ŅP����80��4|5�-N�00��5�v4�W�Zj+|�� ��}���Z�g������ı"	~���@$(��{�(^{�-Z��ؑ�����K$���3d�cd����6#����i��倡/<��7CF|��X4m�Þ�A�xb�WP�D���O�6h|+��W(�p�՗�⦚@�^�#�H��CŊNp�
�'�%�x�ջ�y/��;+� �ŏ����V��	�!W�A�D'>x;����a�����-&VI�S[%v��b�b6� �,�.aE>Kgc�,c��A�_��o��8���K8��,�O���CX>�N����1	I�����������l�j���д��7ǰৃ��*�X �6IE���x�#��>s/�+�jg���شu?gb�,x�n��q���
bB-���D�1��Ag|�u:f~���6�˝+����ps�
��A��1�B-L|�l�y��	��#F.D�\�A0�������hy0x�R��p�Y�:��l$�|���{�ɗ�h�AԬV	s�ނ�Na��D�D���[�)(�e�II�X�p�ˋ�T�I1�s�B��m��,LO1�m��Wy$���ހ�cּťf���.��d�h3�q�DMg�J��N3���B�=���"��Cg� Uv�A��q/݅� P�$8�X0a�/ظ�(��ZX+�Ч���vR�ɦ)�/4��y*w��O��~���20k�T����6��H�y�� � o���G>ޜ�5�5o��g�`��?�L;ܼNA�uQ�tޙ�֦y`�;�Ψ��(;_~�	�v�+>��g�ʨ�Q5	��\���Y	7��wc�̧���6��\����~�;mʅu�GdN!r
��*�����e��ja�;�Κ9�*�"�f{
��L�OC�|����g��w�|sؽW̕�%�f�hz3�o�f�"��Ҋ��:Q�H�Xr)�E�X>�$��S�!��u��T0aP#��t?��v5���3a�a`�K�UD�_�hs��5���H
��,�ۇD!���y<=�g�~9�.�ۛ��E���' �Ն3g2�v2�>�Ʒ7��N���Ե��ޕ+�G�
���M7e5���Mj.?mZ4Ľw�@�x�D�ikp #��tB�$�g��V��^��
�r����[��Q/^���I���������Q
�x���P<���STMoVә݁��~����D3;M	>���:� D]a=G��L�&����o�r���`~<K���-�|7Hc�L,�W�k�`�#
���A�M��qmp����o`�������8�)>\r�mގ�BZ�����������-G��*2����>�t�����0���r.�!���kÞ��{�v�>��V�t��We@�B�T�F]�D�֩�W���7�bO����+p}���5�����2�(X�~�"�Џ�n����S�u��Wf���=��7��}�3�Z�U��)D�X�%����M�xuc}�? ��o��>�qp:y���)�JYZ".�j�X�~0�μb�ӹ0Av<�6Xc�S<9�V��בD=��P8}ʨ{��z���c�r%��2��f{F��Q ��Ϻ�ؘ�O���a����1��� ��q[��i��?=�����dx�{�oEy��>�Wۍ��  �D�5zMrb,�'1���!��bb,`T��(��Q��J�}o�m�5�f����f1�lr���{��/?vYk��{�Sښp��Ǡ[W��ѯ��աP�H$��=PC���\`!�t�2�b̩G��6�+_��uM�z퉨��z�ch�I4�X��-z�ի���sg��e�������b��f�Y�q����n}7�ѬőN7�[}5�LNf���d���٘�����3zcƓ�1��9��H�����8�'&�p�;��"�}���w���,��s���و�yD��lT�
 Huv
A�qw$m��{(dp��mb�)�V+J���9l���g&�܁����RVo�ō��"]KS`����pbpCj�h0ۖ��~�ukC\pǟ���Ǟ�\}����u���"�t���ڽ�\8�	�>�U$�	���������c�1�� �M�vܾ��Y�_>�M���>�L��� ᷼��2�2��ѳ��Z�i�/�-¡������'~�W��k�
خ:����%���X�`Z�w�Ǳ���}/���]�Љ�s����Of����������|�5�/�L;�j�����`�7i���f�8D�)�k7��+�}�1*bs�Vj>%ĢP��#S��'	XKo��afM���ч�{�ɟ�_�^�#h߷��A���CJqF1�Je��(�Zгk0ᢃ�ry�_�0m����G�\����S��bA��w$v����N39�j��f7`�I����ѵ�Ud}`}+�����ݹ˰^�AU2�[���p�	?�N;*��������}
�]�~;����{	���mo����c�	;�Gf�/��G�����L�:��ޛ�O��v��S͆�p�ч��ú�*4n ���	��fu7�;ءg~}t?<��\|�,#�	a9/�	�.�궫�}#\A�`���B�sS�E[�& �H���JIP�m���`l�v߸M�z��^��-%
$j-�R~{#�����:#W���,�N99�M^s��$�V~��c�S�(����Ba�n9�B!��]%����L��B��j�Վ�ֶFxe6+� ��Ч_����-L�d��e8��ݽ+��V��oB}C'�c	��[��Z�e�䠐P��A�J�V�mCn�h�&���_��J����:\e��",听�C{فG�	�w,Q PmG��E���A��p��X"H��E#z�J ҜiT���d���ɷ�:��ߝ��wf���mM��H��ٔ�*�3E��@�z/�4�vL�ep#�74��H�P�\�^��"րnZ(�J�c����h!�%O����8�b	�W���V�%�h��ajUx�e�ښb���2m>���t3&���Dܹҏ���X�d;��x9�c&JtR��(����F�YJK�P�G:��lG��!���x�$�fR�|�ݲ���	��	����Qj�p����'��L-E�dmR�$U�n��1���1&�ҁ���>���9�����y�d��$-�N�+'acȴt��dWA�-�mn����
3���G6�!�Ƅ��#l(�uUӰ'ס�x��v�|*|�Y�ܶQ�J�S�6�@��]O�4x��\�\l���<�I�7��䁍�z�dP`K��""�<Kn<�<bF�ؒ���U:���(�]L��T*�#�E�"�� �]S^�	�� �u<(� 33e�Q*�?C�1Q�d[M�s���!�������7�CH~��e"��7آ	-����W�oƶI�-��!��u��x>�)�f����6TgMԷ�	9I�o���p=f� It���/�1��K�G�[3\yR��!�nh0��O~��9��Z䒭X,J��m0����.�E�%�տ����!,g�f��R�@��-@gG�qHt���'�uHPY'��Qd�P���E�;���|^f�cJj%�M��tb��N�,��QN�^�ȖCՂF�1�kW���c|��h�j�(R���K%��ǶL�t״b(]xAI���'���Ϫ��L�$�.�\oe1Z�IV@Wz�P��u�✘|�i(���h+�$C9�	![y��W��1C�AQX~Y�wT[�ZaHU�DL�e'��t����d�"D@6>Qi$�9���Ǫ7�D2[�Q"��V"�A�U2��䁂��#V����y
�<	�0p��3�U0c�eP	 ��ј�R!/*ER\:@�'˂K{�h+�u������|f&�|ɖk�)�>�_C/������!���	S�±SR"��v)'�1W�c�O&�-����8�����)�D&f_6�B�3����(���#H�g\1�q;�4e4��T !z\�.ȶ��ݾ��:L�$�/R�N�W*"��(�����tH\���ֶP��4D�e��W��u(�T��ĉ%%��R �%��c��]Au�A"��b�E�ku�ĥ
ZK�����\}+�C$j�F�at ;Y�t��/���FC�����nG�ן�~���Q�Z�+��. ��z b��5;���Ү*>�~A�V]?�=IU1�s\d�H�e���e�2���B�g�@	����6����L��;�z�=�tx������.���%[ذu9rm+�Y�����(R=?��J�Z���1��}7�2Pg�%C�l����X��2�f�`��T��mҷ%D�+�E���kuEu׾(���ld��I	�-�L��.A�V؊��M5��{������P0�P�g����ڜ9Њ�Q��,�
ꊆ(�_`�`����m��&��D��bB����R���>\h�*l��P�{ �e�%@Ls��rff��/�EˬH���ƀ(N�DgY�`x����]8=�����Ku�G�9W�e���p��b+��J����1P΋X�D��=����s�bS��?O���@1�������2�����S��/ zFv7`w�@c����z����8��?�4�1�W���G	�s�E�O!Ձ���$Y��I���f�E!�p��Opc���Q(�b�LԘEH%9J��1c|zǿ!cXAU�&|6����cp��=�d��|�vL1�\W���$V�g1v�8�<���?�F���ܷ�P��<�|�ƣ�g�8%�(f9єU|S8�=ޞw��{s�ԋ�q�Y�b]P���!08����8:mh�x���q�Ǡ�*�|�m%S���W��e#!�SO?�O�n�.GCeyƓp핑r$�"��,v����G�+�����{�$z=pᖋ0l���'^�����Q�E�Q��fɑ\��������gb�������
��I���S%-�G#k�����%M�v�c����T�� 4���cף)B�JIԇ-�=����5�*%��h-�u�E�`�Iا�g���b��y��ȼ�I���/�N��A��P�네3�����������1��?�� jw)�(k��m��%�$^�KL��"{��)�,��z��~�~V�}z9M8﷿��0bP��,�T�B�d&�1��'��7-���+����Z��.٤�N/�ӗ�Ð�&��ݱ�9��C�84NwI �4�\WP�0�x�Y��4���9��i>0��5u�$^Z>k^y��]/L�
�U�]���CA���j|2n�n*���.��H����2��C�ƽU��i�!l&#s��K�<ߚ���s}y5޻uι�D�kI��ܒ~ԨL813m�/�!�<�*�=a,�>��Df��������ܗ����0��?������JA554���o�|�<��d:������mH����t
۰���7��O��� �BG��XX��bP���G���K��㗗b}P'��m��˷�������0(���c����������%'�(=�׏���=�qH$�N��P4ѫ�����������a�%�����A��(��TU>�|>n��A�7�����#ű)]�(橮$��-iW?�cx��ؕlm`P���	W��O�A�v�
[�8�}��b��n��n�N=�bl�a���@ul��ٝ��r3
_��E3�Ľ���sr�^!�G�w��C�������ć^��LC#:��'�&�Ð�7�?V̺=�\z�)(�R�G�l��lT��-<��ۘ��~z�zW�%�a(PL��b�[�`P|.<�h��,J�{��x(�B�(�D�������c���E:H�d�����!j�,r�����'�����Y٥2�i$( k)�Y5�v��.ĵ�c�K�Z�f��y��F�
�CK2�nz��Ç.���}+F��U�o0{�8�̟���n�R��J0d�� _,�w#��N'�n�]���/���o=����.����U`�&&
ӌ�+���G�c�3��Yw�I�8�F2։K`�Κ�[�Əu�O9^�����nR�������k�t�p	��C��rXF������=�]��8�!Α��L�GG��G���'I\z����W%��Yh�(0�Y�	nM�An��X��$<0c<�0#T���^�v��̆i��}�?����h:�esVS��9ͷ�C7<t���;:[#���训�[�/A�6zVs���8��#��T�$�d\�m��9+����a��[�&8̒�@�'�d��g�c�돠W�ZQ���O����a���L�T��M�7�1�tkD��*�0c4|���h��%���E�n�-�uM����$%��A����v'��Xl(שVT�(߅��]w1���W����@)��g9P�!+.�Xt]l4�6]    IDATZ�G���=�d������	�*0���#��N��$!8w�]" 0��eőI�֬�2����"�r�g¢=�f��Q��#2�n�|�@���N�2��倷��ӈ8GC9"���'���7ջ��(������>���� �44��$c0�G�Mōl��z�����J�1����)��7�OF�{��K�
�*oL�����
)��j���������(��B�́[���/_�抗p����e�2��t�n�$�NSs
�W�ÂFk��߯G"�Q���-�d`�m������Nئ��BlM 5�RZ=p�$�����Y�A܇l� �=�Jl. %��g?W*r���#2Sƍ�2�ok�:�RcL��Y
������P�{u�D�^�\@��2u���y��w�ᱏW*;�$qL�����}/B�d5�$���u]��P�6,}{Z?z��6(�]`(�;Ճ7�1���h��Q�Ff���Z�c�;c'�K��!�٪(d���1[pc�����o���6�S.C[�V�y`�-�-x������
Ze�*�@^�� =��ɮ��kZp�3��ЩhM��zEށ�HW<X�>[S�B2��!c�K�A�o��Eӊ�� �E�/���t=n4�|�|5�C]�@mЪ2�_���xE�>c�I`�.�V/����tc`p���uT��X��T9JPhS�+Jn3d�o��p�a�?���Z�h�Dƽ���Z�a��b��|�8��\��v��.r#�IUk�������C�þ�C�슂�XJ,�J�+X��x��?�����f�!��F�k�1|�]x��T��pK�:�)_)V7k�.�:̾��ck����G�Qbjō�sN$%}tbYj/O�	�l��$1� �Wc���W��lW[T����Ӓ1����(ql��0m�?̞�k�#hһ�d�Na�Д��1mt�rX��$���� �m�K=u7A�T`��AWs�C���c$0Ȱ־؆%c�k:�H��'$AL.-�?�dZ��+K�/{<����U���E8p�uh��Q�و⁰]�`nn�_��������7�U3g
�W�0�V.o���ߏ�gޏb��pEԅŪjUU��L����%Ό��_�Y�������F��hYf��c_�b�fg���eH�t |���\�X��3��KX����%RXE��'��(�U���$�%�e��֎%o݃���_6Z�o)c��<J��NR'>Da�:������-6�O={)ӤӵHʜg�{�rM��xa�R<��2|�x�h�ȋ|�rT��@������Ϸ������\ps?�M�!V�FkW�1�ҩt�d�v 9z"��Y�$,����l�J:[C8����������|�΃�=�.<� 	���M�h���!�!����K��c+qȹ�Ь�6v[��6�翈�/܊�R���U���I��r ���&��L��
C�ƣZ�ہQ)>�gq��}��{�}\\��#z*0��c�o�c�D'���*��V�]���7���'W�a�eW�)c2ǨC�
��o�\�����G�dZk$$0�����}�Ԯp�}*cc`�(��O�1�&|8�5����'��Y`l�^!v��o��Q�Q}��c�;ӱK�s?y�L.��SGh%0���3�%0z���=�Dʄ�oC2F�(QNӢ�-���}����r~�!d�v���^�"5A��*��%�����*cl)0��І%o�������of=�]b���S��S��.���&Vn���-#�g�X���^�μ�F�ZLىs���$;�%,z�VL����ƈ�π�-�-����vu#.���{xc`���f<�X\	.�v�0|[`�;���E�?��x��r�hp���ܩ������Ģj�x�k<�\#�=��#�(Q`]���7����W�A�ƨ����/��ƚ��(r�ChO@��*���/+̐�f�(08����qS���?[|n���]"-�h�!����(����ͬ�%1眰?b�n�$ ���R���T��*O����ԂCϾ{��0�!���ƌq����I`DXN����5\|�r�	�"��� �U����c����jծ�WG��q�TsW���x�Q�nǏA͎Rn]�Ս6!d%����G��g����sc�*����yMܮFʽ�I4�����7�`���C���f��l\.�L8 �0w>�~9�A'AZ�vՐ�j�YƂ����g�boh��"x��U5�㢫H�.k�x���x��=�FlM��Kl�.]I-T`,~~n��<���;�!s	�j�F����hn*���f [����*��H��H�[�0�%wt0clu`���u˥���׮��
�D�@i���Φ
�@����	c�;��D��Q&G�z�Da���������̀p8�D���� �L����P���^8`��X��;aœ�������q�0�E����J5��X*:)�X(�}�tv��H�]a�`�� +�8u�,���ͺ(m��nQ�{8	"A��ϙ[9Qt=��8=!:�$o3؜@C����YX����(T f��m:x=��*��C�`uƐKF��[��U����&�Lc����P���1<�!���|�yԖV��)�����Ñ��Ќ�4�0D�����}�DJ1�`�̳Ǣ��Q��"<V�q��d>���.���OM��i7�*ge�,�]�����cq���LL������bu��0�sՈ�4b�<"�6`��5}�+Ǝ���%]�D%���2�MA4���<�����Ϯ�t�d�Ő/;���JҘ���(��Pn�n[���^@X���iZ�(�C�z'`�ð���G:��lR�}�cA�xi���c���&�8�%J|��.Ǽ�1X�eW$,�FW�>�N�]	Q�X_P,(����C����FW����/��'���iׇ�,S����1�D!���:�3�^��'\���{��ɹ,&wT�R�x+��WON���7���&Q�m|�Es������[31m�+8l��X�s���+�	��t�f��wr�?��7ހ�����7��6��$P٘��s�˜����[�5�����<�q�bէ/!\�
���2.��8
W[e��{ �F��W?���b�翇"���)nw	��׌`�{�������"�N����^�!���������и�<���06X=�JMXW�*2��i���d�E��[�]%����s-~w���>��0�O�N�-Sp��G^	?DU���`�IW��;�:���g���!��ފ���wb��7
�U��h2P	7��ƛo���z��=��t����Y6���d:�����B��R����:�nM�|Y��1L�Y��4��^��F�b�������ki4��+�_<�i׏j �°�
�Vf@9ЌLC�$�>�&^��{��9(�c�-M��@��_��z�VL��F$��rW"Z>r"I�$�S@��͝����C.{��9��_!��5�%�a�n(.���YcL��#r�[�J�x��
sf܌���$O'1���Җ��%��ō 邇sG^��']��n0�<i�-�Z�Q����]�}�nL�~���hW�5*�c���)+���x=��>���]ap�	��j��Q�7���h]��p�h$l�|^p����@��`Oa"``<�>X����^�f�q�\� �]#��x���9o�<�\{�Ŝ�tX1d�98���� �g������
{��TC�E�s%�"��E�1wL�Ն+�!&��`��D}J+-`���q��ǰ��I�$���hZ�0�Wծ�����gv�͗oY�sk�:�NF>��z��ȁ8���D�F7
��ȵ-�����$�<�Jl�eH���+��LS.\��
2(�x�w30�c��K��z��2�$*q�iZxc�'x�Y8�;�����?d��P����P���/x7����F�����`ծ�M�l���䳘��Z�s��h	����h��^��z��(~����r�6�P"�1���J98Ҷ�¾��ԛxc���q6�<e+!�L�N��O�[��>:�M�*��R�n�w����Z���/>����u�DdR��Xr�P�&�3c`H�U��]I4��Q�52��׺M��;��z�B�{��r�>��
�F�1�k��/F����(��7����OF;r+>��Oލߏ�f9#P>���� 
1z=��{}�'��9�;���e��� �8t��zvγhZ�.��L� �`(-�1p�LN�3�^���Vf1��ñ���G$��47���_�	w�L\s���͍�M��x2&�~>��GJ#q'	����xk~��rZ�*xvJ�	nbƬ
3pW���L���nAJ��&��h\��|���O>��w=�C/���ZvJ
Ve[�D�,,�EeC��H|�ٻƏ�ѹg������?P�ٚ� ��m�g�4/�P��\�7��*��h�����w�����"����5��kHy�W~��OL�,@9A�0�s�����
�ͦt�{�~9�5ZY���PS�;�e�9����y�)�
�z\�i*쳍>W��ό������3�E�������O��Âw_D~�Ӏ������Y#�+�wJ>k�w���Yhu�(�D��`��D�5_�GJ,>�AQ�d�.�]�l�M�����7!��A�>?$mG���䐋-�V���W�(��_�PfI1�*1']5"�Q �ݪ�!w�SP�����p�6X�Cw�$C+�JǮD�v��m��I&�Id�:x�S#=O�O��LCa���3(�����Př:��� $7��L:-w�'��������H��ڡ��dh&��� �K�X�{ ���q� cA�A��,�X��6Ӣ��+߈r�(礫���RS���&
�r��%��V�u������T8��3�>F�Av%�]ݚ�PMlK��s\�E�vQq��"G4?�c��Z93%�����dh�	�D:�t!��%�>DBHɂ��Z
�h,�(g����F�r�f4Zbmn�'{J\��4	�ȅ��
�h9+%�9&��X�j�S�G�\D�C�D�R�VY��5���j�*�[�(MPC�5��,^U1�4�*���G�Q��5=JF��O��K���HoDv����F����N�����KYT)Zn��ۡ��QZ���O��dq�)T�@���``�W�GR�\`ZaF�!'KD2�7�!��vI�óU<\I�*?4:-Ẁ%EYC��5��*Spefǉ!� �d
�� s��nW���Vv&JF��7C��L��>8�si���wM�2�4آ����
��+�X4VG&�Id�DEHyK��B_�B�b�A�N�&|<���qc�lή�a�8N��LJ�GE֖�O8J∁$fp*�q��񆋰�����	�;(F�h����E�1A?�5��Qe&U�(?CYw30x+6mJ���r+��H9Ϡ���d��qE��d@�x�"'�x�����H�Ӕh
	?�A�h�G?V>,q���SX�>W0��uTΚ�<�"j���=l�"J1�;"Pi��cgS`��K��e�q�O�9�w����羇r��^�p���E���+�n��7F��se,���QN�܍��<�B�r� ଟ�H\�g��cD�YX���� �y3U`��T�/t��&�b�RA+�e�j����<���Zo���yLX�|<.D[e�d�<�|���`�̈M�q�������J�F�|VTT�#Z���f��k,�~����U�%�kb���_��F�0�Y�D�v'�:Jd���?0$��jW���RW��M�'ʶ|���QGwm'���L))FUᤊS>J�J�C9�#�J��O�T]��U}Q+N��h��Ŧ��V���C*GG�1(���a�5��H��V��,<�� r��p�$yE�"_�~��<�f/Z�c_�1R	�cS��UQ-���QD}~n����/T楊�P��7�j5_��m�*>͍��%0�]��0o�|*K�
kL.Nt!7��Q�D\L�F��H-��,�<~ʏ����0��i���>E�x��,R�Qe����Ճ�o��0��]P*�D��v�v�8:�虁�T&=<�:\I&(}�YI%}Nf
�xx|H���[&��F+1:�YC*�Q�I�-�3k ��{��M���T���Mq7EƔ��*G�a�{D�I�ԋ�Ht�5�>�L��2~�k�i�fy���_���$z� Fda%$ y��gy�� WD@9R"־ �&�|�����B.x�RE���UlO�K��At�J9e>i��������.���{�*y�6�n\Ή�w���@��ZW܊����}��V�P}$�I^f&Փ�5��B6�Fbv$�������fS�j,�U sr��ḷ@�����"e�����ˢS�g�L�U�*���Z�!hפ���x�'���o"�m�#	��ƿ���N�W7����sjE�&�6�+ ��_Ԏ�8�����eJ��w!�	Ӷ�泈9Ԩ����F����rY%���!G��g.<7�H>�eU��p�u���:M��d�Q����S�CPwӎǐ)����e����ԓĖ��\����J�@��N"��Fw�جZc��0�(����%�^�Ϩے���Q�]�Q�ߩ ��3T'�^�����p��ZLJ�D�+����~��ˎ� Gn���:z	E������)�;��<0�4"����e�w��=�PB])�����/�p�У�gY	����ؘ+�q��P#E'���E*���2��)����Z?�[1�G�"�T��ȕJ(���;�QA���$� vٓ��O���,��*�b�Y������ి�WZ�ddN���rQ���ř��9Q��/X�Yp��y��ٕZf������k�����W
08�|)�):P<�|T�.�&l~��e,����}�y�:t�ɟw c�$�I���r��(zE��h��PcI��>)�Y ��E8�����l�[�s#6��b>+j8��EN�"pRhn/"��H�yT[�ީ�Y�n�RI�VR���� ��D�4��"h]���!i���e_d�S19��t�o%�C=z��rU�0Ljp� �����D|U�ln� �K�А��r������m�U��j������P����t+F�(q�e��P��ކOo?==����)�30�L�q�ЋT`�G��,ʬ���վeb������m�ߦ~����5��D��jt�H��֮Z�uO�n������) Ā ��/��^�\��;��mR3p�W���� ����ߧ�~���g����? ^���m	��~:����g'���=��hhk�@=�a���3b�Ӊ��bI����{�V�dQ(f�b�����؄��
�$ߑ?W6V;���S>����IU��to|�2 �!t�<ЬYX�q�������a�n�h�s�8��-�ŷ���wJ`���<�̟�}��?�;�E\s�0�n�I4���E�[����?c82f-��.C�����᧣*��!�=����m����Ћ�AZ�F,,�����нk�,�x\P��ؒ�0��I���@�'bz�O']�a瞈���F�Ǜ@�=��6�K�n�Cp�1Hl��}GIOS����X�(ss�|ci�r�Hؾ���~�Ѯ���Yx�F^ ��TZ�ʤwk����r:.��P󞲡8V&*�]TQ�4\ɦ�N}ae�0kҘ�)��w��n!0=r���7F,Z�t���q|�.~M�&c�u� ȳk�P`�Ӱ��9��F_�Ç_�l�;��E�;�q��Q*)�5�I���_���u9\5�&0�jd���i|t�Y���PW�I::'��J���>���$h�,���]�\w�Ht��M�b�]�_b��%�c�� �Ͼ�Z5���^JY�F��m����o<�`��$������b.�,�D��ǯ�АB3*Z��T��D���Qc\v-���<�Ja��F��^����)�H _n    IDAT��r`L��5���>A2�Fw*��qѡ4�,¦�X��͘���ÆǳMv:V�p��q8�?�9�-K���`�b2�v�w�"eؖ�ōy���Sq��k��o@����[~��:]z�Tn��}�]Ӏߎ��G��t��Pk����q���SC� di�(]�����.����D�Aڬ���E~ ��5���%T�!�~�6r+���N{��������R�t)�#E���������V�r!Tn��a5_2�ć@=M�\u�����-���F����愑�S�{�g�����.�7md��Hī��K��c���q����2� N��� vqc��D2�hKl��_�p��I��9���N,��0e�p�Tr�MXo�@�܌�������.]�t3��Db�,�4g��=~<���V����N�M�G�.�jmz�5�� ��8{�x:�7(��mV'��!�r¶��J
��KRp�9|3�֭��CQ"�?g7#�P����;	�������h��uߴ�Wˍ��7����۰��u(��%> l�"��D��a��/��g��]�O?f���>i�w%��y���G]��!�!��'5�$P�*���UBn�L�|�6<x��02=A���t��l��އ�-�Ѽ�+�߹��*O)�8+U�|����a�~�$6��	��[���ᦫ���[7�+(�H��bX1\x���w��ж��b��y6n�r(���	ߧ1�����A1���+nĮ�ׯ���j�2�L8�kg"�5U(b�ϡв;>.�n���Y�W��+���X<���+�Ҏ�,�Xl��L��r���"�Y�f��?F�b�YW2l����n���-v%*0���!N�zԉ���q]"A��0���oc��ɸ��+��-]�h�h)��e�q��p���b�����c�_oÌG���#�K%MGm"�EkҸ��;p�W�X�z~>��t�t݅���C2'��o���bI�2l�����:��bָ���G��s��� ��I�z�F\�}~zܮ��uF.�e6!$��إ5�c��O!�Ҍ��OKD��h�(��j�*���\���d
���o���h��� Q�r����2w&�\�O+�O�Ƞ}��h��)�I��w�<�}��1z���.>�}��]��z�A$��q�H�W��Ϟ�.*2J���N�c<�i�c�U7��F���B�j)>Ǐ��,Kj�`�r	�(����f�q�yi�q����O#ѩKW��p���i� �sɕr��ﳏ�-�<�R�r�p��7.#���������O|�Q0z�\�rNg���'��U�6�a��#�܂���	\����Z�݋�W�[�"��ʪ��q+�cK��nį�*"�c�U�SE��V8�72Ȭ���9�c��k7|�?���I���rƘ��މFԋ�,�Ǧ�"�r�x��JM�.��#��[P�P,p���C[��ܯ��?%��r�V|��A�vqF��[HB|��$v�y$7�(|��k�uie���+kh��;}���;�K������y��CUu��Q�.�:C<��y�=���Z]_R�������wV��'̰��ȥS]����E�����%�F��j,�\"��R�������޶�����T�&E�BU�wZ��d`�H��ȭ~k�|�A�ƉM��m��Ʊ�w�	�;�1�~75r:�|������ yq�!��2c�+^X��S� ��a`O��� ����^�h@f���*rT�*�����������Wym��y�op����g��9�Y��O��M:��[�Z���E�^��lK�r
z�,��U�R䏋�����Q��i��ŕt���
�韼8W�Qo@$u����|���H�iV����nD���ĳ�&�u���{�{��3G���>L�F���y|���(~�*Pj�11��!��Ӱi_�`#��T���-�~$��L8�ݨ�Z�ԱPR���M�'��'�X��^v���d_��~������y2�R�sz��w<���*4y5HF�'ї�3c00x����g(j��J`Tgj$��Ѱٗo�P��e��E����^S�6z�S0����QQ��MT�mȯ~Ec�97#n���1��1e�#�9���O��A��ڰ+ߞ�?[U,Tn�T=j��p��1Me�
Eo�����4��=A��Wc��z�	eSs$�V,�D�5V󏲌���B�ΫG�lu�������5?G�
:g��n:��Gl
��<���D_G}؎��@������V�By?ɵvEZR�6��Q[l�eC�yM�Q;r�ȕ�����A2�����&�FJ�^Ɗ/?��a��1C̾�ܶ;o}����E�����!QX���ߏ5��EP���iM��$�@��ʲ�B*7K	H�/b�*�XL���h���h-�D�1sk+.F�d�O�	������E�1�����U�4A����@��� �_�ɒ��A�09J*�d����5��ϐ�E5�ڕT��Y9"3G*Ҳ��M7D��:rR�����_�
C��b�QGö��$r<ʨF��D�I7=���hcq��j��ȶ���ӑ�[P\�*V~�)vv�pwgO�6��Qm�]�z�?;����s�9J�%袷c��w������J�<*�Y�������Xe���:z��#�n��Q2Q��+�o}��n�6
�Ejn������=O�f��@����y�}������������<
%t��a�p���"7�j|^q�L	��M�TA��(�@(��O�Q,{����d09�Y�T�������!(;ΐ+�2}1���.j�k�Q*����]Wl?.�X+;J�Q�GU��.i�"��-���s�~�8�u�(�)�F��vu�O�쬋�v�᷋!
U��X��d4}� _Ā~c���&����6\Q`D ���S�CJUc�������lt�AfxCd���lW��d�=���D w�C��r�(�[ø@�C%�O{��Eo܄���hZ�ɺ8R5�ZĬ�̅ׯ@�ϡK���)heq-@�m��M�Wա�~�~��W."nSۣ���Ĝ�VJ���!�������wb�"a�!��]	��î��������#�=�-0: ZDj&���.��$� LG��Am*���q�b�N]�u�V!$.��G6ׂ�_D�>}Pv������epةK7؉*�3��H!�H+�ǆ�b'KvB5�g��e̱���H`�}�Ň�s�o���Q��|[`t<c���bNc�%e�+-&Qd6t��$@�Z��������%�;%�HQ�\C�i���	͙ft���U-{�L����X5R��a�q�n ǈڬض��ص=`�ꐰ���,il��2ƶ����EdbQ�J,#0���D��Cw������"��:��>GU�ӱ�f�R�.Q�9��T�����k_J<��g�y�X��ֵrĕ2^�K<U��E�L9'lE`�O�e�!g�~ʗ�2��Vc��͔9��3�	����ۑ͵�h�[�ż7���K�h\���z����~{b�;!,瑬������,�[odJ@]�t0�^��b��ڶe�'�5�K�2�$ I[� � ]�t���X`L���qC/���m5FGj��<�E�̒#@!�Ќ\a�����n@��yX7�E��i��ð��H8:���!t��HR RH��X�f-&M��Oޞ�Ԡ�ѵ��j5XղN�
U��H�k�20ȋX����-0Tq�q��NWB7���(#�s��mhA3��%�
��ڴޒ/D���}1��Y��t�2��k�����r��q7�/~Hv�vA��.Ы�Qݝ;���Ȓs
>�f%�q����e�m�gǋO.����Lő˷�n��Bz����n��/�Ev���i���'�
z�ҥO?���Ԇ6<�G2a�-�ʮ��;'ބ��yI��v�%�k֖�������+Jb�ǀ�ʐ�FB��hJH��]|n��{��� ���|#�$��!��)�cݢYh�`�;dw|��,����pvۡ�?�ڮp�	����T�
�n��?�$vؾR�:|>ov�7�7����a��G�h�@10�1������Q񹱘�B`�5~���uҜm���T|���	
�X�~B��TM
u5lw=�~�~@[#׎�{�C*Y��m/u,Y�5vݥ?�|��;�X,�;n��=�,RH�-��yTW�b��ň�vG[����T�G��i}�X-��pI�)nޕ(��p�o��]��G�F��j�ge^�Ѻ�t�3�塃1�曰]����j`��siT�m̝?��&M��rp�mwcƣO���3�V�/+ee��_�#~zjz����?�����������I`P��(|%I��%0��ķ��ಋ�������V��^�����57��Q��in��ӧ��v���HC�|�,�f.~pȁ�a���6�A���V<7���\Ĭ �����W�m(���OD��' ^������D���@qy�T���1��Vo��X�+=�G"��^3kg?���<�r	5	wO������N�z������KX��B���ؿ� �KG�/�tt,\����wO��{�~�����p��GB�h"@Ae��E������Ə>d�5ƶ��x`��:a��Cqo=V}�:���b��W��n��X2Ҿs��x��ѣWOh�rՏ��4��B/�Ìk�X�p!v8wO�S���୆�_zS&>��G�����^#��[�%���m��q����U2��p�lW��liٴ]�pj�N�
��2Bz�S���Q��aeW`��᷿����XP��a� ��q�ģ�>���	a����!�l���F�f�B��q�u�4�$R(�6(�����e0�������Ъu������U'W�1�*�@b;h ��G����[F�ő�^�Px���j-��x��G"��.>�z^��L[+�f�&���r��FM����^���g��]+�懯�	R��*�m���ǟG���#��R��8�X�r%z����M'\����Q*�D�xyc�=�|�8�8��;�A,=�T���j�AJ�	P�N����0=jpu,0�L{�ء����H��fx��<�Za/DÇW.��ϡ�����FQhCJˢ�q��S��:)GC>O��j�	�x��'0a���ڥ'�H ���͵��@{.��+W��_��]�r��N�8�l3庐�}�I{8���Q��1�[���U�db�*h�B�3�-*G�1�߄��,����,0HhA�=~��Q����S��tX����CY��y�V$�~�N8nW;�(���P%aHc���3q��Qߩ�D|�t�@L)_D"V/��_-���O�F�w�L;H.��6Z�"�l����n�8�0�Bہ%��}�H��|Z��f0����m��OP���y-?��~��D�n��$v�bl���X>���]�{o���&��ke��ʛ���?^�xʑ����#�+#��(��T��r��`���8�����s��%?@��{�K�>�8����5B�jS���QW���1���a�؏'�߱��=�=v̙#�=��(Q��{�Rr�)W�����ĳ*$�:(�tۑ^�!�~����}��-$�$f�������Zt�^��rG�������跣�a�FOk�҅M8o�i8��(��$F\5�8�~����6<�23���ZEE``���u�l�`>�;c�8�h�P�\�IA`�!R�
}]
t8�!SJ����k��_��d�r9�{W|��,\~����E}������NҶc�U��k���w�{��B���I�
� �+�b����8���p��g`]&��:����{�r,�2�vĲd,`�HuY�%��m��]��� ��A�;Օ�S`N�V\��22�Pη�q]��6-��~�4���#q���ѥ�u��#T%Y5�<�����ѩ7.9
󾚋;@�/H+L%�l:�5+��1c��1�'~]�9�H%��RH:5���h�
泂���w	�=*>�e��g�
J��t%�(a`�e��u6�'i�C�
i���
��кA)��d'����2������Q@���I��!��a��F�iL{�>���&��=࢑���/�`��v�C�PSǒ���u�n?<Zjg�M�����������V�0�-��7^|���S�}��]��N��9}�Y�2���n��V�;�'X�Q*`��X��X�L$�<J�s���;�`=�î���Ʀh-��࣏��Gg�b1�Z2�IT�m��W'au�Zlק�N6��Wd��G�.G��.��d�D	1xAA)�TT���d&"
;¹�-0��v�bJFd��� ќ��G`�f�+ۈ;&� �}V�{������4����+��@�����|Q�3J���I����,D�.�L{�k�d/��o�E�a��M��(+oڍ\0����C�S.����Y�F��\!)�%EAS�#�+m�����(���ˮ�QhDz�B俞+,> �g܃~�C!�G�U�l[;�S4��3����1삑X�p`uj��ǀ��%�h�+��U���f�N�� �[�wQ�����dE8j�P���Z�m!0�T,v�k_�Ppې).B�!Z�Y[�̪�X�����y眂�T́S�P.`;:��툧��vsXٴ�~_�nB�� x8�2y��6���n��B���6�]��١��������1Ó��2n��u*�l�9�SB*GG�U|n�+��E�L�$	�U�as�ihI�E[q9KC�n;A+���䱦1�� \C^�0{����llhX�҂�\y�qe���>���]Q�Q�Kؐ��"i��.]�"�̒XT(�f����&��VsW+�Q�v<0�+��+��E[��h:ׂl�
;�e��)Z�#,� �~|/-���6�X�0ӪtA�����F�^�D����Э��ր����iȕ��PLCגH�I��d��|^��
G��#c���Z����
�o���f�^�����@;j{ht.2�۾ȱ�c¥�L�J��mH��D��Z��8VI<泅"z��߷�[6
���7ÉU!����T���D6���DcLi&�"_-v'�B`�9�#RKӨ|�K���۽=b�+�v�7�9���T���*�"U���
�S��x"���FÅM�����~j��6�AP2���O�B�?yM�v?�Z�Aw �MP���3��110Zڰ�?�*�Q)�"��)4/5�Q)�b#�klx����;���v�hȣ{��0�N(�<z���s}t��Kp§VƲ��E��o��Q(�g�$Cp�B������9�)�U_���}�U��\}��8tQ)bP{ID��D����E# �t�b/4iV�I�����X��Ac56l�H?e�U_�����A�9ƛ���Խ�����o�D*4�����pp��;>[�s���ɬd��=�|��aL������Z'�F
��gغ�Q|��@�$p��t@�Z������lJ{�$�o�`P�l��P�l��'�B/:&��2-2��kCiᣳD[AFGb��o9`E��=����M]T��),��;u���g_���>�=EjbP���o��j-�w��0�[r�9�L�Q],#J��-����!����4GQ ���b	��B�RSW+�B8g�l�Z��ܹ3L3%FB�%~��i�02)�LR(%�wa۴ќ/���R2��:\TY6�n1��(}��%���kW�8�8���o�Ըtᴣ�H2���>y��e؈��2�I���O���~�[Q�4O��	q�h�)�+ތ�C�,������$�P�QsT�D$�P\\�pMPuȐV���S�9�����C5/�s�-�'R9��I��0ۨ553v3bR뛰z�cF,�{��vJ�7�XDb%������5���u"�I3T�E-ơ�_q�B٘���Js�ZE����AnڼA���:����P��#�!)�lK�hD
���ɩ�}!Zr    IDATj"��ޅak(� ���ס�<�v����F�c/!����7p��kP�ұr�؆�g�G�ye�<|�2��4B=�<������'� ��,4r���ي�Fi�JH��b��%>Q�{�LD��\C{��Nhs��n��NQ��X�r�[��1�\V�%���ka�E�b�'�iH�%��d9�>Ǎ^�sRB.���dV�#4��x�韢����	��nC�bT����Cc;�,�:c2�XS+!0QR��c���Ii�567H~��f�/"b���J�4j�E}�!2T����F�q��Q	A�sX�z��'��ٹ�lh��Z��nM?�yZ�?�������n���x����\0���#.|��y�`�d~��76i�1<T?ŧ�����X��3�C�V\,�Z�J�J֜�[�3W`Ř{� H�UIO*��Q�$HH��,A�����4ũe���:�*�'�YʑV���,v�s���p�5ȥ�F�q�/�7��I�T�7�ݧI�ք�π���0���Ȕ�"� �7�2!������	�u�X�3YqJl��V����6��L���s���Qc��7�q�K�2�48�V�4n��:���S�d�l}g4�}	��~�.�]:����?jX>��^z����{9�ҩ~;x�
1.�v�6c��?��g)Z�L�l;����u"���w����X��I�.Z,L�b�Bj�^��d&I�`�F�4a����Z����\1���Dah�G����D�����%�6�>�c��3М��J��[�y��4s�&��_�Za�%D��8��r�bK��bPI�Ee�C]���X�'?�&�y?�kN8@���0	��g��(|�7����'����"�����~=�{`%:����7�v�[8�2
5c�	�o��g�P<��M�بu����h�[x���h��v���J?���PY�#q	��Ɯ�%E�J�j�>:�.�.c/@"!�R��"��1�o�y�B�R��\/'�=���>�y���͘N�3����<�*lF���N���n�ZcU�2�A߃�*��GEf�al�S��]�*�`1A�B�)wV��$���/f࣠�R<j�J�ÒԆ�S��N���b��	�ϛ��	Җ
U|[�m��`������q��}kW����@mFów�m�a,}������Ѝ2RQ��#���PD�[? 6��C���,d�<����%��5��kV�԰��.�?��E�+�NW�X,�6-4=|��&T�7�ȁN��G�c�^]PW�UR��:	]�g�a�+o �Wo�U]�IYBF������Z%�#�Ym����kk��� ��л�~'��f���	�p8 υ�j���EMW��|T�5_��";�:�ݫ�nb���@�$��*���B���$��T�(8� �9���C�ք�����3�ǡ�:I��n��,�nC���}�p��*�}�uq�lT�����x֞=Ʋ?�FOX���/_&��je�Z	�pa��3"�׿�w���͞�Դ$l%��i��E�dS#���f���S���5����a�U��0(�+�S�j�ç[��>uN�t5�tG�yr�T,Zp�w��iQZ�q]rz�6�N���}6����񻅓1�4�ثtS����*\�pp�sp�)g��r��.؊p���a�O��6��w��
[����S�#�D�DAY����P-V|�(?��
 ��nI>U(�5p�����bOĤ&,�P�0$f4�]e�%+_�߆N�Vl�`%��9�׌������6WF*��>��^_�A��$�}�s\������|��vH>������4��G_~���
^	Y;�XD3D�����_nŃ�_�BQ1�f,�b���m.��q3N�trF-�������Λ-(���g����?ؐ���ޅ�_~���T���E�1o�$t�I#�Pq�D�lW����&_�#�}>r]C�����K0�dt�Tˡ��&�ob��M���N85}��Mn�Q%��|"�闔G0,9���(�K|���1ĵK�h�Q0e���p���H�n�H�͗C�*dZBHk�XT�_W�=t�Aa�:h��H�p��Ǣs]=r�2�ٯP�:�G��g�J|��5�q2v��n۰t�{6��~��.7�_w�FI�D�M3��<�a�5���g���y�����Y[��r�J�̽�;�Z4uȯ���~�hDl�H#)%Ib���ֺm��{pԴ�تף�^ċ7]��7�E����x�#]�@Oa��Y�u�w��_J�X}�E�oҵ[g��s���=�U�Kf-�~������{Ҍ��+��bpfE&q�
���5O��-[��E�D'����+Sb�J�a�e��l]���b|�{�y�'2Vb���f��H ��BQ�yL����	6��'�|ad`�����ա���oF������8h�I�_����ƍ�8��Eبգ�
�vP�-�P�|��>�w�0�Q+ՉC�t���j����믽�\v��m��-�_�1n�5J�V6l�#�"����<���n3mևu�E3^�w���.���$&�R�t���ԫ�����A���Î�xc�EXx�t��M�C]��G"�9��%8�ĳ��<
[�l�c��Z�J}��N�#<�[֭E�#� ��3��Vj��<��	�+��V��Vd�w�w�{�%C���B�t��;�e=�7�c6M�m�nwjPpT�>y���M^$t�/�~y��ym�J����GO���._��Z�f&Fa�=�ϡ�����"}�X�a�)��]T(��[p���PHw�֏V#������	pY:<^)�k60c�8|�4��BU،Wg_��s�a�n�%���d?�UDhW�҉W���磴�I�Z^�sn�=�;�*��I��N-.�6O=ѾG�!L�$�I�Q
)��X� nhH.�a�Q�t-:�_���q��:��FIr�\�l���Y�ɍ�E!��0!���L�72r�U\�-�e�����'� �����+(~�	����v���>��1q�Ͽ>n	���a����&�{mڀ��e|��p��W��K��b��YC�N�'N���hX�.�=s��8yW��-#�P�t�R;e.6k�P�f�2�GX|�4�����R�F=8n��3.�<�>���Kxe�0,�?��v�N�&�އ ]���N<��ǠĘ��(Q3�J�LA�(Sn�LW�����~��ʭ��3ɮ4R�@�XϬu\�C��r��%��]�N��Ft��sa���"%)*�3�JDۃ�?;�,�>��g�dt����m��.nC����'~8z��=�ipI�5�Z*4�4���M|�?����Q*�15���i���<��'8a�Ll�jѼ�cl�ۃ�9f(���S����G���|ڈ{ߏc'^�u��m��6�_�����W���^���0�;������(d5/�5WL��{�iS�̇�a�Rȕ"\y�:��{�-A5"�J4\y���K�xv˚�Z��m�6��P��˔�Th,,ɧ.#�$)��)ZN2"߳��+��
nYVa:*��4��_�(xe2��]jhȗ����ݭ����t|�<�]<v�e��l��۱a����c�;o�h5v'5A�YB�¯���3u�ƈ�(T�5o����/l>`nLшJ��{�V5fp������BԼ	o, h�8���
�2`UZ=z����m�[�_��f.����ZD����W�=c:|�l�PҪ����3t�غ8�Bd�
Bt*7��\4Y�$�F`š$�J4�����.��G� jvg�3�f�r'K��L��<�"�4;+�)n��?�5<RY[��v7����5,]0��=NW���������Ġ	J�^&8�q(��P���?����,� �˴�NJ $,�z
�Z�����Z^�]#5|F/������k��B��b��.e���]�^N~����2uxF
MZ�T-�ЭC嵫�5}��r�8t����G&�$qR03u��Z(�5p� �\�ݨ��ƘGY	X�|BW��=�X�rv(�L&����Z��bq���L
㲶����cIӦăI����a,�n���Jsg5��R�� mZ������%N�a���m�7������?z֥��=>x�]j�J�P)V+ ��z�$��5$Q�y�� ����N6ZaR����
�/!��?�S�%�)Z��$�/�B��n�(�l=]*
��tRI]G�L�͗$�Ϧ�'w{��1E,C,Sig�Q�Z>|*7�z��H�$ϰ�h�[BZg>	P�N�B��������\�<ߚ�;�bi�x��}$������?��vJ������l�ǃ5zv�2��)�ѫ��)��B�h3�q[�1��ѳFL�����!1�x���u�,Q�T:��H���2�ZYk0����"�mnCJ�0*+v|��\��i��Ȯg I$���d��'�?G�ȫ�	��l�0�x
(D�{.��O�0� 6o���J>�˼Df3>0���h���|�L����K��tV�	D4��PG�v�4ĄuM[��wx�7�F	�
��l�K>���x��sQSi6�dh�Y脍b+�_1dԨ����;�Y�c�d�Q�[�j��6����6�%�i2I���>X���y�]J[�P���q:L�Z����BX)n)�n�˓��SKOk���؅GZ-�/c|�|/�&O�f������\ض	�+��<���m�ek�^��h������j���吧�x�>ue��}ʿ4]YT	�21�c���'^��_٭a�}�#g��<���x�3���5�a��C0c�.��.<�n����)W@d�ҭ�}urwuch�,�q�Γ��U�R�N����=Rv_=q�K�X�R�`,'�a��
����t�e��'�g�Zm|@��fg	� =m��c4���z7�C�b��7%���6e��R0p�$��SQX�+r�R˴�|^�x��7_q☑C_ޭa����3FM���6F���-jq����<{VTF�U���&|�H*a~�'�8�e,�[&�q,��-����8F�!-��	W�Q#���"��ƀ��7QCU��)i�/�I�
x�~�s:�*oD�zH���?�c�����<��3�ﬅNT�����P��7[�<hV�
Me�����Z\��E�b����|6/[8�ї���=�#?5e�/�j�"�a�mM��r�FP�4�ӷ�C�k@�cI^ �c�ſ��������?���RS��h�x$�Lx�\ghе3IV�Q�;D�h1&bw`�=�1M=8���֎���o�m��""����@I�3'#��.�� ���vu�c1<��lGr�b� ��ѱ��p�K���!{3�2�7�+	��BI�1b��-[8��=�RQ������d_�Ca�f?����x��@����m�k�3�J�.����s *��{��VW���{�L�N	������x_>V��P֫��G��ʆeo����R񝯖������\8Z�oy����,r0�&�RA�mNUʛ	��cP��=����8�(J%��f5M1�7W���Ο{��R	1�1�'Ti�&��r8b��Cy�����,���*!P�,F�W@my^�c-�=��0�+��R�mj،��M�&O^e���a5�C��5S�'�T�?�\d�U(�K0���،�/���D)�/�����|�7^!�iIN�XLOb���n X{�� �I �A/lDgm+�����=������ҵ��0�/b�[����,�vVD�c����������{$��'ޗ�O�>Co��ϡ0m��C'�u�-�j���0���%m���w[C؆#WV��8�d�E�]dc՝�p���ثc��^� L�����T�|�t���2�F��'(c�c�<b��8z�5�g����!й�A�+&�1��b	l��3)W�򐽗�߈��F<s�L���Km���`��X����`R,�*���롇��F���;>r:�:�ރ�/�OY���%�jh1��;X�%��b���F������=��Q��������0BW��$�e�ni�q�=w"�u�W#h�{7P\>b�T4��Wk�P�� �7�6u���:�z!o�IBC҈S��\5��H|�Y�Ӵ�����0d�	�]���ų0n��8f`/^I��P�X8w>V����D�����a�3X�a�~ElT�qg�!L�@�h^�}\~��i'��0*�mhp�f[ҍ�i���7���5����a��I�֩C�W�E%��KF�P�9�N�����u���p264E�b��8b̵�W퍂Q�*$��\��R�������q��&���M!�`v�C�h3�_2cƟ�c�F�g#O���ebѼ�X��[r�bt����܇|DF�N 5���GLG�����`i���=��%܄�w��0dEqʜ'��1�&�0D��E���T�(,�3];w��^K��p���O��N���=dȉ�B	�����3�.�c���Y�����z�l�1�I�]�<ŗ5A���v�n����DegK(�d7�&�ml����7b�*���T��[��v��y�Gv%����2��l��X��s���1i���dInO���<�J����U���ѹs�j���	�K1BF{^C�R�95e��,��]�|�^(Y�`�Q��	A`�K*1-���~��8W%���zzVP����%31n�98f`_�0�"<±M,�{V�Z�89��'�{�=��c؈��}����,�P2
s���u�s(I<F�c�}}k���h�a��C	�1�4��蓙kT>���Fa�܉�Թ{�����/�a�㹫��x���t��]�u��rfM^��hJ��	�gF�d��c:"����� {Z��C�a�2�����lØ0�,;��pl�*��[�Pr�\�JA[ƞ��#>$a���
�_(�q=�8�������+���y���2rҼ?��0T��鞮sa9�,K)"������F`��ɨ��M<���ɰ)�#GUB	�4�{����O��KGHKPTL>s�O^�c/��l/�*��M�����KbY	��'&�_�0,;�\-;(���9�_<��� ��%M)��0eo���j�W�{��|.��JP��a#����ֆa��v{�6Ɗ�;y���j�a�a�^=�1T��:�1�\��2̝;]:u�K�{��#b�h�+WUɨxs��Æf�'-��/��L/A��&��$S@B$�e�QC��;��v�-ư��w� H�)2�j�~�B��w��/����$��m,�V�z'|U�=��r5f
����/��.إa�Y��QUI�p3V�qyn���C�8D��G�9b�ܧ�b��P���Y$WFd6�mF��1��l:�q:�Lnd���0��F��tT<���Y'�de�7��s�i8��d�@� �|��}L��z�8��ӽШU#G!�te�k�#LH�T�S�J8�a�T6���vu}��q'�9���L&��،��zl�3fa��q��_���EQ9�O�馛��悔ޝR(����~�1�8�7l�5t�$t?�:�z&FW*��8�!��k���RU$��p�%��vø���O9yޟ�j:�N@.��%�!�/n��gxeŵ����9EN�"L8p�Uh�7�?<�1Zݡ�^E�E�
A�AK�n��à��(,���	��&V��o8�G���(�(h\Z,�{5z�$�P���k��P�ʎ��ŋ)#QH+5ZQ�$��8�r#:�#8�6�����e@o�ۧ^PhZ��]�^�����o���JV~�μ&O�����=G �+W(��?��ngM��� ��p]�7$���{�kk�1�m���؉�L�����$� �M�8V��	�x��o��A�l����2'�B(�Co}:c�
�o�M��\����gJ��􀓿-]��⺃	�
ƺj�1QT����I�P#���![�c���H`}
�����l՛aI �Qqh�z�    IDAT���_��@�d�-\�����m~�GT���.D�Yu�Bz[��T[ �:�u��0k���|$�&���0�$�4/_4��=��v���q@�d�+`��}#ȣC*@��`��HBƜ���t��bHJevo�sۊM���Bj��mo���Dx�03Uȗ�l��I�0��I�������A'���+��Z��L����U�CgF���/�1#�V�^!}�+P��x�3�*q�2�
~��c�^��A��Q$a��g	L��6�hv&n��}XE+�Ð�Wo"M�,�f���<�F"x��͟�,�ui�E)��ga!�D���#��,7�\��!�/�LjP�CGI))<]�O!?�0��&1 ������)gU���9�{镴r+���*A�:4M�\�҈i�g�[H�j�c|��j�ؾ��g�,����6?=!#W��Ie�FI<I��\i�q�;k�|��}��F�rAC�)� Nt�Q#Ur,ͤ��y��l��(��%7���![�fkP���?K�6�} �t�pG���2'�݌�܎������??	I�)����"�|aK�Q��G�c;!�8A�DȈ6;�b�x���R�>����+8"��{��q+v����x�$4
�z�X��uJm�6@������0ڄ�jWUR1{Ob�Z�Qw��{&�+�2d�c��I���Q.Tx���(V�� ?R	�Z�yTF�����.�X�����_p����l|4��7�#Ij�O;i�I�T1�ib�\�?5*{�X��%����0	K���(r΂iā��(�[b;3�؃%�n4.A��Z��\v�lE�m0�ۨ0���+�xbl�c(�yk��&�h_�+nq��i��#n)#����f�Ҫ%��!��̡x�=�:�L�S����Gy �V�^*���X̋k%��l�k�ZO��c=*wGMg����Crbe�!�8�I�+�Y�0i�'����sɼDȢ��Ğ�>1lz	~�xO��U��k�O�?!k���%��Da ^)`4y��z��%$w��hLP�x����7Oo�-q��J�t�+Hnl�	�I����O�ѿH-�<�J�8�����[��s���-�S~�1���l9^Ib���mx���-�ɱXFȄQ���v9ȚG쩨%ƽ?R�
���q�{'�xw�bj�4}al��"U����h|��]�֯����cH����ю骂ޫ�͆��bɆ$�'#n�8����$i����\kI�*�H������_�Ժ�3$V�5�0�¸�&�^�k8DV��	h4�c�v%�xr���Q8��p�̟a�+y�R��^J����7Y�ja:n�����!���M����r��GM�G|�$�k���oF{��u�j��Ee�-E� �zc���B0�`�Eۑ}ng�۟���M$y�� �a�?B���a�aҕ���G��� �Cl��&qd퉇��J��1q��i��ai�����~\�R�Dr8Z_�T9�G%{}�o��j �S���{�>Lؾ%�r��x�v ��tQ����j�I=%� C69 |H���sw������#_�8f2]�ױBH�[�Z�&�=.��	��!���7��"Yud���?�*�/���]hh�5�RQ8�T*\1�������D�5)��sԿT�Ί-��Q��ѹ�����i���%� Kj�4��%=^DR��� �Klb:�|���x�<I�J�h�{��H�2C��[��S1h��e�P��k@]M��7�(l�WjĖmM��J�lMg�k:	�g!�����0"�?[]]YH�]=$Uٴb⑊C}�@�Z!�X�������
ٶ}v����[�ў����D�/u3x
�z��E���!���FO�|�r��b-yF[�dL/�=���Q���lpe�r��|Ԛ6�}�W>|���V:=�b���PW��|�lY��"��s �p:����EIKAKנ�(p�>�5�@k�QM҇V}�=>�V_�ŃQ����`_��a���}G���2��˜C@0��|+�B�$S��M0��	>���J�RNO뤬-��g�B�LF#iH��뜩�ѻS5>~�oX� o�N�C�9��?2�(����T��o���<�L�|*`T��w�G�����ed����2wQ��˅�(UM���V���*��dUA	ͨ܄��%�b�P@�<�����ٴ��5�$g��)�+w�U����ln�)UwT>/G��IC�|�q���m�z
��ADb��ql�?��*-,�n8�����r�=��A/�?������Ko��OEV��hI`��#n�y�o��\���y	g�v.��0q��[���g`ejĚ*�q�h��jy�Ʉ6A�WtYHRO]��=(
�?�+Ir��*+I�e�̕�Lg�/���wa)�9�P�V���/.��'P���z�s�L�, �ƢIĮ���� r|R�U���^�f�\�V�JbFd�7�ؖN0INI*�5�%��n	�TVi#��>���/�A�{��A�^��|�����8J*���x�u��w�Mx��_��3�g�ES�F٠�ԅz�Xצ��LZh��*7��L̻U���DtԷ�[��͊m�u� s��?�.S�(f ������Yp�(e�~��$6%gUj��G�l��앴u���7Q��B�D����	�1�����q�_�~{w�
#Ij �8VUa�B|�������Kg!_u0rf�����_�� w�L�M9!ZT�_:��D���t�6���3p�����?�S@A�n
��KQ�����c��]�#�&��Il�\ ���ab������p�����썜Ü�BT,�4�� i���B"q&$ơ2 �2��HS��o~���z��z1��W�荰�֌4��`�y����t���+f.�~ρֽ?"�k�1H�Cq������q�=YjnSK�=9F�㎉X2
:v�(�x�iȌ�;���ΤMB��0k�|{��(��-A*��ܹaȅ�E<�� �����b���~�c�d�_.��tQ�	��U|�e�Ðe|�ylj`�S ��H�	�-Ǐ��)�6��}�L�N�)���mt��*aAP��(��sE�.�QS��m�]3V��!Io��~G+,�y��T-�����a�x����w�1Sh����v���6�q���׈I�~�6�N�<�mKf�W�[#5�	���J薘`q&@��isp�%W��?Mz�"\߅ǐ��������۫�����_݃O��A�=�8,�,�>R�'�$7R{a��#�SÓ�2��m�p��9_�*{�t.���vE�PVd�%�?(+��D4QRV���e;C�� j^��<��*��x!�8pX~$�y�XK�Ca�:���F��}4W<Fblʩ�u`��6������NB�q9	�j9s��@o��L-�{
���l�b��K���>�2Y�yD����qV�9���c8���Qs�D��hLt�<aq���0�fv�K�{%1U(O������б8�F�kz��;�H�J�TX�e)Q)x�,qE�<�����̒i�l�0֯�0�����.���Tʉ
�����𑳰߰���u���a���ѦPr�̾n��o?�I��� U�lI,�t���\u�m8���1�r��̮B	2��rR6B7��Q�������{�ۯ/�(�u\��\�����4�*M6��(�"Xr��u��1@fç܀��y�8l���,n�U��T�Y�HJ,)�w�Ie��ft
?�P2��0�O��&��S���)�:m[�����=�&�z�TӐ�_B �r�Ģ��S�Ю�+7�[�ᔓ���C����7Pg����&+_x���	��`l�2�T��0X	��rK�2<8����W���'7@��,�=ߓ0��_@�i��f�3[��q�R�_�#���z���[ߌ��"��Z��\K��e�Qs�Ua��a$ɧ��Y6P���Uۀ�,��C�; ]�j,E�O�!S]+B����1��_��E���F1Jn����F���Sy�Sǎ� �5-�(���i��
��f�N9Jw�c����CGLG�n����W%1�"˴z� �ӗ����!,}("�"qMv?�u��P�Jܔ�&Y�.RQE [�Im�F.q�X����<#�����G��'�1�J�T�'�妆p�;�p�1����UF\�)Ɩ7��7b��a���0�PE�43�|��!o�*��e4�������a�=PH�:@�!�_���ʫ�[�y��)�^[^v����&iZ��%�T��(Wc�3;�Aя�1چ�K�`@]�~��iP`�/5�Pq]�S�'��G�N����W�Jꪥ靌��G���[~���?���3�e���mT������d+�&&9Cd�&����ܭ�����!����o������,2��`��iZ	f���9Wi��%9��~��_�EU�e�%mB��}��?9i�Ͽªą�N����j�ap4E"�,t��`�/�䳇�ic+({�M���b�Hش8�-���dd�IL�֪z\T�4��o��������a�ᆊ[���2�ފ"�H�iőE�7	��7�9�R��V�4�?j�a�kS����14H�[p}�:d�?�'?�+������:eɾ�<IO�j�f���_�lF,�IB��k$i\k��˯��y�>�n|�Պx�n�BtO��+ K����&�G�v�fcG����X��4[�ߘ=���\�����E�2np%-��z���rو�^m}nw���� ��Ð:ݴ��`�l��>O,�	�;���I
�x��vx�U٨"_M��yղt˸[��Tǵ2���~��50�3�^�Ԑ"�Ꮠ@6�uGu8��jng��Ƕ�"Z��a��0�bzU�#+�j�P�/iKc��+��#3���=r���s�
C���l˫�D+�|H1�[�����n���Gc���W9��1�V=�u�\W�h�]��n
��P�\��X��/}�����C���Iw�!�C؄�%/��NƆ�ȑ�Q����+���!�ǿ��[����a4-[8��ї\��<�#珘4����0��Z�.�d�2����F��a������.?�/=Oe�0 �yp�G��8�`I��ۣW�mC��r�/n�Wf+��x
�?gMX��A��+�r���sD�p�:�Q&�9CSp�v��4�� �M#w����WV��/��6z���7O�Ƙ��ڭa�}����<�_�aD�ZG��-�v�����f6��o���ϱ�+`�]�d�Z&�n<�2)�^��*Q�&NB���H]���O��VǼ�Kqǯ^�ާO�'�j����/_����<M�`�(i��cH�о䳨A{0fh���?k�>z��)s~�V��4X���p^)�
�9E�����1�����ֽ{�Mm��}MҢnG��&Q�t��X
l�� ƥa8�٩m�H��6����Ŧ��Dyh��R�D=t[2���QU�s[r�{�8U�+��@��媅����A��4����C�Ƚ��%�S�*Q�A����
�����'x��Yx����l{�9=&�� �l��{k���Dmߣd���웴�iKF��n5lT�w�s(���헷�c����ᣦ̽�m�����M6V��i�BP�����;�G������o��x$wi$��ÃκL��>e���,9�⍕�t�yʓ�G���-˔�J+�����r5~�ԣ�α��� K�jx&s3�+Q	�a�Vj�$��S���;��:<Ɋ�����}�ހ��	������ݐ��M�jn���H��՚QW��,����z'5Pn�TO\�;J4��ka��n֜}���5U�W�}�7�]8]eK\�z���a�(�勧}�ҋ/X��P���#'Ϲ�-�����DÐ-3f|&4K�Ϸ��Ƨk^�|�����X��r��ϛ�a�Ð�;��Q�Tqf	�o� ���v�� Ҝ��O�W��7?^�,��5ٕ����H�u��Đ��7������rr{&I�QW/�}\���s���Ƀ$S���-�TrT���
!��(7�R�6t�>�SKf⅗�/��Z�Y��0"2*aek��{��Y3Q���C�J�b��!�S1S������\y����ڔc��0����`�.�*ӸBHè-|�ՋG���b٪�z�soCS�Y�q�z���o�3�^,au��Qml�y��t�Xh{����T,9Q��]�J���t²ZLՠ�i+:�BT����f�/�_�G�2KpP�c�	���G�1z����W	�����Z���ۊ~}���.�N��2��9��ٚ� �S�D�V�!�C3`�[ѱ�!^�g6�!��5a�|�x+np��#�$�d_�P���OB�3f���a���V���=ޤ(�O�Z��T���e"DI'B]�#��e�؈����B�Th�a���������/���� l
�����ceR�Ls�!��-"]���et��	����Q~�Y������j��: 5CH>Bq�
dGa˓W�*�/D�� �H�N�JRړ�=����3�l	2��!j�D��8�op��*�@���FM��ن?�t9�"˸(�}|��L
�|c�Ks���g�B�ϑ�.׸-�V&x��R�hO���,���2s�'+/����:�Z<�&����K��,)S��GU��l��Tl��<�F~��#�ڧd.�1NL���������SK�3���F���c8吽���"<Q�Z��
����Pf!RnqoCT�X��/gl'{ �����w����q�������1&�b(~�,��Pq~{sk
gz>JhTkE�4���V\�	��1��E� ꔃP#q��b���Y��9��Q�x��Ͽ�^�Ǥ�VL�~�b�I�<�%�����^à��*�(q���,���닆a�3q�atw6��Z&.�[�a)/�O�Ic�W_��OE��`4���g�aPK��t��R���Mq�|3�j��{y����?�+w/�/<�/���g>{�Vӱ$�y���J
 j���Kzs�҇0�y8f�upS]QD5�	�m	�!ق�y��D����Q�����fb���qD��Đ�+���(K�Ͳ8�[:硗LG���
�g  XՈ���0V��M��6b�ڒ|��ÈҒ ꑇN�:���"\5c����2�l8i�\�@ΦӢqFؘ�0sҍ8l��(���?%�Z��� �� S-g�<�n�kR+,*��N	G��1���Y��[��G���	�(R*�H�cW[����\5����W�u`ظk���?ǠS`v�m��HO�H|��4�H�����������:� Kⅻ����g��=��q�� _R6:�Ӗ
9X)�G�Dߋo��c |�D0�����	o�R��*�l�a�ݎ>���TʄdV4hiA*Q��s�+]�i���!��E��B l8���{�42Ӭ����+P�P�b>c�Sº��wPnB~u[})�z&�&��CD�Y�&X����ۯ��?�í+c���@$��ċ(�:�PP���~Ç�:��#�Uݱ>�ê� b}��x�����"nC�e��<^h80�[�����2�ǜ�c�)�O��f�N5B.NŬB4,'e���	�N���X�kx�����H��ٽa�Rs�]f���!Z�:��8�'U��y#q�vXF'�_<
�ǝ���<����OJfˠ�L!W��W56t�C�,�����[���V�|4�q�3�D&�Ze�N�@JREt�����+����2#'\��:�uA�\[��:��/���}�u\q�B`�����#N��&_�Nu�rQ���0����h��C�dJ������e�L��1p?�,�Ejy?R���pH�����G�B��C�1PV�Rg�$�D�uC�-I��-����&�Xq�CGM��`[BI��j�ֆ�	ʨ�c��1�t��8f� ��BK�p��zI���L����s�V�~��<|��}���ʴl�'$�����Q��/���c��*��	��6`�'�b���QX������_��i+���y�>�Px8�>��C���5hU��T�@L�    IDATv��/j[�|YÐ�'ӗR�ݍx�q���#���n�t��?�I�R�%�w���Y���л��KY5v�cm�|2�n��ضy�{�o�-�6@e��j��*܌�n�p�@�Iy5�F��җ�q�&���b�������y�NZ����M�v�N���d�@�i1ތ�����(5"��r���I+�a�6��W*ɺa�_
������ �,�"85]��)4�
"����YxLwiINQ�!�6�e��uQ���f���f��yU��'���
b��oy�3�j��+<�I�#�DS�uh�-ø����9y��m�I#�$�$�gV�#P��6j-]䤂����#���k:�.қ����0�ڽ��7kD��8M���1��*E�|~���.I�uN�q5���eW���Dl*�(-�2[�wcU�2�l;KXI�H�6f*��\�L鴃b!�T�VDg�b�Ȏ4K�)x�D�7 y�������G��v^A���0SҊ�����Q���l����Ɗ͒����7���8a�x��?z�Isi�aHqse�9�/]I��V/�aK�wQv}�p�TZ��n�Uf��e����7��s)�M^�@�	U+\���0ĿDj��xϗ)-x�Z�a�@x�Iƚ�����2%"|#�J�*��jh*9qY�����%�({�+.SC(�)�B"��i������^]�2T�`"���҆�D_����0�4%�,J�}��P����/H��F������E��l���\*�o\�p�=�1����Dn`+* �x%�)���[�JV��(���I-#�c�z�W-%��7�+aS�J@��@�`�l�/��YJ\���c�8�Ed�iY�XM�1����lPF�hq]�G7
�!��s�َ��[P�'�<d3�_c��-��n�3��=��T]VAɲ��	˟���YK6��G(�x��j�RN��H��*�P��(��0V���٣��{�����"�3,)����Q��R�,d�Q�U�M+Q+Hq	�j�t�|p�4t�!�����K�-���*�)T�.%���ϝ<��|��z�ghJc]QI2�(�6��&�@,+��Mtۅ��W'7�"6a�)�*'o����s�PQ����w��~.{8�c�ՠt�(OxL���*I���>��-9���B��)U򲖮g�c��0��<��6 uڮ�|�����yLɖᯠ<]�Cn %���{�*�bY����IOD*'5�J����I�9�O���I
���~�����8�I�TU�A�'��.zn����JA��Ϲ���8�5uSI>p_�]NI�ZA�c2:E���U6��A��[11q'��/:|�ra��Y�}YT���vF	;�dُ�eΐ�0�ސLSe�[�S�>�T�J�/���=��ۃ.��$TJ�"P8Q-���"5�u2�(�p]��Д˫�C�k��#�
!��Qln�ϕ8 �R���U�r�I}c)���u't��l�5!���GVg�Z:V�_DZK����;#W�s�0*
קw��`%
�+wI�It�p�M��JjE'�	p�����P��KlYS�_��JO�PjY�đ!��,�[U�7׀�AI1Ű^P�l��Q��N#�z�����qJ���W|��A�("��bI�%���dm���TTjB�Y��aC`��pR5ꁺEX��M�$E������VXB�a�{�Fs���	���<)���q_Z��Q�b�,-M��*�JY�dYF^N��ٍ�A�.��r	�Cɍ&ľ��d�#>������_B�LŇC-.�������+�oǥ� ��j���-t���lM5�%5��$��D�v)�3�BP'�7cl+�<�n I�%�r�H��������D�c!�J�c��X� D���*�8��\��ݺ�Cڑ!N�4:o�/b��*E�y(�s�i*GH�����|^Z	ZA<�DV+N�K�	�S\��+�2]�d��=w�l��x^#,ǂg����&�i��\��|N
�b���t�A)�jH-V�|G�%a��'�����Z:h��fb(���$r6+��0@���s#hl����,XF���Q���"��(A�oy���k{��C��*}S��ɤ��,&�erZ;B���6C3#)b"�M9�BH�g�34�]��r*�R2m��!� ��u�䉬�,j���؉T@6A.�T��G(����t��ư#zL�y�"�� n䢙���� �T-rVHY)��y���#��p�ɕD����p�+8_ �+�'*[�Ԭ1|��,Sl'R<;L��������\��Y(�Bx�S�\�衐;��P,Y����0ڷp�2k�!koE���L`*3-�F�F9����7���	U�#d�.̭nIT!&#���pɱ)�<ܮʺi�2Bu�٢���"���	�R)�~lp	P,�^��Z�\>&�
q����p#���b�ơ�eSY���c��)4E1�t�B�P��R7�Ur��*�&هm[s�4�L#Dѣa8r8��Ӏjzٲ���PE"�#�@���K�BB}i�E�?�&���P�&�ؕ�X�p�W��P7 ���F������&��0��'aӨ��oF��	���i�:��YzU��CN�#t���e��\C���
��ѳX�M�Ig�d��r&2`���.�ha��e갵"
�m��nظU��u���T�[���5Ǉ����a�a���(����1�����Q<�L�Z���zҠl�% a�C�ə�B�sa��<�xՖ���|��W�P(QۡNr(�����\tѣ�^H�r��l]�X[_�2����پ���|*:B���b�Qx"��͓��B�ۄ���ǡ�Bm�Z�������+��ߗ��G(4n·���y��?�U.oP3��zϬ^O�@��p��4��طe�ې��r���W=�[��;��ף�Cg�|�x�w�A��M]R.z�쁗�[����c�늌��J���{���O�0�����*ui�������L�]Y���]�RN�����s͠���c��zⵕ���ǀ��q��A��^��	��� �WF��0��1x`?4or��k�fK[K��/ۣ�ve(��1M;i��h흮�
��*�4�f��_@��Ƀ:�_o�<�V�
|��s��n�� �Y�a�]t�i�k�:|��'0�4�[?��}7\�����!���%Nxc}�B�湗�i<�*�IT�KRjVa�bȡ}1qTo��%��Qk��o�����⋿���	=�6�TzX{�!�p�/q�Q�b�y=�֫e��� �����;؝��h0P�\��ȕ!"jϬ��pr������G3�E��
Qӧ9�����{�O1�GCq�`/�=Ė���l�r˳���p���!p��/oA���e���^�V"����Si�k�1�i��3NڳRs;�:I��ت�Oվ�����}�&e"�o�ms��+n~~�%�Aˮ=/<�1~���y�yx�X��x�ݷ�ǣ�OŲe/���`�Kw����7�?��&�u�,�Q�A�.�uK03���������O���4�P�fk��z�zv��o�}�æ='?�� �&���&�C���ptg�x����p�����b՛y���ߠ��P�!ym���zbA�"M덫���s0e΋�|�m�+��߽Z��F��� ��|�࡬G��s����Q_���?���A)@�J�>[�T�!�7c��Y�}�y�hm[;@Lڃ��a�a(JQ<>����5�,7c`�z\x� �h��t�B���ۀ)�5�t0k�Op弋���>��~�Щ�߼?�w��7�ޔHےK��-f��t�s�˿�՛�j$��������]0��>�A�k?l+z�ׄ*�N�����o��Go�����ƕW��{�1v�i�h�8��#q�{bܔ���v(P��C��o���������0�(����t���Ȕ�a��`d��Kđ}�a⸓1z�C8��� �ࣿz
MZ/�4�L��'��ϋ��{��#��R���Y�w����� U�EDε�+��b���G��`����� <����۶YI���Y�ڔJ�*�GCC�p�)��ē:�򫟄�aXv=����N�|����Y+p�Q��ck�v�68���#�����^�S�d4~��!X�6��~�
�N7ԊDX���Ȱ
�n�)͍ͮ�p�1�����p�#(:�6�[ؿ�<_�z�s8x�!��I��}�r�y�x���b��0tԷ1�ʟ�SO��'�b�5� �=K����8��#pѕ�0LQ8����4�SZAHIM�oވ>=:b¨��r�
�6T&���ߏ��Fc��?}���3�����em �~7�$̜r/>3{!��yW��,Æ�!#����c4ߵ`�ɗ���n=���>r��)s�i�a(�E����I����3~	��	��Maܘ�8��G����M�*�0컇�G�,��	L��,<�Л����ix�mx`��~��V��-�p�����5�g/�OwGFKJ2͊��`�-s��T��{�`�E=1}��0;tG��ѷC��c��ᓟD���q�=qͬп�>�1���ﮧp�ȓ1lگ��O��N��u7��:[7�ǹ������a3�v_�Q;�Twdc�8� ��G@=ִ-�qż�q�-´I�`�m�����̪�Z����93��PFA�!16�r��(j�I~#�Ad�� )6�WQA�A��$�2 خb	2���9gN��f�ooa�k�y<O���o�o���U�������ˮ�h�_��폂�C���hށUs/������� ,�#P�H"Ef�^R�j��|�;��,
=4�_'�|��lF5��&^��lĶ5�u�ނYS���;_⩗_�-�]���X���֡.�桤���؉��(�ɜ1���h㞧6�t�f��D�T�7�@�9b*sp߄JQ����s���*6�F$�Y�%[8nZ��8	���7O{��è���
\��Ӟƙ��E��;`���?�d465`�X���Wo�)d���Ty�H����$R�Ԝ<�&����8��/ ��|��qr�1�:|!�pg$lb!���fa�Ⱦ��ۘ��i4
:uA}���i����w�+Y5��T���dT&$;I�q��ۋ/����w�植�N��l��]9�3z�聑����{@m��~��x�=��e/B���j�6�\$����/C	���5@���WS�:�.+M�.��^��/���kZ�9�ǅ��":�U�:�L��7���=�`~'��v���D�;�9�~֯q]���C aǝl�R�c �,����&�M�g�'�OC�)1�@N�[��_����_�� ���8n�Gu������/�@���]w\�ʝ��-@^PCYɚ��G,�h[��A�h�b������?���x�<J��F�����>5�t&o7�P,��%e"VW�ӎ;'��S�s�lM��w߆�`j9��4qF��(������a��g~->(V
�W���슛H��P:�+�Ӊ��M=I�yU�����il7"!�\t�! Yc`��j|�����'�_|�vN�]���rQTt$_�ݏ��~�Aꯨ>���d{�
�
EE��A�� %>oBN���\��t����2�G�>��O?a�?I�L�`%�����X��Zl���d�p'��D��g$-��u[�O�.֌PN������V��c��C�0���=sU)Ȑ�=��a#�#��S7�7Z�P��H.o����Ò0R-h'�nG�D
��|dH�D�3
�$d��*�����,�]e���P�ށi���g"9~�$�k�!H��$� O�Y��h���:k2�0-)�x��.|2R��P��Ɍ�K�$�3$�C�ɢHc�g/�t$`D���#�!��`�a�`F"[63�8`��z:Ú(�t>Ӏ�hJ�hױ�Ob-[��Z\͖���,�WXۢ��j@E'������I,����S�1�%f�4$�..�O� KBʰ�H�Y��:dL��.)YZ������=A�I��_h����Q$�Is�n�M���1H���a�SU0�Լ�?�d�ivj�z���_VGtU�\�J8Sj�;
�J�+����룣��b�ϝ���$��}�D"P�xV�	^�t�NӤ_J�K�=�ᙓ.1��~��č��L�#E�J�%�_P\�I�E�uN�3`mr�9V��S��G �hD�~^i�����iK�(E\�J|�t��n=��A�Fe�!�q�Rw�J1D�#{�l�4���N��7��*�ihhDT5� �GR�<$�s�1�p�Ej��bP��$b!��4!�#��ޑ���Sy�&��V~��AR��X:}!�u/DP�{���1�5����o����͒2T��Fm!��4L�:�&�i@*�+t)H1UN	�)�����P;:'Ľ��� �cW4fd�dd.���E�r���
� ���A��X�6��,�6Gy"�VEgԃ�y�Ds-l"f�izNw(�����<�"��$�!��7�0�X���Cد ������)��Mք���@���}P5���BGSFB�{o4e迉��f|��+p��/�q�o���q@�X�xŐ!��~��u���<ڣ&b>K�M�r�B�I2����&Rk�L�KuDVO%qŁx�|�D���PvҁBH�KLx�� ���[f�F�IO h5��s�t����"<j6����oݠ
�C9��~�<xD�<��A����뽨�	(��P�l&Q�y=��z�A�
�����T>�z<*)�O�r��i� �
���#1�I�>��4�KV-wׂ���]�8��/�:�;_Bp>��f`��AX����hx���EZɛ�"�[�E��ۣ- a;�G���+��I�?�I�a,���&�@��rX|:�:7㍹� f=��`n$�H�o����Ť��Fd@m��Jq�)��QKF�ʢ-�w�s/n�!�(��D�R��jT���J���Sg<�rIz󎞡��AHw�^�g#�+�e��&�q?�W�+1֔��E�7�c2��G�n�@a�
}t�/q7L����B��F����z�|�r��@��:�o*���/�Y��v�/�NG��)���v�N��=Q:�UR�%oefP�Ϡ�ڃWg�dvv�}#�-qc9�<�n��K�N���'��[�#����x��;Pc�:͊
_��M/a�ߖ��i1��j���9�����<�j�1�aĔ#��d��1�Ɣ�]�{&_rݐ���1���l�]��j�=����G
���$��AnN�H"�I�����������V�G�hE�\(�&�i�Y�G��Q����
ӟ� w���Q��4m/e�\��#�nDAf'�?8�l����+�-"F➠6W���Px�(��	;��,(�R>z?ϣ��qB5bϣ��ֲ槫Q�z)T���\2��E�m�SN��~���Dq�	�OX�z���l/�^�Ѳ`��K�J��,��~脻l�a����]���*d��i�J�Sȓh��2v�0�ټW}�{@"#�%T���$��΁T����v3)�������8��(�[[!��2��jtqvc��I�̯�'Jw[���d�Fb2J)�.��ec��� ��c8v�M�����yXWI��9zқ����j�3��l�db�Q�~�M�DW���^�}&,D����L<�����y3'^:|蠊{�%+F�������`��#���?�\�d�t�eu�[
|��1����^5���9��AWE"o4�A�:�R�T\� }�Z7�=�nԨG0��x�i @d#���$�G�N9v3
t"Z���=q`� �m��N]q^RC��G���Ǣ�	�!-�p�U���*Hd��<B�6ȨLGF;�{�il_�?P�Z��G
�b���)
t+-T=�b6�|��a1���,���<y��g�gM�lXt�ڃ��c���y�bh�����2���
6��Q����C�l��b�s  �IDATFِͪL�9̫�O����nGn��ۓ,��	c���+� �H�=�N�)G I�*�]�(���3]�`q�a�|,-C3�_a��ɀ���d .}��%�qR��ИHs
H���=��-_����j'^6��)9����<N�x�]�tw�����齿b��_Q��4���i��B$'i��k�][��̀e�^��L-DѠv�ek<}�*���0��gM�����p��qC��5���Ὕ�C�C�TB^sg��BQ������nA��5�[u/?�{��*�s=��B�"���9���$ʮ��
���l}�ށ:�I9��*�àݤ�M��J�Ŵ����x�̀�`6{�7L�������$��h2&���;����|��)9���^,A�S����a����"D�8��]�]/-㬈��4HE5��KW�b[&��(�q�5�����7,F��6Iw1-D[�.?Ʒ�h�y3�\6|h�k���ax4C%Z1u�N��o.it�g Ό�ͯ�n�}�Y�����N3f݋�Y��F���rc3�=J:����W;!)繴��+ܹ P�u\�#�k�l��x�-�U��l�d�c&��/N�	���-U������/�~�0.����EF��`(٘���<��l1F.ZP��*�~���HN��^��=�P(���pn��FL�2ŕ�d J�:i�#�X2$��ګ�������ߑ���c<�h�ء����m��
�8�:/t��n�+��v`�Q��g��(<:T����.��nhsH'���Q7s f_�d��^툤�+��jyj͕�o����i �đkVc��[������N�8}N;����"5�n��TTn�r5MX����@���c�:�^AM̮�0���[B�(Ix�����a5p�̌�2p����ɇ����ݜ60��1"���.��	}&>�_� 4��<]�	��e�fN���磋W�:����b��9=e�m�l�@P���IL����"���M�~�Hv�p�6�{/��LI�SX�2"8��<u��q��Q鈔,x@|^̊~���M��l�#Ϩ��{ou=F���ɓ�3�N�͚�A�f�uL��fl۾�5�L�.���aPZ*�ἴA���D�{A���%a�?�]lM�㟞t��#77Eg���`��񮖊�j��c,A��H7@���U~ �.�X0{��MW�Y	Sr�H��/	������p����QQ0i h��a�z�(N����F����E^$��:{i�h���PF�낳�ގ�0Zȭ�}o*g*��pD~b�a4�Q��>2�� US1f�H�:�'�3ҀM�O�6_T��j!
.��ǟ���m��6E�Dɉ����.�,�� d�a���M��B�F����9�AD�~�-��il�1��[�j��`��`*]�{�c�����h�oo�2��0�g�E-p-\�l��3�5�Ԡ��y>x��H}�(��"���3j����>�OйK�)��2"]ݼ;V- �Q��������Da~G��I9��Dݣ��Z�;�N��af����
���^����yX'��݌\���a�vL�q��ĉpꩽВLs5����4m**+w����^� �/��O�+uk!��%�'�*hH��->Z�J1�~�<����0��н�C��8�&��Q݀&L� �|u���LZ�G	���[ܶT�@G��3'�f��A�������1d���:f1��B� �"[%4�jc�H)�$2v�8���EB��x�ILA�C��+��o+�[#���m��~��ܾ��& J�R!?JXr����Q� f��#�[�`��k`�<ͮ�1����(YM�:��D�8F7�pN<�R���ɓ��˯��Ћ!��oJP���#��ʫ�z�5�����a!�ɼ~��_���|���WCs��~����׎'ۉ�1na܈�P�[���,��g�{�Z$-���j*�-�د�x`L˼{n�p��?���hђ��f�;u�b�!�!���t�N.�D��# 9̚Gmwj_s���W��p4��+��ހʏ6��:���D�@e�4f�1y9y��Q	9e��~�.|qT.k@�N�f4�"X�|����KɃ�^��8��g0:-��[K�si�L#�"��O�N�{�Yl7�<���?�v�r�(:�/�\�L�EMTQy���� 4�]i�(�L7 d7a���hx�9 ���W��W%̝>EyH;Ҏ��Ҙ~�T&���A��:f�+��˹/��5r'�����W��X��RR!`G�<<��~#�^u`������J��=��腨��9�XA�H�
zE	zBUO:k�<%w)PGn���72�US'����4�15ۑ�݁�_�q�m��|�C3|Mq�hV0�ɷ�)
����t?�$�I��a6\qxyi���T�aI�B��V-��ћ�h�4�4An�`����[;���)��ၥϠNꈌ�"��1m���w�*h+A8�#�bQ<INQ^�c#�qXB��d�64�4+�;*�D�ބ���F��iX�j�<,{�%Ȏ���g\
�[�~hQ0����b�i�6\�+y^nⲼ7Q-Ւa$�Ϟ��`����2��G��^�Z�0�����|��xR\�	�G�ܗ�Ӄ!"[p�A@��Y�rXݝ���P�8|�ǥ�uC'gBH!c+h��o6�l,[� �a�*�Ĕ�� �i*�*n��%ua�rFES�=̀^�j��'�x��_��_DpT ���3о+V��5��Ѣ��&+H�M�ׂ|}2�Z�Ȫ���b�7��N�L`!��Q��Lq�T�z9?B�j�?%cd$ah��Fg��h't҅�#�|4�R�\�LT��V��X[>�c�wЁ�K�K���Xt�臱G��L9��vQ�d��K`[����e9�V�!PR:쾴9DWd��Aq�����?V����n�nD�҆�X�h�Y_��Dn�%aD�C�0!�e'Y��[{o�%u!yo��\U�M#�To���A�b@�؃�����SKӬp"�k>m�6�H4�aPe�1�d�Z-n|�``�;:Fż,W��`��~��A<]�%�"�AH#nA�@?Y�Z\�S]�j` !��Y�7+chrr��Tj����ԓ|?���N����?��X0s�Q\��ɒ�	w,9cԃ�E���Jf�u=�bN�Ĭޔ�w��kx�"3/$��QUQ�1B�0�ڨ'��[m����%�B�ӄ��BS�x+�Ӊ̎��6��@wJ{Ncm�Hg�P뷇���!��OT@ɿ��,�X��HT�z��Ԃ�0�p� �C���1lu�Y��LC#V<j���%X��� �hT�1�n��qPA&4oBG�_��'<'�nu�j�n-8©F�6�R��:� w�V����P�v2L�B�Qj��Ϸ�4�F��ϙ���4�=;p�����9u����kR:J�!i�� ��y4�ď3� VR&W+��(7\)
⤢a^����
�=�Xa�@�"�m���q��հ:�Emb�ԋ!��R���0�.tq!�(�%�����ꋄ�th�@q^�$��MBK7C�P�/�+��?2a�
2@�.�uT2E�)��OZ�:�G"�h���O�.���,���	K��Q���I�Ȯ�߲A��NG�zo;��G#)E����� 	��j$b����"Ø;鬃�9�[�������s���!%^|"��>Z+�)�oA�����`0h�T�����+����l"S[����'�ev!OR��R��v��]ð�f���ԗ�!g�2�K܂�[�̟H[lK��k$���'霐�[Nz�.2qR'N��ĔBT|^�]Ng؁�0b��]�k��\��Y��(��@1�"�3�9�KA"���Y|>������F{�Ჟ+��ԃ�S,_>vJ�x���P{ �(6���H6��Ȥ{&�Q������;MX���g�|����[{�o�1�_�X��7�|���	r�׎)���G]R�GG���������X��"��@�K%=�MkIЬ"j
����}I�p$��=)}�v�|��7D��,�a����baL�����a���� E)����4�:+�I{����"n���g�Qk	�.�a�U7p�K�C�Ik�R6E�����D�d}��m���]����6h��io�)���AȖ�%�������:́h�[<��j�	[1�8���G�~�u��r@Ø����aCG�_���Upu�!�^7���&:>F@yT�8$�I���k?%@p�t���J��>���fh9[�E'� ��Uu8���p��I��Y��ɓ1��
�Ket�# �����1����Ҙ�S{��h����ѓ����θ��*B���+���D�{\�s��Һ�b^��E�Y* V�<cέR�<��dd,q9�I�ǘ���縮Q��������m����_��;������>x���_NsD�ḧhɧ��>��J�O<x�Fh��l����8���{�Et]W>�l�d�Q'��*�5ɤ��q'�0�w�ޱj��W�8�T��'a�R��;/���^�2�(��<�k�C���IP��C��q��a���85�����"[��������K;��Uv��=���Ϸ���_A��Y�耴�-��{03���8tȈl\�ڗ�;�zϞ�[2FWJ�e+u��訩�X��X��c��9cq�#Ѐt0(4�dI����:��a�u�i�C���2i=S>hH������믽�s�����G��T�u��*6�ߺh�/��gg4�j'�B�#� ʝ2�ʁ3���am�/���)SK��A�*�x�����������Vm��9�8�	��oWvq6֦5�/\�(RJ%�|����3h`tB��?�cٲe/�'��;w.B����ß������y��WJ?���Ej0�I_S��MCˆ����i��O<�L�/oQ�J��}���A%�Z��6������-����X���������yc����غm�i�T���%%W����c,_�ڱ�I�I#��+���?[�ֆQ^^�aƲ{R�K��۟�����ͩ�xm|e��\��ҷiVF�����]�x�0���RD�����0p������4���P<�h���'g��TTT������+��vdn�F�?��ڴƊ+��u���{6�yqq���Z�p�����k�0 �[RR�'��v��몪��2�O��hV��k+u]���a,)...�ƽ�o��*]-//�4�KZ�[%%%gfcs֭[W�u����cS4�Z�bŊe����p=�����ٸ���x�4�K[ƛ%%%����ُ���FO���n���0�b�0��������QB�eY"�YUU�@+��m�x�0�?�������o�ˆa��*�|cp�
\�	>?�F�=��ƮX��)]���c�_�|��0�m�16�������SQQ1����V�h4�+k�+W��K&���ceqq1-��s��kM�����8뮽�ھ�ؘ�k׎������0ލF�YɈܬ�]���0/..��{�O>י�yN+�������llNEE�����٭�h4zz6�v�Y]�/����=1p�@N_���˖-��,�W�b��|^66���bRee�V��v4=#k���뗴�Os0z(>��a����(�5��nݺ��n�z�g�e�UZZ���k�u]��3�@ �Ԁ?����(//�4��Z%�KJJ~��7f�ڵӪ���t�]����...�2���c�d���"]]�n��[�n��%kt]�x��?<=`��+~4�1�Y�Z峢�bzee�M�0�\��:g`nI����bN_��p�1�5M��CT���������0V��P�yXƲe˞�,����&�V����5�\��^Ɇn۴i��P(�m�T*�NYYY6�յ�a��y^E!��篺��~4�Ix¶��4z�r������|޲e˖�Y��DjL����Ҭ����� �G��~���k��u(>���X�d�R ��(�|��ʊalذa��͛gAZ:�&5�#G��e�ʲe�^�m�"�G\�OF���� V�\9'�J]o���ܹm�ϖ��e�Y�f͠>�����;��pgհa�f�0V�XQ��'I4k�����,���+'fk�o�sXy����Ζe��i�i���e��nݺm����ܹ�g�i�h��b�f�QG՘��w��A����$Ɇa4���U�=b�Z��6���Q%�H~��8�<�!ڃ�����92f,    IEND�B`�PK
     8p�[��/F��  ��  /   images/0c7fd013-2f4e-47d0-a46e-2d19cc1fd6f6.png�PNG

   IHDR   �  w   `�3�   	pHYs  �  ��+  �RIDATx��}��U����קd2)$@� �����T\�����b�����E,��P�� ���R$"���H�(� 	I������=��޼d2d&�̲^>a޼y����{�=�{α�o�oc�o����7������a�mlpL�X�h�2{���;��C����vuwT������M_r�G.3#�7���{r����S�ryJ:��l6���^:���4	�V%�;���+����_��W:�݇�xo��<^�̬Y�h͚5�������|�~t�Yg^~�Qx�����n�i�뮻��<����Ţy�G�iQ��8��>��J����EG}����z�U'�x�[c�[�0^xᅶK.��w/���S>t�G���_h~�c��ܹs�������2���$��r��U�VA$�ʕ+m>mg���=����}���a�4I�y�w�%�\�N8�����{  �"���ðx���Xx�]w-�߃/�˟�袋�ݒsߢ���/~����2�K�~�s睷��OAX�z�J�P:cӚ��3[M�eT��aX�:�Y�g��]�����y_Zh>��C�O���3�������y�{i�������ۿ��M��ַF�oB,�H�;�:����x͟����o^�/|�7�cKq�-B�?��>����[n���V�s�=ȶ]�
E�811�T�O�G�kS�=�����p���}��ߵ�#�M�_Yb��GWg�(֞w�9�����O[y�������%�a���i&�7����'���3�8�ܟ��'ߦ�<6;a������΃~~�y�O}����I�_���~�dSG�'�Q�t��~�_�۟�̙���t�9��KO<���7�p�?�V?�p���[�x��)8���8���E���i^s�5�~��o����1ڌc���W_�3>��;������~����W�d�!C��Ü�cvj��5Qlx�4�+Ez׻��'�x��k���eq��%�\�Cڂ�Gi�o��z���;�^���(0p�DI���QVL_��O�����f#�~`���8���{���ݱ�ڊW����5oGDF*���6zF�^W�"zz���6���S��<������k�|���?�����Rɣ�O���F+8��Htp&�f]�7,�~C�al�`�#�J柿��������AJ��S�d��XB��@N������<�0`"��R����@L����4m�1gΜ%�C�b}Bh�H��燿�c�l�6�(�_�hQ�����	��,�q�Y�����6�=���a%�f�����,�u(m��^k4�H��T��(�ʊb
����>�Z����~��G?N�q���o�Ή�MK,���Ot$Ću��j��q?&볟��������r�`y��~��w���[y ,�G����dR�_�@��,�I�:�@8I �bq����s�Y�r�i��}������?!4/��%N�f�)k(\����?8� ��9�y晃|����r�2j�h9a�t�qןq�)4oގ"B�@��⹖-?+�
i70mlݒEM	a$��d�w���ݎ>��c���_/ᏜH�a|�+_9��/���KNwB%��"�5A x�������κ�?�j�h)a<��s����{|���Z��+5�>��w�5�	b#�⍬�t�^���H@H���t��O��s��i3&�����4��$����L^��%K����vۭ5f��0.���?����B���j��ƺ%+b0Z�p��'�e2._���}�s�Y_����Q���_��'�l�$�h�����-3�[JW]}�	7�t��=�V�9E�w$���R�U)Z�`[)ל�j)a\y���$W_}��4	㩧����=�n���;f)ŴYG�)�3QA����}��ٳ��|��ߟ�{k���Yok�!o��④���Θ={6������6��ʛ�c$�����s��丆u��w���~���������`%&���"�E�'�x�Zqݖ��z�#|�p�χ��(�ٸ�b��9�ݬ�a�
�,�ŋ�e��`%o�scJ��\��w��ElOO���'''�Q�eaX��b��R܈^t�A��CصU���|;��ΫV��@<��cq�i�5[FO�����9waÆ�o!=1O7���''X�Cs�8�9s���gvn��V�X�GBo��Römѩ@�K�.ݱeץ�cƌr��`��6E�Y��&n�vp9@<��N��ݴz��Zu��^{mF��zk�D���\�r����n�k4����n���v�A	�ʳ���Y8�r�I�1���3Zu���y���	CɾM��L|D���I�ܻ����fx��&�fs�&+a ����m���B�44�u<I�8u"RxN&�����e����(��0h+�u����M���{����I<ĘDb$��y��f�ey���,:F�Di+G�y��l&�ɇ��,�Z5ZnK&hnِI�~ɢ�� ]C������G�\t8�@��c$��pQS(�b���dA��fc��|f�@�1"[[�4�AFK&�RQyE1��5���
����300H��J̈́*�O �	W�8��H�����?1<����Ds�K���2+-�}�hp����f�ϙ8��3o}c}����\=�붌0���Z�!#�-8�4���A�@8q�v�����^.��.gC���9���r��	�ɐ�$�0 =��,˥B�P�c�%�#�$
�h#��l�ha�p�+��P)�d�-�n���E��b�,�q,�cK/p�;OVrVK��q ���4�<�!�`n!��rU�pŃh'1�To�s&9��$�J����i�ò��G�iG���pY��J%l�ǜ�䵵A0�6���@�=��N�)�O���;;��B��){Z�D��g����9xUIIĕ���ʥ���N�9'��9ژt���D,�)r�J@:�E]
1�F�o ���c�Kϟo��_��;�h�5�6�`D3�T��{"�p�iӧ�?��:�5%�ϻa=�S�d��-�-�1�'@�mSM$.rȾ�����|;��|��fϞ]?��w]s���9q��xԑ�w�GN���;�8ꨣ*,\^p[�nV�8X�/��ne�F��D2�ň�Mx��t�mw�׾��2�����p���W�"	H[s`���[r Z�c���ğjU�=t�O��m7�U�t3��4>�K?vʩ���k�������~�/���}h���{�;��v?&�4+���=������7�y��@���ض#�H�8o:�pL6'W2Z�i���&k�*qpHM�G��_͋��,:v��W�.~����¯��7��v=�����8�?�o��Ƅq�㤎�5�/)�9L�n`?�tJ�D�����f�6)ul@rj�i;�/��8��aۺp�O�-�e�Ϋo�麅�v���+���/���1������ʆa�`�$u4p'�d�Ԣ�-�N�g2�|	��d���c��W	.b�h��~3�h�X��������q��_[�^��/ް�N;�:��!-�Gn�V����c`4ńZr�͇��)�dd������;�v�u?y�G?vƒ���g}�/�4o���Oc�������;bƮ�5�p�U�!�}$���%`�W�a�7w�r�/��r��xξw�}��]��/��?劯~��Oo��дz��L(��BVV�M<�8Fw+���	#����s���=������Ww���;��e��Ѭ*\��u;I8���u����%�`����1��m�}�{�\r޹�]��.�={�eW���oY������1�b���%~�@�*�?0&��1}C��'?��3>�i��?�J�6
,>v�����u�ǎ�N(����ئ�@���ͦ�~=I9��������0�/�����s�����Cl��L���PTA|�u0�ZEbu-�7%a4ڙ|�!�F�W,�0ů0�~��#�f��a��'�p��Sn���w.\x����ͯ��l֚l�)��?���%�.�a[0�:�rW�S'{M>��5y��?9s��#�Ng�V�Z��o~�۷^x�E�IE��
s��խ��shp�֪�1�6Y1��x'��~�����A����.��9p�8�1��JW�Y��c�r4��&�X�=�9F���Oj��s����s���=�<󌫘����ȡ�������<�OB���9��0��D���G�͜9s���5�;����n9s������)V3��M��F�_$DӼc3r]�b�i����}���p]�*����n{<��7�Xr�Fͮ�̥E#^7�n��[9ZKʌ%
�y�<O��bq�����M�z�u��l�o���F�VϘ��dN��m��ZB9E�1Ls�V�PEl�g��9�m��.L,@�nR�'��ko�w�̖��d�$Y��N��Y�2�2��);_�1Fw�01���Z�㴮�ũ���e˖e�I��~�'�R6��Ea�:�C��δS�7��sX�R)�OW�ߣ��[������3�<=�Ѓ�����a��0�D$�E�b�?�R�Bm��F��ߴ�%
UK��8����������k��RƧ>��k_��SN���SNy��]���o������D�*���Ȓ��0&��3�o��V��R��^uC����oe���対��Q�}�����NZ�ti��;�8nqk`j"�)s.I<�5�MǞm+[=6��e�qI�]�,tH�Q������E�_�S�Rؘ*oZ��0Y�S�_�٥���?w���y�G�������s�����b��re�` Ҕ�S��M�M�16��L.� �@nj&���d��"a跿}d��~��Z;�BVG#����Bt�i��p�����?�~�d|���G��bT�������1g�Li�500 �o�m���Z��e�]�p�%�Ă}cS��x�)���'�J��A��f�1T�WZk"������\�믿
�DU���@.{���HED5�u�*�EIh�������ъ�C�}��-�@�R���䮩�b�������A��
�a{{A��_
,&�䁠�	~?����z�>2�E�d�7e��IŜ���*��ۻV�%%�@���(��fh`܊봮p
�$/��v�$�K�'���Hg$ҟ1�j�ƍ���˚��(�0�p���5�؍��0WenL$�\���	�8��c4�1�S��jPK��~;Q�uO8�1�J���h����8���8~����`&�k�U�u�!�>�ĸ)R��c�j���)x=���uK��Vr���I1`";���̶'Al�oܦ���ٔ�k�o$z�By�ιNKJ�LF�h�WM���uG�Ҟg�>��0l�YՊ+�-���O"<�~=��U�o��#�h�Z^�>�c��Sa���cL�X�dQļ�-9�X�x���-�Veܵ� l�^����L���X��Y��Wl�h���s�d�+Y�¤s�� �N;�v2I�Os��78����
è%�d2�f����i{{�@+�;a¸������ř�>��<�(�j2Yq�o)te�\Τ�����~��ex`�6a\|��Z�j���^{�<<[���':����UW]u��>���o_�`��M��	�#�Xj;Ԩ=��pR�@d󛬣ӦN�J���B8�?����p��_�c�׹�;N`>�T$?��{<��*�-�܃|{��C���#���?���i��0C	���8�t&�/7��,�>Dzz�!�7�8�+��leSn�H�:a��$��$:���P(��Ƅ	�Z��(�b�{'�K��
�o�N o8�Ht��cpp�mS��Nr:'�� �JUBMz^�D��&`C�rH�q�R�\.	xk�4@�X��k�x���r�f�Y�(�[�2I��V��'LȎ0:�<��@:)�R�,S�M@�^_�]�1i��Ġ�F��[�ӗFI&%�L�HI��tOE��e���D�1h��1�@�J������iH�#Al ]g$����0��O�t�ϲ�U�'��1,��@L�EO�\�%����	�sM����w7����,@ {ǟ�ST�BJ���}J��3?�,N�s������HH����wS9�����\�s�ąw�YoX���&�a����&?K����D���g����#���)ND?�*�)Su��b�'�3��L�;�ǡW�S����:H���xA�`�a}B��'L�m�N�u�������2i2� ��g��d6�c��	�f�!ʘ)�{ȟ�MaP�Uf��R�n���ɷl�XS�w.��_�f�đ"�Q8F�"z,e��'�I�Q(VM����G����uV��V�R|6Bз
���xD)��a��cC��M��Z���.�X�0�`���Pd?�C��a�:���EB�O�0�8�>����l~J*��j�Sh��3x�[)?��v�ƺ��N	�gx�"^�J�L�c�x`��0�+�O\��:,�׷�I�*Lm��̘�*��e&�����:>�`̵����Z1��e��aa`x�n��i�j���<0$��P��q�S�x�@��d���ab�ۓW�2��	�e�vT�Lc�p�g�͟*g̺�W�L�$�0a\�݋�����|�s)'���Z���d���~z������_�P�^ه�"k!4�����e�[��^`���:`�[5��&ˈ�}�&Fd�S����a��hC�D�k9�m��n�F�U��2�D��,�4��BoQ�^����C_���ڔ�|���O��''c�3V�Cx�s�]{-}����ț+�`����\8���+�h=����++���������|����Ь^�����+_U�}&5^��yU�_8�4�1a�8���y|�������rՊ���N�M}���'?��<�����[�CF�Ȼ�������p/M��5cƋ/�Y]�-E:��(���ul���,5$7cF[��[4���#�X�ݫ�Z�:��k>1����V�~Xd!Ϝ!8��&Q`T*7�s*�T'����a8�N[:AնxU�-vg�R���g	1�ޠ9'��y�rW�^K�Лc��k���J�8�2���yQ*��avEp[~���o��Lyh��2�N+��]��SO>��1���ʹ"/m�N:��N��u���o���z#������&<�|⫞�5��a6���i���cPkPF�[�0l;��e�2�Y���E����~߈�]���Ӱ��(2*�遨�S,v��I��������l�a�2���A4�e�6&[6�Ҵgm�1�0n��?�;�����:u�df���%N��<6��5����AZe�������wڐ�E5��c*�����Yfª8*6�{�:n"#e�3FD���15�f��K���Ղm
�TM}������B���H%Ū�;N��xm�>V�q<�Ib��f�v=2~z��~��j�H{��^s��7�ڊ�������]uH͇�{vY��ӴE^Y<Ł�=�Rۜ ��+�� �5n�7z�7F��l�1�]z�7?������O#�/N��q[��'��s3��&��1���t�)�GFF�����(ӂɏQǣ�l����:r���L;��^s��6yٖ�ڎ���sh��������>Y��Q��m�o��T(l�m�{��]�2�,�a�ෞ�e���J`K�cID7
׍!P뇬��\ެ�N����j��/��y�5p4��>�v=��΁0GE�c�v�1-�@����۳���(�e��ݨ�{�r�Ƌ<�۴׉;0��]��H!��M{6	,����
�A�ӑ����y�в!�R�y
����:'�`k�0e�qVN�6��z8���1���9�C�
a](d�Q�Lo�V*9��08p$3Q��4����<~�i��R���*Q���M�ԫ�O�;�����l+�E��0����5>-q�����.��h�.;�`��`e�ژ[�\�VU�{��S��R�����G$�v�ܝ2�IAy��R/Q���Y�y����e�yU�8�E�De��jmE�&F.\��ڱ���pb'O|�뼉v��7�9���Z��z��[��$�a	�p���K+�Ӯs����p�������P�_O��/�ܗ�A�]Z��E��TIt6�l��l��LhU������������p㭉������yÝ�M%6��TF����ub�H��z�H5w6Kܜx8�z������,����A}�=�LEU*�j��6�9M�"�?���akǕ.�&��}l(�APhR/�G�bA��iȿR�'�=��I�=���UQ�$�A⼍A�!��x�^�F�+ejgkg��D�gH&?�K�O��(*Ih��>?�_���PY�V��o�� N]lɬ��aȵ���R��<d��L�� ������FיS֘`�8>��e
m����2��^�~�}y�u�oh�,�01��L�Q*����ג��S?�bŘC��f�cJ�0���Iq�d�m�R�F��ވ�e���(�����"�%?m���]B�(G :�	�4��g�-O�R?�%B�� �hC�7��,�l҈=F���ұ@�G�
�#0a�g�̚󹙔�����	i�0�6"��X��ux��������ƈ�2F��U=1�R��O]v̧Y�P�;�?�A�d]b5مN&��{;��NN6Es+K�PVd�V��m�_��=�}�T	ҁ\+`�� b6�z����� .'��  T?+=�g�������r)
�a&eD�j��`q�C��D���qX��+�Y`�e�XD8F�O�"-��wl�~Z�6D�2�E��&/�̈́P���N�ya��!6f:�(��Ї�7̒�`H(*�f�XBw- �d�� L�ejc%���b��/%<^�E�����KT��M7vRi96�P����ׂ�����%�ʴ��R�t
�R�qP.�F�؇�7�y&e�GT4�� JF �G�����`����+��,X4~�]���l�͗0M��K�h�&�v��)�����x��L*��>X4C�
;)�^#r�<_���o?��h`�� AVȊZ�#VH����5h"����w"�G�χK�]�Akʒ�p�y,F|�T,f�>��1���+zP�D�C�d��"�L� ���L���X;,ZB_�"�!�m���3��I��2�tA��D�
0�V�b��9EԄA25GQ8sɄ�BJG�� ��e�?�)�J�]�����X"�J��|QF-��.�j���0D$�S>/�
>�7d!Գ(U�l,�0�J�r@��<bšDgRt3�����q�r�M�F�T����[�S��V��;�&%n���6���Ĉ���G��^4yc�Ԉ��6�$���(�6-�\H'�p��P�
�MWēMUb ����WFT$��m=m6>D_/䟞(%���D�Hq9C�|%>#э�rMj��P�91�y���#���{C�Ew
c��"�_���ޘ��|���3R8E�(�.�Cs:\_�|Yej��cXcG
3�5�Dk��^djq����;�R%��0�ݑ(�"!��9��P���'�D�C��W�/�J_��{$�(9���,�G$,�l&�	W?T�b�sX��
y�9e�B�
�iQB��}�ܲ��`��1��Q}O��8�|���(�0�c�F��(W��:5�Zdَbq��WT�v�T}�g��}@/*`G�՛Ĳ4ʊ��Uiu�;p��5C�e��D�	X�����	&��(9��f��p�^�H+�X�HqAc��J��4��v��H�[�8�1��>�d�����G�m�,�S�u'�>b�����BP�q}�R�5SDф�|V���x�.j�#6�M-�#q�Í��F��5�U�]�+�M�/L&(1g�������������X�bs.L)	����(�b7�[�2��B�ն�;��w�S$�Ѱ��~�h�T�,��<�Ta�_�
�{SX����8 n~����7#�,d(�4�h�4ŬS;
[�����xN3���"�E��j�ǉ�9�a��8Ƹn�(pvf��7�T�b���Q�Y�ld)U�PրUi�Y���bd�1��8���x��q�k(=A�%W�.N�9@鸇��6��6�H�~"1_�=\���&�и6a@y��3�\l��&��GyT%42��`�q0ڢ!�`]�b�ITi��xp�0O%�n��[X��Ӵ�G8m�1��q��NciKqb����	c\#VR���@�66��g�����O�� ea�D�(d��q�dL�K�&����/>���b�6s��J�T��UWe #��w�*�v�4d�4e%4N�F��L	���XU뺎��*:1�� g���i�h�9Hy��sfQ��$`�cS��aJ<@�a�邖���%bK�h�ڃ5��5��X�-�s�����#�g�Y�0aq7�{&0 I6N�8�bļ�,Y �f�E�B৞�z�Q��t�OJ�Mg�Ao`����Y��<�ê� ���������Ar��^��!�� ��'mJ����2q���sT�2�@��K����(�-��9�	,,�D��4k�:�<�2�4��I��< �: 8sr���T3�;�c����fnQ���i�[}�e����"B�j���w�b��mJ,V=;�&{�Z�Mִ�@F8�R=�aċ��J�.S�]y~�6f�i������W'7��)S�O��DQ���m�PDQ���xd;���xK��d��A?�d�����+N$J_�(Fù���P��fã;�!q!'��������H�O�Kވ��"T=�JL����
|_&p+�'+,�����aQY��?��3���+�e��,X���O4�ﻶ8�&:�h�$��W�'ɤ���9�M�ޫ�rh�e�c�H��H$�XIq�b#��0qYQo LS+ ߫0����+�H�Xs'^�����e�\Wi9��i���I�E���$M��	8�T�8���F��� �jHWg��Qۜ�C���"��:�ق�Ļ�(mz���ɅŐ%J9��L��e+/0�ϊ<b����	�X(s�1R�g���$FICX1���@�c��,�W���=}T(��*�F�
��,o��� �j�)�0��1�ɫiժ�|BJb� �������R���7�o��Z{� �IT���$�u!6I���Sy�^[��A4��K��1qx�:�9C/K��	ϟbQ�fh�LY�2_�.��:�N���(�#�f�N3����>�Hq�!Kt�(gieSG*C�ę���@,�b�����,�"�&�cK��F����UQe��㇅�Jj-���;�#�Y����W(�1A�9*ȸ)����;h(J�uR��X_�q����wS;�D�h$!oڀs*`�XW�5����l����O��sur&���Rm4�{��,�||��2hwQ��x>X�j��!�'�A��J�T*�y&�
�_�bT�c6�� J��1�'Fb�Xm�#*� /@�����4C^,�x9,V:�[%yRBA��X����	��Z�,k�a�5r�a����]1a���ڌ�tl'A<���iPܘ��}��t"Oղi0.(���q���!$y�E&�
s7q剗��P�]��\�N�_�����N��>d��C�X�*���� �o��&�Ԭ=���YN�<v�I"ǋ�:ZL.�j7j��m1�P��7S�6�S���r9��g&d���Krt�z�-`B>M��i����/1q�
��f��9֮s�Q�aa��FcP�L�����s<ǩ"&�&]�V�C�R3i��Aui�w��$��_�TYl�G�%L��c�e�N�)����}�,> �)��0��z!RO��56QbF�V@��i�1'OE֜ײ������s���ryuX��]_��ꄋ���^���*�;�l۲��>E=QAN[��XD �v����(�ǒ9��9��N	H�CQJ��<���F���	Ew	"�1aDl��R���Y�xc#�Zz�.�]L�Y����{2W�dR��fѐ�c������k�#�ֳh�W��Úc��G��D�&쨋��h=ǈt��j��)��Yc��'ކYa��~����L�U���@S��.3G���8iz%��o�	Wx+QM�O�9��Ma�s! }"�P���	#�,[��\
�T��"�Ֆ���32$Fo����x7S:��f"B#��b���u��>�F�:EA�0 ��u� )����(����U�_N�oX�QJ+��j=d��#��ۈ*�ߘ��U51��ŏ���2J�K�������ʬj��M�I�\�I���F .���zVEW��H]�H�F1��]��j�Ni��u�GM!�
b�/	T�U棸J,
ewF�x/Ԡg�pr�MQ�~���§��8u�W>�H=h(1I�B2��b�a�U�C!���0�8��L��= L=��5��&J�5��G	�N���t�ر������2���c
�K��]�K%)����^���rRH.S�bI��aE�"��Dj�L|�����Ig�ћ$M"V�6��� 55Ľ�Xob<B���3�1�B�u��g�5R�	_j��G#3���&!*xK��c�J4�h����$�@�{_��u���RJD�<�OLlDԌAR�K�B��j#"Smr�)4~.�HGx�i�@L�d�k�i����e����hXE�Òg�@#��"3�֐�`���¶N۰5��z�T>73�HF�s$�������J94����������a�a�cWU�� CgV�-�G�hK����6�c��9'��ǖ�M𼂫h�7�Ok�(C�.�M�Ex�r�)`��TF�4D!A���Ñ2UVL���%�BHEmC�)�J$vMPǰ���ݫج��vA`�á"- Ԃ�fɡV��u�-Pe>�B�x�n.�xf��@e�+(P�;��fJ`"B*��RJ���R�l�&z���@����:J�]�~}E4��E�w��|&U�-��s�Ɏ96D۬�$6��]�la�n��%2U��V��g�d��H��,Ca.BC��f�'p���@R��Vk5�]^ac�K�/�7��4C��" �%b�R1QD.��&���r=��|�8#�l��gR>[sE�Fl���:�9��G�ceu�C�� b-zH�*F���'��6	�3��6��uٮ���H>����QO����OB�tq�H@>��T|�]b�=��Q�[��K	�R���~C�Vt�0)3I�Y���ua+.c4�9��G��H/�Dt$�*��<�5	?�!bn���5��'�X�0�cC�������_]��U]JB��Pu*��'�~�ծ�C���C%*2���i�s�CQ�Ė��W of
KV-Q\-����g��p��@��P5�ee��بD#h`*c��K��Td�P"I<��b��\���馩ce(���U��YA��6�Y�9Y������r�� ��^�\�@�rI�c]Х�����t���|��m�i�	�75�GV<"�m��)R#3�K�xQw�;�-��������L�Hsg̢:9�3R�R�����ry�"��T;��p'^NW)���i�c�!{���w��uk������U��Ux�r�i�P7��c�)��ԙs9)�x��ixs��>�r�5��|�,���bţ0�Pn.[ ��VA
e�Y�dޥ��\�t�]\�N&+DЖM���NTJdY���Di�ζv���g�à��6�_ˇ���*���`�*�%�I�����ja�	cc�.I�x�b�Lg|?z�e�'�7P
������Y9{�fP��3�|ǟ��/�P��)���R�r�H��}팝��K3�6+ǚŮ���]������3�U�pTS�\*נx����R.��b�`�S:;��,xa8|��^@պ'Չ�s�Z�*��(�L�" �2b�gsm�;��5R���4���V���LA���v*R.D晋Ʈ4P*Q���JuO�7��2�<g�#�B*b��զ&��h=�����% `�o�#́�/jh.��57<G�y�L~o��3��3OڃY:@�W=A5�sYތH�Oc�&��A����e�Sɢ�5͞Ӭ��i��i4��#�u��D��5��L�u��a�`������6�������I�:�;�8T��y��������=��C]S
⓱b��������S-ɯ�T��ďA�j�ژ�Qq-�S̩�}�N>VS��w����+��)�E�P�Z�klvQҌ��U���T(�,>P�J�b�O@%v�hM�F��<
m�=����]��󎦽:��������Oh�L�����f*�]s�3��&N���g�C���V3[�@�4�4E�_�5����7���1�{��Ī�ۦS�u�����wҒ����;�F�z����^�ǖ,�߬�:+�(�]G@�Jo{�|�6�[�R���2�˫=��s���A����6��޵�n4�};Z��rzt�2ZSdn6c��F:�s�Ϗ>H��:�FE#Cw?��E^A��b�*9�/eM���;�=�@��	c>�2��$�2LV���cy�tC˱� wb�O5!Y�ev�V��%ϧ.6W�t,q���{�dyfO�z����TH���נR��U����B�$z�L��^��v���o{����_,"�0��2��3��ϡ}�a�Δ��Υ��w.�{�誟�KSXtt�N�s�NL5W�m>辍n[���0K�t�>�h�;�q��4�Ŝ飴]t�r���%T��m;��>w�,�ޟK'��?���h{�]�ɺ��}�mM�DԢ��K��C�jLS�X�o��u1�sR��xuCխ�ݩ��P����Þ����O=K�f�@eF
��TDَ<�q�+��_�N�6�˶���n�1+��n�~��(CCk_�?s<��D��@O/]EUՍ?L;���^T��*Ma֎�co�=EG��m������S[@�ٓ���K�����N#�+g|���O'��jƌ<�Ȁf���`G�&�Ǘ�x��.Ru���}���鵥���DN�j��D�ͫ�D�|��5�)�1���'&�%��8Nb��T�e6��gd�c�Cec'�J��.E�L�WV��j��rJU�>�߼�������މ���V��T���Ot�^�U+ג��A��p31�����=����)8��t��t����>���|���_)�wSG[��Ţg]A/��Y*t�(Up������Bއ����Rɤ���G��ȓ�ߖ�~�`���=w������~�`0my�ӦvRƝFC3�r]�T+�N:R�q��p;���g�a���.��t��С{̡�|��W6�7����>�gr;w��U@�6[=�H$Ш�P�D_Z^e���h����H<��M���T���c&c�-rT_��,>}#���K'���t���oK����CV�2)��E�jm�X"��&�,��;�?��~������_!�}Gr]��̻aV�	�urbjZ�n��g��wn5h�C���}|;�cv�~��g�}j�fg���:���O� /��"Ųf��X`���=g������&������W���<��{������˾y
=�2s�_<NO=��ܮn��Y9�E��{eo?��S%9{���K˗	G�u�)R��ηK��g_x���v&��L�
�$�}�e�R�*	��;Q�vC�j�nc�4GUhA����C<�JG�y�$�ꬿ1�Jƍ���Nk�B��O��=_��6Ņ�*��zY�ɰY����>�	H������}����NL�_�yz�Q�Ko���A��LA�TI�R��葕颊��H�m����u}�����L�;�$č�zm�z�dQ�Γ_���ZCKW������f�B\b��������VV�}�ܛh���л�K��>��g���C=���)}}��Nz�C�C},��R��M�*���YJg34X,��`�:��"+�[gp�	�(�E�P�W�!�C�FO��=�Di�����,�H�(���[_i�[@���]�3R���VO�
�%��03���̲1i�tɝ:�V+���W�>���nt����1�?�[j�兒�5Xe��k�f��YNէ뮿��z�I4�Z��2)F��*��7�G~��t�G����ffS-T�.L�[W&�Jp���8)�'�*�*�f3a9y���ӭ�Wҭ����oٖ.:k�y��韮�9��uLgQӖ�� �M݆*}EVZۉi�V�؄-I�:9<�+�XgE<�fn���W��Т[��ſj8B$k�u�*cH삂��m)���@"k,e������g!,��_<a*�'��)��&"nqKN��e%U1���z�CA�ewz:���􁃷�SNؙ~��+R�=9�٬@�C��U�y����֮RT��>�@��˯��5��5D{�-��c��S{�@��O�7{6E�L9�(Y)��&��,[E�j/�Cm�5[(��@Zߚ54���?��O=F=����N�V3Kx�W��mK��so�颧�(W���#=PD�ݿ{�RLxq�� /W���1��L$�C>����pB1�"��L����R�0��4
.j�b��0b�{A���oF�['�W"8�並�*�@$�t2L �����L�G�Iz�C��R���H����|�?[����˶��7<E�|��t�GХW�GS�fP=����Ot�ns�c����DԻf�,����=w1��'�0�X�L�MW��t������s��ޗ�^�mfmO;��AW^�$�i�R>}3�d�Q-����T��9�O���Y;����h�w��I䱂�ڒ?S�����hG�W��˄m�ѿ�F��mK��z˜����>Ms�sz�M�����WXL�ie����X� bf��0'AV�ҋ�fPcˌ���d$Y=*4���*a�t<%��a��.�k)�16s5�6ݏ�S����$)EGU��zN�i� ѫ��t2�~z
=����f��LTO�iy碷�n��l.�؆�eJ�w�@�����
�|�4�f�c[*��'���_��=�2��N�ryz�%t��K���^:�sD4�ġ��Ѳ���A��
���Y})��ζ.�f���f���c��N9r�cޮ��S�_K�_��D����,�"Χ�^r}����C����'�f�r��k��w>Jv���c�;OO� Zœ�����S�4"�ď�RcV����ƪ4�I&���^(d�ш�*���!�	����F�%E	�3�S����.��`
T�M��s�J6���`��ѓ���w/b{{;�U�6���x�T������28eZ7[Lrn���֣~���L������`����g��B��V�C�C����=�)���W�be�����P��K��U�εI���`���^���>��{�k�j�nz`�tσ��D��NQ�Q��]X5�K��k��ϟ��n7���*��<�X2 �e����^��K^�+���ɢ�g_�;R ��JRyQx�(��.����+�N2O�hbH��e������p�&����g�~A�L���� �����S�PQWVP���uH�j�/	�>@	Hf��w���Q�!h�Fqp�P��FTc�5t;�$!��i�WA
CPS����)TD�8+���`_ޜ���b�L��,6��J	'B�ӻ����_���i;�[G���HY�q2�C�mn�#P��$�XJO�#��k,G>����p�Ä���!��ܬ�d �{K��b�l��3V����4x(�b�O���aB��Gg�t����@��q�p��o�v/�k"�
�S���ME9�5/}_`.���B��À	�C�'9]"�,S����P�[ .*�,-m
���*�WbK()m���A�=�m�+b�s��B`{��Ҩ�㤔R͛�+�F�g?	3�����������
Ѻ��<�X�%��B(=���ʉba�l�j�l]��a����*.p�=c���Y�'&VR�-䚘�n�
,���_�V�RA�H}2�GUAccI Nc!��U��G�e��J@��7�AJ?M�O�@���T=T�A��T
EN|i!)�Qc��P7(.����Cĕ)�{2�Ȗ������n��Mq/��#�%a��s1���"���b��(�^�RU��������� ��!PB�-��,Sk�MJ��!�rb�5' ��p�T�J����Zj����G�A[���yҗ�?���QT�ut5�WY|�'�<��/�k;��0�y1@��U�S���wL��NDo9a[�п��yA�@��*a9�eE�/R��Q����X�6�t"g�)Ś���V��/�`��'R�l$ʲI�Y^ &D�!@8 Ѡ{uʲ�$ռX
Jy���l��5\�y���8�R@N��8�9(Ub��3�V����0��t�s�
��d�mR����8�XԘn�P��V��51E�Y�x�� ��͵���<�����T
]Ή��pe]��]pٔ�P�֕ �X<�K���<���(
�b���yUI�����C� 5��U���	`�+tba��	��v�R�+��,��eQ���	��h��I��@�����ErA�<�j��rA<ӑT��-&$p+�l�.��M: �D.��1� ���LmF�C���!��݉�`���	��@8�ͬޯ�s�r��t@2T��@O��a�5 �
O�*�T����e3қb�R~X1��@2oul��\>��t#I�,y�A��٬bV�PJ���׵�(��6{FG�8Y9ˣ�W�P��*�_���f҂R
�jC�h� ����8�N�ιT���IʋfI�;X�S`�Pz�E�{��L&(xUQ|%��*W� !@�\p� �w6!�)����s1,0�[&B�yl+�,����Tx��[$Y�!0���y}͛
L)����!g�n������,:@U�O�*}+�//�bsHǄ��e̛��k�G���*��<Wg:M�>�� R����gB˸!�X'q��4��%�mTS�@w|B�^�s]�H}Op|��v�ڶ��(�Tc=��=��1J��1���U#��+7^I�Dk���$`(]@C��A$�
�w4��mw��Ա��T\�Q�*$������釩��Ս�0�+T�.��U�V�-�l!̢]�؎��4Q! .^�s��O�-�5��x?��TH�*u�G���z�#s�&;�N����̳V�����]�C/>��'���ST�~K圲|ϰ�8F5u}��#p�}h��?C%t(w��D�c"��x���??I�������v�K���!uN��5P��/���?w!��n�i�������A�o���@���g~��e�����(�0XT��-�4��L&G�����IauP���l�y�!�A�'�v�9��y���
��{���B��N�QřT�'�レW������_,�c����\CJ&�L�Pl��#^�iوf�;�v�1�Y�R��k��9�)���Eǭ��AO,롔W!�S��<s�|�u���\L��wo:e���5m�A�ʞ�,��3Xl�T�n��b���s��l���e��0���Ru�������fNTa�H�/b��h�DA.27~�5t�od�X�����'}�bS�3"~�'��1�5�E��\���6D�n,09'@[&պ
� �D4��giv;��� �Ѽ�	�w�芹�O!��Q[.m�������󑥓yP#�9�\�)Lp]i���*���7|D)E�;�i�	������+�E��iR��Y�E
���H~2���x���# i*�ZET{����M{��Ւ������b���b��כ��� n���q!��q�c�YA.�/�k���^#�Q#ҡt�cBj��F���*K��|�����pC�Ft���kؔ�H꧅��}��iC�e�uO��@�fٌ�E�2��{6��rq���4���3a��|���AJB�p �ԅ�&f�_3���&I���9�p�C�ur"#V�Z�� rB���$B�H�M�	���TX������%׍'u�F=P�bCu0lG5�&�R�R�M�+����q��|�8Pu� f��bԓ����F!:D��y�9N�)����
U44�k���5���yD��bh��-�_��÷�z��Q���~ �lE�ե�)C&�H7��m 6���cH G��(�v��L���-~~P$��R�����n�@��sǺ�f$VNzv�=���4t���2Y�W ��#
!kZ�����bV��L�)1W�r�4BK����gJ��##����瘽{��=� _��-���T�3y$���`H?�x�j]�d�\Z���J<��T�*�L�_I���t.��1p�2��=ߴ.�y����etKJ���{�:�M�Yʁ��߈Ԏ	<ޤf&�� l�*���}�ڵ�7����F��]�d@6By��,�8#�k8�$0��,�\I�'�(p�pU�$����K�Z�|���Hm8E)J�d�Rg�@�#I@B<:���T�"!vd���ä��@�Ռ���
C����J ��b*M�:��T�@E��GWrz-d��򘉠�x�̭`���)I 5?���Q�IٮqA��[8�Ⰱw�y'-^t�,8F6�j�~��E����˧�$�9m]$o��p�.^�.���
���:f ��iB�C�It���ZU�P`�H�_��T𹧞x�.|�/��N�J��}dQxA+v�WgQ�1�\ fE� .��"�^��sK�H�ܼ��H&rTsa$U�	�b
��z��]Ya1���Ɛ1\�UED#���(�?��ZJ�C��tEUX>lt�d��M��\P³&Y�9o�����5��%�!<�._Nk�RcS���q�r͆	
�){���]��c7Q�g��Q����^~��[Ջ��\%��~�4.��F,7|��R!2��¢�� �4ܲe�؊,�e��9� �NA�����i�+�C�T�PA�j|(�lGC�����ء����]R0=f��w��(��দ����a��Ǥ�[�,��T�$�Wzı���֧�s(�h�ƕ{`�c�ch}e�S���/7���C÷�:�&i!jd#`%�I}��l"�憱�!l|����7��-uC��b�I)�O)g���M��i�?��u95�>r�x��-�v7gش���t�q�aȦ&!p)0N� 7 ��=G7߷f8�~�ah�/8�'�8���~U��P}\��bC��J`Ѫ�}t��h]
i��n�f6,�&|�F�HQ2�lwY�jU60�\uBI���.RM[�H��}�D̤R���e��ͷO^�̵f�1��IZ����{:�3Ho�с>(���@�MD�noXA��'=�M�8<GC+¢�e�&�,4�Q��U,�()����d�|H��@�tD�F&Y�h���EJƽ./)nR)P��zS:Gi���T���b���+�F�
$��G%"{�j5N�p�X�G�ԼF^/f�����hː,r�g$'�AZ�l���=4T_5�u'�l���9�b%�ћ,�cP��O��zC)��q��M�Xx-�H��b��*�I\+�8,5��~*��V�VR�]B�Y�YI4�~����'8ҏ�DY�.����DJ���N=���L��Xz$l]m*563�UJ���aqE��d��6�q�Z��78�*����5�&�����Ł�:�(D��'�o�������:����A(�X��$��֩���br;�5G��i�u�HS�DFb�V�+)�I!�ULE\|r�tbQ�j�XR�Η�R��A���]R����|n�\�kl�jQ� wx�MK��_���F�"��Hİ�qZ�L]K'V�U~���|�:���0��Oƨ�����olA��S�E�tm��X�%f2D�IM�XNw�X���0�D�$AB�����7)
&iAb͑٤�5�X�r�H�q�J�׎�EL#=.ɻj��O<��-BE�5�'�
bڊ�%��F����b��0�M��#H8���/z2�eS�8N乮5ּß3�T��M;���Z8ĉ&@�@b�(����Nn�7^b=ڿ�|�GҬ���$��\�x	Qp������Es&���Yqn�|�5"�r�?#J��@�,�z[��@�Z
*a(΀^1D|F{mEq�_ƺy!� Z�|����4�Q��x��{��ـ��3}M�\�ډ���xƖԝ�8@�eDB�]�E��<)&�>�&�$Wץt:K�(%#���$nr��f?�'M����:�ǆ�a�s���~�+�r��ZO&�����M����D4��������f�~mD�%lisyx>�k8I�ў�X1��F��9#)�/(�f#"�ՒI��A��-5��X��5���ؔ��:I��Γ�=*b8!۳��L����bSߔX�/��0󖕇|�~뇆����8(3W~*�qC�S������3����[h��o�nh�=)��?D_}�K�S��Bۡ2���+V�A�5���[��W.ن����UOc �3���W �4��j������ت�$��_mW���'($g�hY��y�9��o"t����R,�u5m���l��wI��ύ�(��I�l)t�����I�H��:�ee�����q��rP$y5���>��8C!�%�,�7ְ�8P��Ke�cO���/^F�G�Uy���"�,�f�T���}������]��Im!I�������G�%UC�Ԙ �� �y1~��o�k��{2kub&�����Z�i��ZV��q.}���yC��	tP�L��� ذ�.ʼ���~�a����ӨR.�:&�~U�8W��+#e��������c`�D�2�Q�X���^we���G��:���t>h6^"�����3im� �ӷ/��D~����R;Rj�1a�wHFv��M��CC�(P��q��d��j&�Y*JP-A��A2U�����Te"�{��l�[ �:R�q�LS��-rR����s(䲴��QP#_��
^�z/�S
4��ç^�fT�&C�
b�/�@��K锋lR�yS�  �Ђ
���󔚳-}���h�\�t�cD�+�ӓ0�}O�@��8ڼq�.�o(�d�am����>�)ʙ��³	�#P�}�Ȧ]�Y�:����ԙ�P S@�i��zdk����#���qX%�+�@R����X��)}D�TֽPp��ՙ}cC0$�� �a�^�veG*�!kCu���Q�>M���-1� bº�<٬
�#��Uw�$�\E 4\�m�.p����!�P�sF2S�l��<�"��Yǔ؋�Ĉ���r֘;����$5Da�tB%j��d��=�|���I-H��*�-�n�z[D�� �Y���C�ֆE&�Z�����5�Ni��@�!pB�ZC74�z'	ϛ�*��V�T\��>�S
3�UA���
��)���Y� �am:���E6�Do�q�8l ,�i�]��a��, �ZI-	K�X��Ѵ]�y��{�U?�5�c�*/�a��Î��c	9�ir�4���(#�<�J�R���YY&B�9+�U�k�G��7�j(�r�(џ�������6�"T��+��"E��G�H����%�2HE$�7�xk���6`"o�0�[#ͺ9���2y)��0t��ʴ�Z�x����](�	������e)�e�Hl�Ʈ '��,VA
��Ϙɦ��pr �N��&�j| IP|� �C����AҸ�HR�IԵ�@��㴊^�VH��H� 3pS�/�X��r��{rr$����h�R~/a��H����\L[~5T:�'�A�JAL�ؒ�&X]Et�W���`��A;ɿ1�x� �Κi`�jŊ���{�[�U��
;�*Wu��PMGRC+ �(�p�>�
"���lT�\L�- ���%�D��n�s���\'���s��ϩSU�T5��}��+v�s�^{�9�s��? 6P���{������j4e
�� Gd��zm��tݼn�t���[@�.i)q6�0R��ܥ���	�Mم#m"�@�:+^C�xl����2!�����ma̜����J�,`,GS"��5� �\l����u��! W�\B�0�e�}"�p$���1HR�E�a�vN������H��S�o�R�A�K���d��bcЛ!��������إ�d����5,e=٫m��z\�ְ^_%��5�l-\���We�#|����O��2añz�\�
�S��p���VD��J�b;���v�u1�F5�,���J>�wi�BS�f�X��!���u�^(�U��He!�q�\�\����b�¡�߹J�m�AD����H�n4����v�Fq]��~o���6F��P�����������gMT~��螰{=�v>H{i�����{䋍��)<��/�6�d.�OCTkl�0�����g��U��}��U�Zް׌l`e����'�"��ᨅ�v�x�-\�l����#+�	����Ae���ρ�!�(Ҧ�����p���H桫;�R�nӊv��d�<�����L���+���%�XT����%?��=J�=+�<�K���I�F'�k/+�v�U��9��6?��}�Zg�*��[Q`�La�XeA;`O/V���U�;*yttȩ�q�/]!��U�"���tG��/Z ��@&BW�3��|9���Q�B_�F�-��X�Ќid�������2,O�.�!w�K�A�X]bd�Kaf#�ʀR��!�B*цQ6��q��ܴ0 t��U�A�:A�� �fcQX4�����)pH6Q���Y���y�]��i��.Ϣ��f* �nL-�v�%�]��ZMVJ����T�����l�,.LmC�,�'wQI��FS��_�8c��^Vny�Y�RL�GDAe�i5�5�W����p�0ϲ�<)̂���`��et��� 4J�><�1,	�6��)Ѐ��+>0s,���B�Y�m:AQuq��w��yV�oҎ�»i��*�`�vE0��'�ob�@����+-����"��L����H:F�_�"��mjC��\�{[�	��s=j�LG�!�BZx�z��8IՅ����.���Պ�]T��Ŭ9�ՙ��υ�}&����j��)�s��	(��UXw ��yMթ���؁μ�,i��PP���16���Za��U���X��������+���M]����(�o�pK�z_8�Z(åp�8<2��ƁұN4'{�_��)��ܒ��z��͒.�B��#S-I}��al��|�ν�

�͊��/8_�H[��.��>�,qU,��k7�3�Z��k�l�؄2�`H[�B��,k��y��T5AE@_'���I��m����	5zi��Н�Y1��3#
���<��f�F�}�;��L�����8�ź
8��C�ݑ��pz�b'���Zp���3o���[���1*����<F����-\f�}/�@εF%�Mb#� uc��}X��ݷ
�.D`5!�������G�\~�:��8�q���P�h�k5�.t�[>4��Ѣ��otR�s�	P��깎� {1���s_�,1NRY�s�ե�8���u� 3��֪����.SF���zt=�%*"v��PP�{�Ư(��5qWݼs$a�,集
,�P!��K�ّlKo����4��Y�gӧ�Wg���K����T>�3~|R~�ޫ��0�Q��XN ��˂�Gi�-97ͱ[h�U���`ߏ�j�	DY]f0>�&�XPL���\�AI�� ��|�C�|�v�Y .T�{�����[��Z�w���pж������5p��l��✹��Zs�9,r��!g|�
��7v�T�q�[H<�׀%�Giuu��PL(�TG�vY1�tn�,׶ �5w6�-1��q��~���7�n�=A���]�ɰ�%�UQL��?��ی[��������D���wcY��E7e�n�Ge��TaƲ�쮪t����:C6��J5hf�N5��@�����ӻ��j#4�5LF�wzd�w��r�Li�̭���`"�{鉱��(\ř~6T?�` ���**�V?��ĥ:�X%k q:kU�;}ͼ�Z������HS����}ZGr��!Υh�u�l�$YҬ%� �l��F�DE"���
��L.��X���@�x`�af���<�>�h����`�ff?�����A6t�^U�$
,:�e���a&x9L���bh�
��/�Ԡ��c�2���:�Y�`A�9��/��$a��硆l#n�2*�r��瞑ZX Q��QW�Y>�<�`�A�nQ�UH=Gܥ#��Q3bx�:��I���*�D��պL�����D���P�N�-��6�j�g����b\.��ws��2]�x�C�p�D�����C�G��%��pp�v^�8�yO�7��
0�la�]���!��Z��0C�x�WG�P���D�I��>��a%0��Tpa6���j:�қ���<�s/C�3��x���J�|�g�>s�΁!�C��~���}"��� u�-�)f0��`��X�1V3EH^W���Şu���ݕa��IbB��w�^�EB8��P�6ѐ��;�W�D�z��$�A72�@4Ks�z�|my�����Jn���%�����!�4!���WZ8(��iny�^�D�ZD���Yw���u����JS�� !�U"cĬ+mm�.��R	�
J
gZd��-3r
e4�4
�g�<!q���,���0�%.��dlTDd4���P����������P3�)Q�������j��������/w�F��6��?��r���b�G�%��l����`K$�I��eW�����\��7������������!�|;�>�v_���|�&.���!AA̼�l�O���%z$ϥ;L�Zv��t�V	���KQg�,�(��T
�\̾�y���~#�'�Z.[��W}6m�6�sM˻ ]
;+�@��
�}��f�9�f�G�j��1&�A���
4>�:�>�tSm�^q�B7+u��^p�mw�o��>Te�eH_5u�,^���zo�B(�bb���;����mh$�)4-�܋g�}�F�T�$*.��ۡN�W��-���,��.��Y�*v�y�\��
9��ݻ8ğ���0-����i#̓d6d�YS��Q�Q��w�43T��<-�{V�x���"DY�����OGd�q�0`�42���������Q4����ް��~������ŉU�m� ��pWDJ�ߎ٪��\U� 5:&�����T�a&i�Ҙ
/��̶���z�E�����~b4��/�E�Wg�R)_�ٛ+���5�C�7�ό�شc
�c&C�����Ǚ�6�s�U�E���2�-���aT��k(GU����'��T��F�`�o|��ȿ�Ux$3\�9&J劓����>�pn�]�	ga�1D ���9��N,��	>�8��HW��*�}�,�|�`��W�m�O�Xl��3 �bע��}�f�r���+�0�@��͊,L����{r�K2�K ��c���i1";�i����-/C�N�ZB���-9�d]Qrj�2�9N�&�H��̊���=�ϵ�4W��X+�G���0%�ݨO�{�n�v��6��#�in��$��5(
�?r���쇻H���E���1T>���Ԙ,�����6�g]!��}t������|O���Υ,�!��xJ-@5�"�*ɮ�z�+���'�S0ږ�΁½$��՛.f�3���"{C��I�B�}�>�X��ϋ��`h�ܣ��E�
�/h0�р��QXÒ,��K_�2[�>h�7�Uq�D[���l4�:�Z���ܠ�!F(�B����=����7��n��;�F����zzSvZ����fw���M���0L�T���Ȫ�#K���j�3��f��v��ڝ��wYp�G

6��c	� ��7d����^WR��2�hN͡GHC�����E0,��ʼ�US��(������5F�סU��R�)�
�X���*e�(_N�b�0f4.�>���Tm�HIIe���Нi^��M��&[���ɟך��~�\��w�Ei-��i��k���Sb�,n�<���F�sT���w��-�$�f1��s��4 �tM�Rr��b$uW����*��|��iw-���.�Ϋ�
��&��:53'�`�p2u�%#�!������ה��P���ke`�Kj�2��n����a�C��,�%�J
p�!u�W��P�$tY[U �Hw>^�cÓ������0�B�M�o�>	.�1��ݾO��!`� �1L�P�0\ڨ��r��ah�AUl"�ϒj�v�u1ִ��`=G/Z��f�����0�0��K�Q#�Q�ѓ�C��@��}:�=b��	�Y��\f+�Wt:��0�PC4좑�P4�p�Tu����,��@p͚�ϑ���a��r�n�|j�Vj^�>�X]0��T�;	]��ik����;�:�p9�xB�qu��C�'�Da�պ�0FCw�裨�������	��x%6B��ev Z�뿎Żn�x	��>tn��y��X諺U�0��ynGq����ð�I1��;o�[���Z��j�Lե�s,�9}|�C�ð�F��*�{�s�Q�j���7X������׿���[s<[<�w�󝘒3T�?�Y6�Q��� W���݊~�t��#?����)���(\8��' �b�Z���s�v�DMͤ>��3�)�q�h�5�F]��p�5�B[dՄ�zwӒ�#c�ӊqt_KTv�O��v��ۀ� 6��\O����-c<�5aF�GVm
�[�c4b�E_��W��K�ߊ>P�G��=���W�0�5��nY���Pc�I�d�k�{�]s�w5��[���'?����"��������ǩ��0+��6Q�fk���5�a�qQ��%�&8��c!�o��@	N�1I'!/W��(lyc�Q�<K���^'=68H�qA�B~���0���ep�
d�Պ%ȝ!�X>��i	�Iu	��2����G����MEgD�g�A%�L���#�b('�,?�C�x\oԔ[�%o�LfM/��g�NL$�W� o����F�F-W��A����z�P�����:�CW8��'�l��ԁ��p[��ŧ��1��,7�f>W���J��J0a��i�c0_��p�9\3h`1w2��/��X��Ɛ��!�e������G�����͉�E���\�z<��;��� Y�2L����<`3��+��+]ݴ��n�s1~Vj&���BSs�D:���� ��!��"��D{Ք���+y�ۑ�H��X�4PF��A^X'��OF�$�(���9��rNj�ɲF��^���a�,L��>sJ�\%>�6���H�Pj+~�J��-\J8��s�*�d*����!{lt���$T��d,�K�����v&�n��R�Z."�Mt?X����\^&���5bEV��H��G�T/#�ˣ�O��c<��h�m�-��lsЩ,�
|
��N}��qҞ�\V��F-�v������F�%,C)�j+���tz_�s����E��=��R�j�0S�si��l�[4��eyc?���Zv�%y����l�0i�\�Y%����p�ى��^��uW&���3����m4�Se4d��j��r��\�ء����׮���������XHá��W��9��r�3b�u�7~@ꈀ��U�s�p����i��3�z-���\�F%����Hܢ�(�W�ԹID���$0ʊ�0�Ct�*6?c6�V?jq�����䮖�ԁ��y�P{�QrG儮f5O�jy�8?����劣�cC|ٟ�/��V��u��:�YK�4���p�d������B��b�����zf���>��3�׺������h�lҠ^��f�S���*Vh��C]dj���!,,�Ccj��h�kDXL�$�z��=�Z�J[	w�K��P���]��13�p�uX8�X,���+wlP��`�Z���X�xbT�:b���a�bLD �a��'�@ֶ�z��6Xոb|wĀ'�wsfN�K�b����Q�k?�#�[��[��.�$��F�k���Z��`�#�� �O��fU�b�V����O��d��M8���H��X٢���f�J�#N��B�ZeZ���μ�"T�ieVL���Q�0��=�����D��AY%cS��A��P�S�qR��5�ﰿ�ܪ�iH�=�B��3��W��/*�͋�ُ{���oV��[�0�q'6nݩU�D�ٲu;��E�sF�Q��Ë��Cp��3l�n����a�����X�N��R��q�]D�]¶3��h�u5<��޽���_�+x���e�y�h9^f[b��p�w���}����s�05C(��QmlG_��bs�Y��Z35�����>Pv"c�����������`����'5�5k���{�`��p�����?���6�U�%.�d��G�.QwX��*��X,����{�w����;о�غ�Q�u�` ڦ֘B��]|�Y$b�(~W	}ߌS�$�50��*K�h��٬e��Cr�����2�ۮ�]����ڌj��ޔ܁ͧ��FA��p�9���5�Hs��o��G����5��3�}݀Ab-�A�2����$���G�	Z+���$#-3��:VP�1��e����p��ؼ�j�ɹ��[?�]7|��kO�G��AqMOd�dh57b4*�I2J���>����<Įͳ�=�sӗ����T,C;�Y��J��pB��R�2Nr��w��'9*��u;�VU��,�b����[����_��?v1���/��s����7݂g=���W��٭h���Q�"m3�?{��>�q�>�t��s������K.C�9����7��g0���	�ic�Қ�5E��2>��A�&j��_��C{P���/an�"��~��ֿ(d�7?��8��]hGm��]���|�tӍx��~oz�_cq� j�Z�6��uo§>�y�&��A��K�?7\w5��18���\`���5��?�J}Sr|՚-9b3@1Av�`�� �W1"7l���� ��!->|׷p�Eg���y��/�Қִ:�t��E�X.��|����g?oy�[�`�E(^����شq3Z�SZ�ڜe��H=��/�?f�؉�����'cnF��Զ# ����*|��r]'2V�DO�k���o�͠ڌ�_X@�x'���g]�{��y0���w���e�k
��n���]���/�Kq������=�T��]BF�(ǵ�݋G���q�/�<���{ދl����3P��&�����2�t�B�qJc��`�D-�`���H�:6NGX�� �q��.�K���g>K������s�t�mk�c�y��/~��睳K���DTd�%w�w�Kv����ڨ0'��?�����w�̳��\�T�2^8s�8Y{�sU��`����LqcZ���b� ُ��{p��b3�G苇��g�� ���û���Ӵ%!��}"�u�%���M
�Y"m'�V�bW�$B� ��oԞbc�� �s����P�R"m{��;w�x�ەl�k����S���%�r�
�9R]"!�r4���B6w�zأ���R�h�����g?_��y����(GG[<����#��h��Zo�,��7ߌ��/ğ��r�v`������.�o�q0���t�����(���O�g9����z����V{	ƂR8LgZ�J��$b~�0zK��P�g��x��]�L�,݃�-m���5���bt�\������'�u�����u�1.����܅�/����w-�E��"]v)�Ze��{�ޡ6G/_@%l�ݚFczڪ�
�q0��p�j���ˑ��T�kR[(敫�����()z�ƬW�<q��m$�k�����eg�Ш��s�]���06��!�i�u��WkX��Y.���L��&��A4�����P������J�(B�6i[$V�	1E8�t�be��)�q��`�E���#�*c�cܒ�5�$�CZhWW�;�f��ލ����E�,uPW$�PqA���/�u�zl<m¦�(DX���%��7��s7����/x�s18�u"7�e�aϡ�\o�μ�B�$�+y�0D��-��}# >ec��?J\9��g�UD�'Y�Ѱ��[eV�(����]���n?�n�zK["?����^�R4ڄ���h��7�WA�A������mÇ�}�d]<���m��#��;�ȽL#I����\õ�f��1�qq�b�e�Ȫ'đq�S��e#
-'�&J�a˔aHvj��g:[����}�k_����0]5\�/|�x��_����y�FYO���r�x�uZַ{�yj�Fu�N�眿��G�i���_Q��T_��7�8W�����g���v�]=��>�1�3
�Z8���:������N~��eiQ^����p|�<��/~/{�+133��7!�E����q;�6o¥��_��c登��Ba'N;k#��m��v��>�ױ��a|�S�ö��������e(d�J+�I��G�����`gxnu#�	5�Ɏ�e���v��ߋ��r4E��[/����ϨF)~��/Ŗٍ����1,�J���n�NO�׾�5ر�\����]���ۍ١�nD�~fozǻ�ܼw��JK�Ȼ�� ��Ѫ�(`�A/�k���S��GqD�y9&k��"�j�H�4���+�'#L�7`�����;���/���z�4ds��֔�]�y�]������w�@��x�k_���J\s�wp���ik�p�G��FP��W�Vi.��_F�ލC��8�ZX�%p��0�v{�5�������\�uō���1فn�������ô���Qco�/�S����'��ϿQ]w�q'.<{7�K�8�� z����`��ͨ�ut�4��׿	O��_��7ށ3�:��y�D��0}�#EK��Ae��ulk�9x�
�D�j�����<�1t�X�I�d\�h��H�6@��j��im
�� ������c�;����o��ضm�x5�Om�:��--���o{3�x�p�m7�='�h��7s@�t�{��:bx��<	�偅:w]k@� 'S�ud�+?��p��eK`t�߭�1Ҹ��a_Q/&C7_AI���`��D��k�����x�{��v��~���Yt�0�f��3ӱ����Y�{!n�I\ӊh��s�c��qסEl:�t����	P�q��%�fS6���qJc��H:�Ө����,����f0�]�<Ksg��o|O;7�3�M�v�=�ᰂf��5���-"B$.�]`j�N��&�/��K�}K=��y�r�M�v���cv�,���xg����5�c��5����\]j����w{#eW&U����&"1,j lv�y�
9fq���;��$^���?y�><�<l&���{R&�O~�����3p��O��܅�hl�s-q���s=�l٩�}ڋ�	z\���Z��4F9ֲ˖�/�-���,�k�Ĩl6�O�Z^�����*GKv���3 ���WP,����@ܞ��{2�a"����1�s0
U+hLoD� ��c|Э�9�S��uO�3������7p������3���r�lFD�򤯋��"dX��޲i��,�gsl>�ǔc���3v*��2 ��X�{ϋ�*
�6�y�<߄F}�V�Ȉ��+\�^�XԒ�+%��/��������ʗ}�(?o�]����0��ϗ=k�3����_�&����6�1d�;2�sH���/���*Xw�~o���=�����(ĳ47���DUm�D���"�۷Ga��6�R6��&H�@N�K���+b����#l��F0�˄�V�T��KCT�R萄�2�U��A�I�	p�zc��5A-٧�Ȗ�$�F�7��n_d�:��~��ZQa�t�K4�������>��(�jJ�C�"����/�ǣ�0bT: �щ�\���ص+��D���*��ـ��H���I�����7��P�C����C�za)[�g]`�r2�d60E2IZj(��J� M�תW:���"�-��"5Ɔ����x��/�Q:�S�a�G5R8�@��=T�M�1%�y6BK��c�F�#�r�Qd]�,C>��>Eg��{�������6�/�}�����/���G��Ncl�4/�**�S����ˏ��WǄ7b�µBy�	@�b��exGUyXe$�L���=Z��]���I�Mrg,.Á�M�،�j����>��.
C�ue��|��#�+]��/�4x��j\��u4�R<;;�o�TQ�Q�D�<*Z󡛉��T�+���Mm�X		Gz�Xo�E�J��.��A4k#�q�5�֌l�)�S��ƍ;Ā��� ��FT�<�ZA���9����)[i$���/D����&5rZ�w���]FH��MA*�̣��Z���r�X��?F-��lT��zA�ץ��/�m��a,�P�_�M�D&m�hRt��V�����J�ԇ�X_�Z�X���b�|bG��x��P�Ȇr��9��W�`�T�f�`�Ar�C�؆UӟS��)*������u
`_�YZɽ��ĕO���y�]����k��M�[�Z�i��}����l�09�Z=2$�9wؖuQY}�Y�c閁���$\��f��5��O�d�G���Z�v�7�'�v
�?&�X��A*$�_�y�AODbńp������O��Kx��_߱(�p�Q���(�INdc�yi�W��rqn�E-o��D�[�LP1Ru�Yjb.�t������h�4yds��q��ɳ��e���Q��_w��tu���������e�P��5]�7��H��}��nwZ6�A;��Lz)���פ1��8��l�-7�X����UQ�Ia |�%#��%��[W�����w�H�g�`<�q�Rڬ�R:M���ڥ0U��3���v�$�i��d	?w�&�ɯ���'��h;�R���1��͡��.��9�q(����兯����(0q�x�=r(�99Y��T��UqS�*C4�yZ�-ٳE����!R[��[ɺ����}���B��[�Tɠ0H;x�/�,^�a��)Ɲb�.����Rɳ��A)�(�(C�Q�VQ8�l^����pUk.�X�?���\��1�s n���&�ŗK���h�t�f�,D�<��Ύ�J�a�:���@��N!J0�D-)�6�f3E�S�c�&�&���Xψ���������í�G��ޗRO��yZ����EV
ő¡~N8QT8\,��OP���8(I�u.�ٝ��3���P��CA�-1[�㮽�`��I�N4�Q(dÑ�%y�G��h]�@,���᠇��ѣG�e��*�M�L�b^�h�t`�C��nCv�?p�_J8]�I��t3���[������(nc0�x�K��)W�=��Z�'�����:�R��>�w\�s�>�3-�� ���t���Ck�9��[ŧ�������.<ː�s{��+�5�������� �p���D ��j,
�+RGD��5r�O$Z�P�d,��TwǎJ�kj?w<���f�zL�<�w־�Ȁ���نc�{����9d��0�o�:���hk;��:��b#M�30X����VÊ�V�Xa���jk��П@���1+36�����%����-�Xh����;�/�e��j<��y*����V������?O��<q��cœ��P�{����=yc��f|��+��>�7��qC�,�s��H�i<��+����~���ص�¯�ʯ�[�:���:���'xȣ��o���n>�#�UG�%qp�R��e
c+K����Dt���Rz1ˇ�'z�/�Y�Jǡ����!F�mPJl�J�`k�����}����'��]g?Y��D���*�E1�?�����{j�i12E�U�8q��5���,��*�w/�Z�`V���3��*�ܳZ2eZ��D
��]���V6�S̠��`wP���	m����n���,�XJ��p�Vh��(����Đ.;���O:9�bY�O��E�#N�"#5�*t�����^���)��F��"�F�C�5�YNG.�T� �P������J�(,�c�M�h�,�6�l~c�3ч�">��(I��,O2��������'��ۂ�X��o������0l�m����>�)�+[��8<�(Z���D�b?Zn~Z
�k�5��Ȯ+���G�o&��z"͙��h�b����C�s�u�Fb\�
����a�3��^�
���U�ᘞ��+˘��h���G"�5��f;�h��"��s6��\r�$@�h
��	ϣ����A#Y�^QE^o����Bc+�7
����|lj?7P������rI��J��1*;`dń���+\6־8\�y�[G��X��,�l�Ao��O!���`>�����6o�푙�Iv҈gG��Q�1��i�dRb(��AilҖK��D�9��P�b����gU��A��F2Pn����#6��6G�B�8� Oא�;��zD@�%=s����I�D,�sLM70/�e�X�$�"+Q����Y=�0�a-?�+�0��ī��q^Tk
�dN`krĈ�=����r������13<'C�f$��10��^K�w^ V
���=nΘ)F���.f[[1�9�ƝmY��y�|řh��ܠ�	���{8e��^X��dt՚�x�J��h�.Fk*��j
ݩ"@���x�6�T#��Ē�n���.
c"U��r�.A@�������@c2�#@#�/i<�F�yU��pc��-��Cr�1
k������\�%�v���&�=��#�h]�jx^s1�I/UK"������N��W��c.��e@�9 5X'��2P//��ɀXbЮ֓=I->��AqQE�'��իG�⣂̧�2h����&����r��즙Y1X���(j	�"(��l�dCl�{ZG"�K�	H~+�H�ʦB��
Y�D��������r<��eh��6:8(�l��G���|OE4G*Z�뢥�X�B�#l ��h�	R��H�~i�dnR��ж��V�3�%�s
�h5��SLe��ĖA�u���S������A��?1w�e;����QrBC�U��P�ͽ>�M��t^��	XD��\jm�0�C���O�ǣq�mP)�l���"e�������/�,l�[@�w��[��/NS�4 	�>
۸u���Ƭ�:i�Ա����%��IҤU[�z8g�n짶Hz�Rk8,�̉�PC-�Q$�<�����F#Nb?��U�X�{���b�ʭ���"�Qè��+a!L3�>�шvz���4Y�$0�&�2�Yi�JA8�`L�Q^��`Иn4���c��˼b�Ǣ�xlя��v:4�������-[eJ��p��()�?�aV�G9��8v;��	�L�ٕIĞ^�����t|ظ6n�����&�3#~��{x �;{������b;��g<N̪ȃm9���t&R��&M��/ޥj�,��f�^�|g��.A��NG��^�W��"��QPs|�EC�Ӛ~��q0Wk�QUW�8�G��}Ypf+C��(�]�F�-gwU<�@Y���⎒��L�	<���(2�Qs��=�%hb��#t�J�͗�raA4r�UU�WmY*���2Cz$�`��N�}��jr� �p.��Z�X�����8�b�{�����"-���$�h��!��vY���g�� \��?��!�N�[��J��� �L=�Bŀ:p��Y��?�!N:��qAA���E^����YK;����h�m6�_{Z1�^��x �ZZ��6W�2n�bw$�(�X��RO��b�k�"U�Ĵ�@���2��j�mlajX�,(��|��.\��de���%�V�P�3���9-ǤQ���%�F]V�#s��+��$��0S�D��Ȇ����,Z�`h�%-i�V�e��nte��D��-��]&�LŒ�ԵK�=��@]�x�A\���fԛ��W��gd�]���_��p�E�;e��C䨠��` �;�VE\�,��~����@��ކ�:��@�SC������	Y���p��h�� %�!`�
�)E�i�x��³(�,F�h4@�M��G��b�*�R�T���a�̆y��)%	�k�.����}+SQT��)�I�+��"r�����aE(� �b�����Y���xW5�™,�-�}�E�GM������yn��p,�b`���2uG���W��r�����8~�B#��4���ҵ�g+�" ���S�x��A�!�Hu٣IA�h�*6EC��"Ҙ�H[	y�e��scW�cQ�����+�ȃb�?��NTXp��b�G7U�4�IHEJ㙂�x�ުB�����!zWd��"^����(�m퓖ss�V��v�5h��p�H�s<�X�P�8�VܒO.�R扆��}��v�s�X�	wR���,�#^���S-��E�D�]�㸳G�Q�jq99��yD/D�!�4*.���q	߉�J���>H�5��w�r��5��hFa�I,��,6����Q8�\���q�VBd��zRdU�x�$o+p��Oȭ6�xc��:L�h�Ck"�$�S���Ƹ�H;1�SӚ�]�,�f��)dؽW3�|e܁@e�\�(5Tb1[U��bYeq��xz�Z�X�`��!�������$��8�1x$0��դ�Bn�(pVK�\�x��ʻ.�'A��6�=��1���A���Z��x���Z u�:��w�`��f0i�p��5 �K0\�^�����9P}�P��-�;$�6��*v��OML$Z=�~W�c��g�f/aK!G![�@'���{-�	�P�6U��rn��e�B_�q��	j���y���P�3����(B���#1�#CS�C��e�X#�h�t���o\��>J9Z1Ĝ|@*�6�ۊ���-֥�����Eq}�u᫟�\;o#�~g���/��̣-F%#�*8bwt��҇?n�X]fkD�Ϝע�:X�9=����]�>T�9#�N��'�e6�����E�u)�U&��8Tۤ��^-p�-�a��Of��A���"�zMÓ���u��Q�4�џ��M[d�&��C��w��ϽL<��z�i�6��Gj^���1ƪ������%�F�g_��~!ww�Es�K�z'����-���i�]Pm�П����p�Tf�k0;��v��X���,1��-��>KZ���U�Yո`ʅ�X��銊�dK^���5[H[&&��>���_Ʌ���(�R:��}��m�g�]��x�����/GO�d��d�����~
ؾ��6�'��K_{�֩,f^�8���dԣ�j���[O�U/�/^�2�6�@D29�?x&�?�g?�J۩�2��^�y�Lm�Q����_�_��'��h�7 �4q˾%��Wc����jaO�
T�G��5l\�����$��8�A!gK3��M3�X��7����G\����Qk��n�����n�\�+)Vy��5�ח<�I�͙a϶
j��~��E3U#��̆vY�KC�h����2N
�KK���}䪲#1�2����U�`{b=w��k+�B��[� ���Ɠ�������2�F��%i���u�#IG�G���B{%7�S�SF���B%yr�ꮲl@ٖs4*U+$�5e�f����T}��j��e�㗭Ze\a�Q�߿ҋ��%�EVVÛ��f`!���ES��H��9Y�,;���^����=���.������o�#���^��X��_)����7Y��2u�NhT�L�z�/D�����Ci�<3�GPZ�����ל��u���MvT�n�����ǆ�ѝ�Ul�l�dM;�f:�sW�r���5 g���Z6.�U�f�#K��]��xմz�aC����Ov ��x�2f��X�i�/�հ鍜�}a�e�{�uZU^�Ҽ!ih�8��J�G����c��	�����۞�o��o�uzX�R���Fk��+n(0�pƑih{�=HU�+��`<��f�'�2��D��7�B��T�pe�h��,�dWOq�C[��zR�86��j3���� ϗ.zY����.>B4�qBϑGG��*6F��-X�6��\���3B�[Ȉ��s��pe+���ɱ_}G�T|qn)%��I�����-������Ɖ
�FQ�wN����윂�D���V�[�����١s�=_�ڞۄ�s�;�q'(:#V���?V�1֮[-Wb����2ʨZ���{��S�6%��O���y��-7��+��WV��<�Iן�5�IL���;78�����z��qn�iP��լ��<w6�� 'c-�k�v_OC3��3K#>aS���
˝T5���G��u^��aBV _�� ���|p�dJ�C��]c�T0�^�ޙ}s2�K�Ń��3�%�h[�}U�c#!M��B��%���᛺���6��u+�(�	'~V�U��:�*7���=6��;�jh�G��;\�N9�8�}���7��0���bh�Q���|��sN�K��h�u�����l%YTKX�HT���(mP�:��+��݊@�D,a�Yq��F�y�(5�9������w�E�(Z��X��aeO��S�XAUo��uP�;�2��Lk跢���-v�l��e��&4���U%�?Y����Di���r�Qq�,+��,D��!���(�4�oB�r��_�_N�Z~?�/�)U7�I8� ͦ������̿-�<�k�"�]�ܮrH�YK�c�M�����(�)���e�Ga�Y�G�]��I�`��W� ��}�}��4�c��љ�<�w%5�Cd��4�����u���5�m�w��ǳ�����}v�z;�[ Ѭ���q�A������w�,L7�ǐk-�Ά��X��_#��l�(�� ��2���Ώ������P+�+)F}DVMA�Z?����ֻ��*4��i�NT�-�����0���,/���|��~��ZB�G�ח��$'uKqƃL�I�-�rN��1��(��(1�n�[y�z*YD,��r��s~W��Qva�"��h�M�ǲ�w{,�>���Q&����O^��m`��ziM༇�S�*'WY��_23Fc�Mkڊo��U`F��ベ���a2V1Ũ�E;�wؔ��Ga��^�v�Fd�&IZÜO�<`�Yl�A�>&[���� �7����Jo�w��+>�[�N �w�&�<L��������`�s-��U��"i~��!����A.G��,!]Y��΋�}��w11Q�V,�.�(\s".�MD�-=���m��d��jv�{(�й��]t��}'&j��-1��Pv���sx��������!O�
:d#U���b^��ui2�]������%,����2L{U��b���N�aZI�f��o:�_N�������c��ba)JQ�aMI���LU��L6��}�6pE�>����T�0ꃳ*e�����KP��;�X�T�βD�<*a�4�=�������>&����W.�^�%[��ܡ�X�#�*b�,��M���Qf��>��Z�jb���F�{U��Rg��+��=:r�d̪��i�v���}�C���
��+Ǒq� [���̝�'
����U���51���`��2.)�[%���Z�2Y�`1+��P��x k7iCd���o��zݎvw3�Ċv&�<܏G��I�;-�W<�������pYH���1Zǆ+6�0��j�JcF����:D'�jMk+r�īh�^��(o��>ܰ%��z�ݥv������Z�����Im�ͱ�
.mj^����la��\���̚��H���Jh�~���
ƭ�c���G)�f3�1��%pY ��u%�WLElMd2���Z�]����N.�/�5�c�����B�b�l��zl�[��!q�f��'�Y����c��E5d�����HG�?ʞa����i��q?j�]E[x^���X_�f�z�5��|�++����ވ�Y���':�6F�6�[E��EI�(tP[��U�D�S�:�y��n1ºz��e�~��p��K+�L���fD?�J���,�8�N�;;�Z��5|
VY��&�J<�td�
dD���ŝ8��]폰�{���9>+�u��AY�V�W�� Ř���}z~����.0'%�sS5Z��Gꪎ�q��C-2He���E+Vo0ޥ�$�U1�3Pau��XSd+&���4�R��ͬ�5tF�.�b�Vv�6	��T�KSm�]��z\�'��h���h
�E���r�[\��v�-6�&������Mc>֠�Q��EaU�
o���g؊}&�}�7��M(��GG�E���{ޕ�-��mP����y��cj'EiN������a��I3$���@1��tǛ��D��(��'2�$����d�5��U��E�^֘fV��F(N�h0�`Ҩ?R�B��,�Б�Ԙ9ʴ���i��H�LB�S�90ΨA)l6g>�vߎUl�����(�x@D����x�q��H��^}�@��|h;�g��(�[-�T�`XYs��D�xP��U�6�ar���!�O<��� w�"�r4vY���uВ3�a��ݪ��X�����;�&�|�f�1�F�q�s�?�fg��.Y,O��X�^^�X-W��o!�~��J�ɝj�������"�(��v��������]���6��*e���H��]�j��)G
���h���:�*��l��#�0NZ�)n����qF}�"��^����C�*�o5��ׄ@xOfbh@,�O�4ǘm-p%y6Af��k����4L~c��d��Ǉ�K�s�����e]�0��m�L�c�*��c��ǸgF�r&��~��F%6W���^g��k���C��/G��/j�k�5���f�M��ڮ6�Ѱ�Q��B����jL�+rx��
i�Mi���Q�.�gv��|������k0����������Ñ�� s���Y�8@-D��i�X��*J<���:BWk�,k��S��f��G�w0]I13a�]�����Y��k����i[q޹�cv�F\�5���7@�kϾλ���۱Y�%�-Z�1-�G���Pm������hh�r��r��������bBN��x��L����Iy%��Yۨ�	�j��qе�Du�S0�D1ĭ�� RN�I2��3���(��.w�Ot�H%��Ii	�6M��W�;������x�_~����ٴ˱z�^��$���V|������֕"YS���	;/}8n;��-;��Qo�����8��4A�q�iC�D�f%,r�I|j��ʚ�0\�D�7J��v��s�@�F�4��¥;���M8`Ho4*�����KbC]�1�[-5�r1�'
UƑH[�p!�X�V��\s����ѻ��q՛��z�c�
䣞���Y?�0=;��z�x����o����}���O�7~�٧�;8�8m*�-�0�b�����oEy�c�T��Dl����}Ѯ#ͯ����.()���_~��#���O�R����@�*b-%?��Ǎoz�|K`7��JW���Ko�����0�˞�r,UN�(n:��,76�a�y �A(F�ᥡxm�%$�Z����8��}�U��]��k?��wnr���թ��:��=d`�������?�?�����Y��F�L,�50Ԟ��:��&a!������]/8\��ڒb��a|卯uu �6;�|n�1�����bg��KQ�r��-2�H�bB1��kk��,��+������`�\����L�A#Ws�+���D����ȣ~�"saU'��v��tw��O��M�۵ �#���,�1�%�R�0�Z�T0מF֛�L��x��G���6b\=� �c_�_f����8d�����W��w��k��U���/�����Tis�ץ+�TE���@0��s�ծNe왠$���&�Ɓ�:W�}�ӱ{Ǵ�0^D,,.��`��  �:�����u�=ޅ����	��,.��,?|N4����:K'�@!������p��	`dq1���dQt��+�VbɤV�"di��S�aK�ŗ?��x؏?��P!&Vl�),�D�q���B �@ql%��ۿ�CK	���7��]��,|/]W
�}0ֆjE)��������T�Dh5�sS���X�$Y��j�1e�]mn���-.��"���K���˰�T�⚆À� �z�D�S�������+�6���d��,ʩB �F���gl�o������ܪE���Q��~�z-���(&>���!	[M�6y����|�3��~�|�s��O�|/GufZ\�B��x��d"��`y����3���R(�>;�"��W,]$.8��LOOc~~KKK�29<6�Ɏ����D+�Sf;�V��/N s���U��"@�{�^9ƕ��*!�}���1ը���V���w��� 65]<�I5lV�bJ@���G�����Ǩ�V:Ǐ~�ݯ�E>�=�hO��ngQ+��j� u��V����	-�c�!����E*\Wq&4�Yg��Zd0�(���f�]���녣�U����r�\�;vh�Dwq���H�$n,�6���w�]�y�'#ɓc^��lLo����Gr�d�{�5x�c?������Kt��0(�������2~����J��Z͚�W�B1b����ݟ�'<����A��ʱب��*�m�~���qz�y
��%��Y�R����"�B,Sn�ZՐ�Xҹ�D]aR���͊��:�_cȍ�s��W��5>�G�+b�h�'�Q�gq������v��!� ��?"�LLg�~�C��O�5Hn�F4G�i#A>��X��s�A�f�������H�!���~�9x�[���={6�G��2��r�I,��]�ڡ�J�ȴ�g?�Y\��������fu�J!��ح2<��T;��q8��v� �4;3��
9 �L���©��&�����׆;7��׾r�^0���Ƨ��SM|e��(B��G~����\��wź�UMQ9�,��	��6Ÿ��E%GV��U(	��2ţ(�;wlBk�6��zl��n�� �S�����ᅿv\�(Z�%Gk�`��H��SSSG���V��^A��v�: �D�)=��� ���X6��Wr��䓟���k~w��\Th�E����Ck'�# }'ល��O�9S�����¡��е9NqL��ۉ�:���P9�+2*�+����_w��fkZ���x��Ql��b��9���}Pkl��%ફ�£x>�h�ǜMX~F���dn�U:-��^�?��G�B��)_S�щ��s����6X�B +z���y�,;�e	����O�����Xs�ꈰ4KW��qѹ���������%Í\� 1�Xͭu�.X�W��TN���@�	�C�4��G��hvW.�ԯ'FZET�pi �0v��c�_Lj�ȴ����~R��s�?|�׷	�]Y�����]�� ���I?j�8��5�4�fx!e%:��k�������>|<��'�����Õ�������*w��U����"Sm��Ts"��ߍϊP��L4|	��y0��6$*�&]Y�ǔ��=�d8�,C�h8���0N�/��ึ������K��+~�yY��cbpM�h-���ʮ�m��4���F��6+��:�����E[�k���J����1�!(W}]N�Ĵ�ߗ='r��a��@<��n�y6�]8&te�_�n}�(ߺg��-�5�����(��&�U-VV�z�&F{����J��v0��J�ܠ�*�ipj��q�rj�D�+
l��D����PR�zlGDLۂ~�ų�AO�\���Z���+_�v����U�A�3ϣ�+�׌�`��>�[vs%�!�[u�z��~������7��O�w�d��/���<���1�Q����W��f�b��.yG���u7`���jk���MOa�)Ζ&B�+yI�ڥ��k�7y�H"~O���q�Rڷ>C�B�;f��M����;��ٳA�c�Z�i�8Q��]GW�b���v]s�r�s�N÷��C�lQa�hvO�=i��U����%��佒��~����C�B����u���B"5oU/a�ؤ:@�Gx|�T큲L8X������_�7�.����遟�.�r��VL���V���Gj�uUz�
����V^�q�E[��I��k&�F	enS3�J�=����Z�kaLIf��W�����˗���<�"-qb������i�b260�7��e�T�r������k�ť�x(~'ݭ���G���K� ��?V��e�	Q���G#wK�1M4D��9����'��߷�B��/����ԅ�vaf�z��Ny�6��5�e��� �#rC�;���P�� 8v�C&<6nj^�a����q�RBS�#�P��Ʊv���Yl����/��.��C�-�}��a	rd�� %�*�rKN�
�:T���	��S���uo}����@�ܢF0��T�r��T�
7���Ϗ�j]t�3�D3�L��4�n5,?prV���=�N�3�\�	L��iL�X���`���5�̯}�B���i�a��(߻�?~���_���k��!q��(M��f�{Y>ծ��ط <�g��e1ІU_�k|%�Kp)J`�������4��zJ�{����	���7���"�G̘D5�S���D�&=Z�a�QK�ԕ�e��!��߲��������[���������]�e�Y�%-f��n�[��;$첋��Bޗd�v��T&���/�G�����d�ғN��=뻡l�R�"��|��/�%�_��(ƅ���:��`Y��XV��h���k5,f�i�$.�]q�Ȕ~���.6o9�����َ>�����=��.6������o�lR��_��P��U*H}dB�v��`�ⓞ�Bl}�Oc�3ppd�ܲ�D���(���D�f6nV���?Q�梫��̳X�!3�r<uʌ�
�̕GM,�����S99�yX�s ���.���������蒋A����L �/ڍ��QhB���EW��NV�yB�=�]NF�2�����T��E�lۿ����E����^�
��߾NT�����5厐P�C�^�2�z�"�*����"�k�	��?~����#��Jt��R[�PQU�м���G��J�<�����\��G/:y�*K	�(���,�3�0�w��OL��o�t�����b|�w��=J�F��4����"p@��2� d�l�$V	eg���S�5Е�Ui:ɚX�����¹|&(j��/gI��P� �Bԧ6���,pѣ�����7_������YNR�{hb�c1,k>#��g�Q��[�x՛ޅ���7�G��=�OCM�)�$�C�Pu��G��k�,��KAT-X3�P�@�GvnnN4ƒv���ڼĎi /�]�6
ׂ��\�(C�c��p?���v����+��
�R,�Z-h�hX�j-��<`����$b"PRa� �I�"Z�0S�bkD0Y�^���/�S|�u���7_���b�T!b�E��}>4�j��V�/�O^�B�����|����H��1�V����u�@���ص��%䑙"&W��sG:�l�����w{%��6�T�v�T�5V�?����S���:�#��*�\w��!;���Fy�l�CY�Ly���RO�>1���� �Zؤ���#�Fz4�!Y1��.ϡ�
Nc�1:�Q��Hda�"�ڎ��<�E������az7��m��������z��
�ۋ����%������`�9x�o���v��IQ��E"�X�A�K�lP���!�C8��*��`Q!�蛲��Fg]�����P���nʤ��\��{�Ur������Z��f�20��&� ϱ�aB;첱<)�	�յ�-TV�*'k�7.u�|F�?��~���)=;ϊ)<���ɉ�]��F0�"�T��dd�!�HH΅��`���~?�x�q6�x�ȿ�7�x6�����`�i�7ƕZQ,�o]{>��k�;��
8l��p�C�{S{5Y���w_c8�g%܂�Q�Z���"涊��xdvI���'ی�,q���B&�R�,,P�ƐH�]�j!�Ո(�#��ȵ8�e`l6��']��+��8�.�RXUKк�X�ьR���Ri�j��-�"gdC�}�mŰ����k탇(�G�4S�E�eYZ�f����[ο[K��;o����x�k� 3*������Q��坿o����z��6Av�p㐣�	�F�11���L�3�9��xt�8��!c4g��8A\ Q@Y�fiZ��n���������<��}�{o�UTwu���)�����}��>�������Y�S6�$��'7?�=[�Q��n<��@�V���[�K�#:�����X�.:��U��W��V��Z3]y�����r�)1L�}��F�y�ݻ��k���UW����/)x��d�u%�-�j2�8�/�����m|��FB�C��O���9'r+�Я��gj�;�뱃���	����b�1�������/����1�-��Y��Q���*�l<��߉���S����ִ�҅�ƙo�0����f�hh�X�s� �tUL=�#D�n��C�
9@SعR�8eۖ�"�g+�
n����_Q��9����&6]'A�-i`�QIٜ�1�K VYr���L�1m�&Y����O�"�%Gp��,�
���|�T��b�`"<���B1�y��@|!�V��vӱ-����V򒁉 koK�MOs1e2�`GC����K��d�S-R���S�qj����s_KۏW���r��Z��o�a/6�� �<wi~'��71����<�M"��
�JϤ-=�>#�v׫"m�X���|7#Y N���,�(�\-}n���	�DcV�R�`�Lf-�r>5��٘E�O�3SYe�FE[�C~r`���,�?�h�\�˼2�fc��v�1e��z��(J�J�kk�P,Y~�,���
�;��{�4)��/�5��cU�2����b��yM�Z�G�{���C�X�Q7%�.������l��-C�kj�=�^�L-h�-�b�pS��4NҾ5���e^��⏃���1m�8�������tn�
�1�.?,(>�5�S�ȹ_�M`��g;yߴ������b����l
�1Q�߬%cA�e�kMy�Ai�vD&�cx�J��-Y�mtd�X"I�E���x9C���&Β�OC�g��
Lr�q��5�{�հ� bh~	5b�,����H����	Ѧ���b%�ܻm9_O���!d��@��Bƒ�J�f69Y��U�4�
�K$Mc�6-�+��s�֢�U��6���t}�7ѥ�S^�d�X�}�z�6`�َ�	L5yv������\�/;�b����-up��r3������	�Y���B*JS������#!MS?��%�Li:����3iS��&Qm�jV���B�3�vC��3JF�A�p�k�.���h�c�v�L�u��%�,�����T��!&@�31O�l;��a�)�.�>ĝ�:jrjU7��e�l���� 7���+��a���o�
8�*��9G�A�RR�����rt'J{���MN�5��d�#6�ݜ��\a�d�D,�oX��;&I���3g���|>Y ����b�R�W�ТN���|[A�V
d��V�Հ[�+���u�Z2�Cc��:-(�؆�^j�����P3ju7;��6�u��!�ԄWC3a7A���0y�s��	U�0�N2�EExZ�s�����v�VdbҮuqX�{E�|�oh ��CՕp�	&5Q�X��e�f~��U'��z���`
����C�,��g:� �5���{�&��Ս�5��&,bm�h��h%�*)lH߰r��]���\�G��y�ͭ.�\��:�x*�sZO��vsm�@�+j���� �3ϓ�|8�Ψ�E=Nlu��mi��,�ew�|Q����r�)�A�W���%	��+'���k�Y1���]��
=�]�MPP�2�'���H�$���Eiw�Ԃ>hT3	�e7Α]X~f"�f��R
;���H�K^`��.��EK�ƒo��d�99*f��
�Ŭd����&���S-~f��XJ��)�f���Z(����y�٘yNgi��&��{�\ܥ�%	'��_|����ر��^)h;�o�P ITS"�Q��Nd�+MA�X$���b�,xWI��]C&� ����6�����{p��g��֨��/U�5�s���3�����q�a �-v�)}c��5_S;#*�}^4aQi��鉐6Zu�Dk����h���B��<�>��M��T���+rltŪ1����QI@�YO�H�S�/yH�eX�wԖgU$�<��;������d־�\��W�c�J�N�&bKw#���^8�5XV��yY��� �cS��P.�B4B�1d�\�2�RK��I��GP7Mz;�#���G���xg��4���Y*:&�T�B��&})���,'�MY�xj�b����x�ٽ���T��^�Xhf��d磂h���aW��]��y�0��F�#��"�%����a��5Q�IꚲG򋤖��H�%	wD�1������W��b�T[y_"��Si��B���٢���!C��G�g���*ʎ���F�HSi�S���MZ>(����ڬ&_�\6�c֓�4�'GFsF�rX^'�$bW[����N�7�7}�أ�:T.�Y�5	.)��/��7ɸ/bkfy��!,V"ylcnF����kI��`;09n�r�����,(�ʂ��y4��-WV��/��r�䰜"ir`����,�.��9&�����Z_�h2L�6z�&�`��;��P����U1�`��VPk����#aH!''psr�+^ ���9���rbB7gw��U��;6�QW��ب��j��ۗy!CEu�T�33"�r֋�*��k��&����햇ju\ k���1�����/�!y��'�]��T�sZ]y���VQ��\��}�w=fL�[az9Vrh�Mc�%��ИhCu����(:��%���"��u?0AE�x&�M��=���:�
9N�{p��c8�����0|�i���-���<�\l}�)1	c�h�݁sљز�Q�|�|P	�e2j��a��2���� ���5�#��k
�a{W0E�1"��W���k�И�����ĝ�������Gy[f"�ΎB�w�F����ry�蔕(��("X�>���{��`���t��L�,)�;1ʲ�W!��Ƿ�<6!�{��?N<q��.��8�����W����/���-pE �����q�Y���'�C�<���"L�\ds8�2R?Y��XL]����"���)z=�eQ����L�8��g��W����gw��t
.�����(�[������_(��)yE=���k���k��O\��\v��j���D��t��Gb�Ƚ�2��;d�����k�;	����������F���������^�w��7��~��r�;X7���{���{p�+���W��ct����+�a�N��f�&Wk3�~�p��+RS�없Dc4�r���~u�����K��{o�[�r%���3����%B��޻Lͅ��!���YGs��5o&��o
�'��ʳOö;͙��a	#u��h�Q&�TZѶ��M�1ˡkhG�J�d��1���P|����ӂ��������o_{>���?Fm�p�ӣ�n�S!�>4����?˱*��=�c�����m?��-�&&�+�1�u~م�}Er��D[��;�߀��0���"�I�"��B��.������L�;��s��-�:�����!f��{�O�Dy���ˏ�	�굸�~w�8(J�!|����g&����v\��w���l�	ڙ¥g��~�;�\p��w��ߠ��l��s��1��k~�
����}��(.��;V1G���.$QgqGփ`��M�D��y�u�Ȅ5j5��qf�8|j��ȏ��^DZO<��%��wn����>Q��h$f��\��	/74�6[CT}�+���(&6���^3��*:/Ml+q�����σ(����+O��:'���~��9�:���ߎO|�2|��7�L5߸ �07ׄ@̱6u|��:�k�|�F\��Y�M}b�E�g���$��Π$�xσ��o��ٯ�ת�������w���;n=�Qǋ(�R4���U��tF'��\���rΠ�Bn�Q��:/�����]w����β���׏�=덣�W�O㸕�䬔�#��[�S<���8���_�"�H���-y�zm�6[*!����ΐ�jc�R0)�ֵ�v�Gan���D_�,�˱t��S��xIP�`���q�
�:���߉�U���Wn�����������D�4�z�E�4��T�ڢ��N�Pm�ͅI0I�&���#|5<�Z�Q����������.y5zH �h��a`�����ȕjJ�ҳYKIN�Ǟކ�_�U���7q�2fĢ��E^/i8N|�\���,����<�� ���y6�����j;vlǘ�m�=M4��q�ƺNǴ!�ã&�W^7gń��l����<*��J�*�OU�擺Y�p���73!]��O`V���Ę�B�%���7ނ�Gc���R�c����0Z^�����߻_���`ƟϠ]$O$�Q�+�=L�މ�+����4�W�*���FPA^ݖuuOn�!��\��a�9����w��:��ΚXh���v����ג�[y�Xe9L���E`b:��RQcIGb,�%Nn=��X���[(���"�ڻ�ֹ8�k�u�n��|5pꩯŽ��BvbGk'�]�m[6c�3L��p��ER��KLy��Zr���u�8�4tF?���X�UJ����b�ú��bӶ]芠޽���J���VKZ%����v��ǛE��
8&&�"���|^�g�h�����q�[~�ݹ˦��"u�%=6@��v~35������;��4�7=���j5yt��wc�Np�l-��gZTc���o^��7�{����X�Z0�Zq�H�\��xP_�Xr�Ĵ��m�,��a�7%�r<&f�f��L�?�p���l3�Yg�ؽ��!^�oz��}'`�ګ�G,�+.��>�"�>|9N���e�0GrX�k�i����Z�ZH��t�n	���؃�}�
��0�v�Jƕ>�NΥ�	f�9Y����u_��?��I&�g9�¹��A]>�����o�����;Q�2b�#u�G�֘�1+G�H\�T��b~7�|>��_·nK46N
��]�㲋�����n��j/��W��y�w��O\���x+yR4�tξw��\���%\�\�Șah
�֓��6BKH�J�,z�����|6?��y��V��A�����<��^��?݅��;kN�㺯��]�?
�z�L�|� �;�߅�b�TG&ЊM!�U��N
�ɍd�c|r~p�#��&�]y�&��]�ɗ��^�-�o����L 	J(M��O}�Q�Ys<vEں{�z�$������	<��^�i��V�1���em��h��h����Mw��-<���P[G�-�?���pʩ'�7 ��~��=�1���?�c�uڙ8���`/1oxRۓ�z~+J�1,�^X�8�Y)_�c�0�����J�7[������U�}���Ҡ
�6nA�H�}�I��ûerD]�{<Y�T&��z�V�{�"Z"��<}�����N�yL2-�X�t#Gf����t�FmǊC��ZA��06=�F�m���y��&�{�!�6b�����>�r�iN4LՕ'
0���P��N/��61���c��0��Ąn������ڔ7j��ʽtEM<�m/���S�L!V�	�� (O`J��]?} w���L;�ȊI89G�[���s�a�B�n��b���J=�.*�5��07�f�&�Lݣ�95I������SutR��YdS��Y���4�b�QlZy���8x�X]�ZH�E����f�V��� M�_!3�=�Ֆ�ntM9�b`�R����{O���k�e�6�aƕ��[BI*5yF�¸��W�8��mkg$Zn�$���wCK��_�Gb�n�BQ*�I6�6�r~(����n�����8>����2Bȸ���TC�j�m���fՙ,�/�P�%��[��$Yu_A$���j��9e5z��:���lƒ��<p0�O�g���fFj}v�����hn�>r�os:L�j ,�,#�VEw~���S7�8��s1XRijK�L��.��[(��+�6���8�9I��+Ô�P����@��*�дgBNfڇ�R*[�]	�ѫ+IM	�YN��k�H̸dȘD��A�f�w`��v;�?D&}/���6|�,1]1m+%��wuA�W��>��,:� �.�9r%���P��"*xn�/0ĲH�%�i����3YעB���1�"_Y/X�i-ñ���Nb�gW+�px4:ME:i��r�C�%�]�ˑR�g����4-k�|6���AH�� MFnv����L'1�_o5ܒ�0^��q�E�1̙��>����%�D X�����m,??���n�G1/��4�5��}�}���[��(�=���0��~ـ����I�Ք:h�<jXGܙ��_�N��=�S=6`cv�y>���{�s�[�����g�M���Y�L�C���Z�GuxT3��-:bAl�n4�I�T��w�ƈzi�� 2ZG�3FA�^]�����_Y#k_���Y��K��Bh�E%�d�%˲���~��k����U�@�ڲh�bT��G2�)CLb;�?��ɩŶ�,�~i<3V���|��	5�[�N��~��:�X <2��,\ʉ�x2��vD>�P�F<��M��^̳F��l�'X�7�XԀ�G��K��YMg��؆S3�dwT�t���|�������}��2{� ��^��J�wy�PALu&�v�Y��ǒ��,�a�t��J�����f�h��ҋ�9�\D3��i󖬒l@�M�`
۪UK����/�ݬ�Yi��l�T�~��lz��m:T�k5�,�\�[�[�i�X�	��y�ġD��L_��L&��TL��M��fǓ&A��ep=��\7�f��$j7�a�Sd�Q�PP�D$$E�m���C����󥏃���1�ť���c֏r"S�?���5�f[i�>;0˫c��E���O��n�8����3� K��h�2��Dq����[�J3h��.8Øb߮:�l����P��hE[�0Ɏ��T���5�A0�\�J~_Mc3����J*3�=����Ũ�v���Psj�\�T�Y'jj��tvvZ��e�Y�+�0$p��.c,�����݁ߘ���R�BFJ�M�S��I-m�vc��u��j�|l�8��i�]*U�7baP�n�,VÑ]W�(��:äh�h'�����I\[39�HLN��&GՋ\<ϵ)�L��h���	]�^�B�ߑ���g����#U$Z����=�1C��Sj�����g�7�I=F/����� s5us�����"�֎��쎒PkRY�C"�?��ۊ�]m�j&��x��<�Y�K�+:U���k�t��f�f��,C��5���c�%L�%���Tr�^ʤ�G'He����v��R{�� c#Qqj��z��w��ۨ�b�G�I7����`�E��8�'aI(�t�~�i����1��uy�jf�.���jO[f�����D�܍Z�wш�9����~Cch�]��fn�5�Pt�&�DU{����/�FzS�jo_�s�xz��tP��Ư�g�!���j��p��?�-O>e�J���e�%�ݘ�1��4�3�d���Z��\DzL2�~���$��a�Y\��s�n|�~�j�l��Ŗ���0��B�%�ϬtP�{te�eT^�bM(ܱS�����SN�\'���$J�1l+δۄ��4=]t���B��	�X�UC,&��f{�+VL`�ʕ(TC%Jcy`�e"������ڂ9���V�1��;�Be���W��>
f���n��L�g�Zt�E�C�d��I�Z�Ƥ��zH��q��VKwp�
�U{f"�l�TK��0u{�ڤ�1j��hʢT��-|25nd-�)��U��wH��1?0�5��G�O�n��<׀�N�!ɉ��P��R!w�[�$�J���!��APNv����Z�S��	v*��FC�ZM�����[��<l�!A�K#�9,<��A�M�7Z���o��p�f�W�>��
Z�϶��rrg ��)=�CH��}�J�{B��s��'iڗM�jm>�(�M��e掺I���	��YE���ؚ٬՞�<K|;}W׿�wA�"��Ts�m�=ǦO:�ݲ���B�S��jwǦ⩊�S� �-��p,ڎ`�PS���L*;�\Em}v,�r����N��_�l�Z� �g������ɤ�ϜI�`�g�zb,&�Ȗ���v���G2�ˬ�h@S��3<���1�*Y2S�Q�iE΀X��Ƭ�����hu{~�Á2<o!�J�@��]���=�6�<ƞɈlNbx*L�(GU)���Sx�hV��v_���a�}��n���ps�0K%����K�kL>�)2��*�%bIP�źP>V���׷�%��d�Y}��\���U.>���YI���j5EӸ�T�U�`9fU~��'8i��4ѡ5e��quc��D���$Y�Q��f����4�~^F=f�˘m� ��1�	���`Ǟ��9L�U�]M��,SW�)m`�bH�*�}z��2�s�d8����KQ|��U��٨��R�\*��@�VIg�"���)���xP&Z�`�I�Q�X޳���S�@��ݘ�������A��C�=�m:��i�����g]�f$ڔt�8gI�.�(a�gԣht���he(��j
z��,S����������ʨ'��MicS�d"Q���A1fيI�P��pkʱY��H�-dHk"�Qά���f�i�bF{e�:�b�ٽ����1��Z���O~.��mHfg�b��"[7c�.R4t�PvB�S���gFN,���4��FMP&�K
��{��4r�u��{�9�t�qfy}qT�gO�56|����~g>�g�����=���
��bQn�>�@�'�t�5�fo6��o�Y�)�\s�k�m�d ��G��f )`B���S���ȏ
���=�B��i��a"�@�0--w)IV�jg��0��3-4Km�je=B���d^[	Oש�B�u�NS�V��
Y]�$0�����ޖ����2�$0:r#�Ly��b�fy���p�H�e=�M��3t�Y� �D6Dq��
�m�HyRR�Fj�����ܘV�i�΁����P�ˏ��t�m	�����)���!i�l9H��OTS�-�Z����I���+5�:cΣ�.Q�����NK&�.�2��_��+�{�pjd��[��\�<fe#EE>��06���רFI��@vl��x~>�D }8�y>'���b�_������J_�fTE ���$,������Q]�mnik�x5�g�@ǩjL�����S�F�l�+j�԰�e~�����*�[Q���\D�*������{�pN�4�:ن<��X��.�U��@,'1��b�9%�˫А��jH�|�Y�c���g��� G��`��t3�4_�$�4�i�D3M�}%�=��E�@D�1fs�����	ztݢ��rSC���RfB�D d��_�
x�����j�tt�o��;��m,]o>6�GY����x,�NytT�挋5|m���pJU�Ϻ�cȻ��E�p�Eb%lD�Qv�f;%��2�8�o)��9���N�xEF6Mb:�XFY�܀����9;���Q��M8$J���&|��;�"��l�*�\���Z~�d��d�A���1�;����_�����j]�p.��e,'����Q��I�I���D)[)�4/�-:2�,��r�Y"V���7,s"�*�zu���� 8���u%{N�k�
�d��'M�O��f&����۠)Hb�VB�9�T�ihW�*h�A�(���ޥ֘�?���$�+0�6!/!���`w欦�65�ɓ�yyͼɵ�^(�/C*|Ij2�� d���u���NL��TK�r��Ӂl$�.�3���0f�%�R�JD�%���s0&���G`�,��؀%�z&3o#G�5�-�:(��+g��/+/k/�'�0ǡ(�f^�C����k�(w=8��7�'��Kר��-��p�Zu+k��t"s�U��O�AG@n>ߑ�5���"��vC��	��0A&(1�SqR�������f��O6�Y�T�+�u���ԛ@�SG�K����䞺ih�H�^W⩮�0W혓�(X�A���`�.8�RDCE6M�`�]�-^�G�rd:6�L�w�ɵ檓�I2_ej�2�s�r�5��h�S+�y*0C��ɤ���b��b��Uu�%a����[�=E�u�[�9����u c8j���cCs4���|�/��#�8$d�]4SB����=�;m�}B�{�N�i�`�+���Hh8��	4��8�<�иè�e�ш-���X7��	-'�̙�Yģ�ڋͳK��Ԉ�蘒��`Q�}���ibx�X	mG1	���E^o���3�Q�T:�}��"['��,�����Q�nhh��:�M�I@�fV�(��\��ȘoZ��(�{��q]ߓ#�����6�v����5�FNO(H����b���z"���Wa$ECО��B�]��X)��2�<�ג�9����O3�f7҉ɸS=]k"g�+M���?��S��(3a$Z����d�b����	f{�q'	�'uc�IO��H9@�U���J��.`d	�����O�V&b1@�s�`tc�\7�ϹCb�9i�T�Փ�CS�x�ߡh��Wn^�"Q��y?�Ė/jy�Q��p�-TGdG5v��D���f�i�b�;���9Vx�DF!���5NJDǸߍ��|�:��sI.g�.�0B��F��]Y�Ey�1�gŁ��j<�q��0����h��>�h̲mu�K�����{�%��A�a��e��1���T�݊�ĵj��YBN{'	،v� 	��ߗ�):�޿c��C���׼t^��r<G= ����~�|�=��m�[��"�yG�۠�.�Fԏga �!���W=��:k��� ��Ҵi�E�p.�̟x�BŐ��ۋ�ʊ������H� I㚝h�b#�^'�B��=O��@OuQҸ�=H��5�����������S�v����Ǣt
�>Wұ�fKE��g�G=���C��Tk0�<���v|�ǳ�Ug|��z�0�[q���\vT>�|Of�4~��|+V3��h1�Ӗ�Ԛ����
�o�ƻ7�MC�9\ks3N�&?��������a�El�LD����az�?�隴��/��;�FF�l6���O����?�p]o�k;w<�X�Vav��7O�����-��M���շ�cc��x�ٍ#pm���6�s�|�������_L��%�\	�\��_�η�������������߽`>Ƶ���^��7,w�,������۱�T������9�\p�,�а��r���߿�'����ј]h+���^�����6��f�v}����N��/�(�l�Y�c9��P�0�(��8��_��:Ђ�a�S]�k�A9�ꄫ
��rX��2/?����A��D�B�GqS����Ǳ��)�1Q��e�x��I	,B�l�Q����c�ޘ(V�rf7��/F6��wʬ���֬Amz�����n{E��n�y��W�57s<�q�K�D�^�Hշ��q�qL	F�T^YL;�3�U2����ɏ_��|w(_*�_��bg�b�8�4ʗ
y��d�/�(�cJ0:����8��b���0q\vC�>�sD�'�v$ʣ�>����e{�cJ0d��O��xK'�\�p�z��ue�JQ��'ը��7��q�	�<��4M�M0r�eJ���/����a��A��˭��֣z�k�����Gl$��KO�^�؟�`���8�#]47�aG{.�0KGq�ɘ7D�� ?�C�����R1����O?�`��w�r.�����V����hjO�G���ڗ��Xf�8��_�c �l� ;vY����L	�Qǔ`�_i����r^�c�1��U20����5�����܂1o-^��c�s}�Dq/}$Ird,|��_��1O0�Y��s]�h/����e�d`̋O,��V�����Q�,�bj�Ʋ�ǔ`d~Vl��5�?D�Aļ&��I��|�M������Q���.'���(��m3�	�V����jy�Ϝ#��.�qL	F�[fa��o��,H��lCCCڈ��l.[ȟ�����5���pS�Q(��Z�P4E�NҞ庶��z��Uv�zY��-��2��cC�,��]�V��Qǔ`\|�ş���V��eq��1{�r]���/���۷�#BY��7��n,���K�X���T�3r�8���6�o����q�eU���8Jc�ڵO�ǔ`d�h��c��W���3j�    IEND�B`�PK
     8p�[�c��f  �f  /   images/c88b2895-5e8b-4a57-9f9a-b80dd50058b1.png�PNG

   IHDR  �  �   ��ߊ  TiCCPICC Profile  x�c``RI,(�aa``��+)
rwR���R`����b
����>@%0|����/��:%5�I�^��b��Ջ�D������d ��S��JS�l����):
Ȟb�C�@�$�XMH�3�}�VH�H�����IBOGbC�n��ₜ�J� c���Ԋ�_PY���Q���Tϼd=#CsP�CT�%���X�}�����ߍ�������k'BLÂ�A�����΂ĢD�33��10|Z����� |�'�8��,������z����j��N��������.j���p  !e�2���   	pHYs  %  %IR$�   xeXIfII*            (           J       R   i�    Z       %     %      �    o  �           a���  �zTXtRaw profile type icc  x��S[n�0��)z^�8~$R��b;^eW�J�ё"�@`H�n-|DI�D��@ȴ�v=L�"�	�s,`�ۮ��z����"H����pz����3�ͬ,9&�h'�tN9#���(���d>CQ�h�|q�k��R�R����mOi�q�6�Z�ܶ=���C�>hrK$>���U`�͚t3�s;����%�S�T�c��\���~�y§b�_"%�G"a=}J�H����|)�Ni����2��yl�c���r�E��|�7$��8��s���.PJ����
��wq�8��P'��j����[ܞ�c2����g�+��|����RM�=�c2gҥl��ϞauTh���҈�\�z���줡㜥   %tEXtdate:create 2020-01-31T21:31:09+00:00��y{   %tEXtdate:modify 2020-01-31T21:31:00+00:00	�   tEXtexif:ExifOffset 90Y�ޛ   tEXtexif:PixelXDimension 1391c�   tEXtexif:PixelYDimension 800�요   (tEXticc:copyright Copyright Apple Inc., 2017���   tEXticc:description Display P3�y��  a�IDATx���|SU���M�M��ޣ {��Dq�����~�V*�~���(���(�"{�Q6-�-�M�{�'I�M������K��{onn���cU{�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!@��-[a츱�aC�5?�q8�^ݺ"���0�
�"���l�a���>C��p���Oo��vn����"��mE�9F�1\���?ۛ�����(:���c�X���_wlP(�ʔ{���=��|+��#}�Y��mo�w��k��]�o�������?�O�0�?���'�Q���W?s��3��"Sڶo�dՊ�}�I���i�f����gf^�t8Z������^d�g`���>�n�q�0K���k|=Ϗ���5�1��}���I0�p]�y��U��'3r��~'_{���G���ߢ��h������1o��v�#�����޵{�I��z�}Պ�ged��x0'""��!;;�߁�������t8�ADDDՎ��4���N����E�l4"""��L�����QQ���ԿTP�UK���	���sn������BDDDՓ}����{�������H/�=��|!'""�c�4a��sh׮ݔ�#F���u�}�?_+.q��p8PPP��o�O���m+�p���DDDG�}ǎ툯0;+k����C���PA܉��\��+z��I#<r䑓�\y���O5�Q�?�^D��R]�]R<�5k����q֦=11Q�s�*Yǖ�Ull,���0�C�Y6'"�`V|֠g�HKKS�o����T���Ύr���������GXd$���(T�:����=3+Y*��D�~2+3K��H�h#"���sx���_����`:͈�����O��;r��"""
f����6.��p�)�ggg��oDDD�����R�7Mgx�'�����"""
n�Cii����p:M{�'��]��QP3��SSѼE�8���,�3�:gOݟ�F��:�������y�
�DDD���";+;ơzI2�kff&���(��j����H�4�L��at""�`&��:���K@/3�^�a�Љ����nC����E��J膻��0���(���*w�^���(@VV���(���*����:��D^^>���(����p�Yo`� ��;w@/;�����FDDD�Mr�0��mPP�ϵЉ����iB��'ԭiՆ.������Q�V�%""�Qt/w���^J�&�΀NDD����m6È𶁴�{+�Qp�/^�T���t""��g߾m�*���6�Q𲧤�H������]��1�'���i��*w""��g����m*`��r���/��Ä�m�����NDD���3��G@g�;Q�S%�Æ����˝��(��3�����G����ΐNDD�Lس23��i�I��S��)U�ge���'{�3{NN�
����%�;Ճ������zdDD�i��K�DDDA�T=&&Ff��Н*�;Y�NDD�L{xD�t�S�:M�~Q��l6;|T�;�&L�Љ����=L��*w�Su"""
^v�a�ax�&�܉�����0�QN	�U�DDDA�T�\J�׉e���U�DDD��.K�|tV�3�|�i�̽t�U�DDDA��%���F��8tV��rK��U�DDDǀ�����t�K���˝��(���K�z���X���(��E�{	��7���t�,��ʝ��(�ٝO	�:��:űʝ��(hI����4�r��YB'""
fv��a�iz	�n?7�)���(�ٝ�sm��NDD��r���SQ�n��^�n��GDD�쐕�L��T07Љ����)U�J8|�r�Nq�DDDA�n+/�K�g@����<����@=?""�F��0;�*��乸ҵ033ii��k�.$'�@jj*>�����9	�QQ��S�ѨQC4k��6���\���1%>�|��%rpq��+�*3��?V�Y�?���Eb��-طo/<���<W�C=��,|��\`�!6&u��C�V�ЫWO0 }��A�&�f�1�Qȑ��i[�I@���p�{�W�܌���X�z5���;�:��V�ޯJ��(��Q�w�{�>)ͧ�Ė���/s0i�$t8�#�=�\|���ܹ��v��D$<�����pU���Ʉi7`��r��s�C��\�U�^�x1�����n�n٬��E�ۆ�)����`�E���Oq��W���GR���yv"��\�g.~��w|��g���;п_?�i`7нN��¹�}�\�-[�b����Gcǎ�p�W�����=轢������i�O��P\p���������O���u����拓�'�S��o�T!����>���2>�͘����3������_��p���T�Y���tf������ذq#��nԉ�cP'��'������ix뭷�|�2]�Y�^�z���'��2���V�{!�Pz^�0���*RS�µ��Gݷg��g'a��Mw���������{���#R�۟���#G���x䑇Ѡ~}u"
Zy���7o&��f͚���8��yHo���;�1��&��ޔ�y~&M�\�f��`�
���hܸZ�h�:�E˖z8Z�*UGGG#7'�z8ۆ�n�:lݲU�TU�[�Z�QV�a����HOKǨQ#� 1�A������K�,��߁�����Qi�tn��lC�C�����g�><����!??�oF׵kԸ1����3���&M��v�ڈ�{o���b�ʕ�a�:�~�:w���Gf ?/~�$��'�@LT�:�Ca�^��,���eʐ�0���or�gf��_�G*��`���9Q'>�>n��V=��v�Z�ϖ�|/C:�5i�H?�~n��L�<S>�\��S�5��s���[h׮n��z�~Y�(�2+&K�"��n�f9U��W\�Á�U	x���s���Űa�p�9�v\-�_+Ƴ�L�׭Kg�;��|2��֮�ù�J������ѱc�ؿ?K�DD!Nt�s����!�{Μ_���~�2�M�!����#г[7�_+O���/�	u�b��aX�l)�36�6��ѥK�� "�P�c�i7���*w]-̀^�n�ꫯb�d�z��L����p�Wb���hռy�Kƞ��u�@����~�H޶�����{�	�_xK�DD!ɕ�۝�i���q����0��)���_Q����p�����FTI0/N�}�Yg�����ǟ@���(�/3p�@*�y�m�4` ��cP'"
9�����rg��#���,F�9Y�.;ѵ[�G�M�VG%p��,2����/�L񲕁?���?���%]""
I�L�곛�k�Ԛ]B����i_c�jo��L������ރ^=z�R�'�N݃~�os�o�X��3��0s�L�{�DFDT��y�"X�X���x�����X]��:Ne��.��� ״������͞�}���[8�2{�u@|�ٸ��K�ɲ'8�w�{���O��������m=�c���xbP�p�ٟrss�����f��u&"B=�ߞ��y�v����y���Cn^���OV}���a+���N�[�8r��!�1�(ǲ��V�Nq�|����EFxȹʵ)p�>[u�rm��ץ���u}]�����OC��:����9�?���"��\}��ˌ���^��Пc�{�hU��)}>޶�R�5RT�y�s�C~J�@~�V�,�[9C�����57"��_@��U�?ϙ��+V�ۭ%cͯ��zԍ�?�7�/&:�^v	�M��C�0���-lطo�-_���Y"v���X�vV�Y��6`��]f��S�P�,�B�Z�ШQ#�n��:u�q�uD�����JZF233��]ۺ		:�*�>��)�f���X�x֩��s�N�I�##"�{hѲ:v�^�{����k�}^ŏ�r�*,Z�k�5۵k���t@����36o��{�@��]о];Ԋ�����u�8��W�3K��t�	�H��r��!���Q�X������u���lչ5m��}ջW/���u�9��a��5X�p�>Ύ;�q$C�����M�4E��ѭ[7$%��k U��{2��3-=[�l�K!�9n۶�))�����C��(�OL�3A��E�ΝѦMk�V���~�:��.�����MIJ�)���+T���6mB�>y��zK�D��f͛��,�u���㐘X��ZT��gVvv���}<p����_�X�����)�T��21g�(��t���k�8t�(���S_om�&���O<�R�>}�]}�������֊����m����ޭ{w�P��螛�J|���f̘����[�nEzz�����u^��t ���x�s�98��S�P%���w���x���٧��U8r%���5l�/��2ڵiS���C�o������
+T�g��>އ�";4h����õ�^�A�����8;U��n�����/�l�2���w/�k����(u�p�)����N>�$�R�ؑ^�/���<iR��r]d��_��*Hz����ᇙ��/�x�b��>>_�͎z�����5�\�s�g[O��J��`��F�ܰdrd�$���q�#T�T�9���u�	�$xUU��\�M���5�'���X�d����Hp�uT�.�6P�]O�ё"��*�W6�{�U�~1#G�ҁ�0��j�L�#�<Rbd�<������ս>Uw�MNNF���zoR����Z�.�1�sp��#�}{���� ���'��o��H׌2*��ґ��,X6�����?��v��#����.�С�)��^��C�`�l�R������;�ޱ�A.ǭ���*�4h�=z�K1�tP���>��U�ɫ3U[����{����z�g����t��.��c�JXd:ܛo�Y�ʮ'� ��%�ϕ�X��$�9[�
y���N��r��z�8�ޭ2�|��~��^v)U�gR�ve�]�b���ٳ����:���q�*w{�6|���0�Ǚ�Zɇ�J�͎��T%���_��u���<�+�ȿ����_�sGvv�_�+�lʾ��5�����y��ǟxݺv-���I�����B��Z�'_�.w�ځi_}�9?��ŗ\��{I����'g�k�|���z9ϕ+W�i���-�����nՏg�T���p�������KGb�*����?�{���K���Uk���̾R�����'[[��>'�dIAa����G��o֙)��L��M�����Z[j�֬^�u��T&��ge�ԯ���(g�pKU0߽[� �=�%~�q�I�������5�گ�GZ����[=�m؀�^{��9N;{$�6%������/�E]�r�Z����5�m��֩��,ǘz� ^U��7����}(���\�;=���}lٲ�����]J������7'��^��=�ܯ��5sm�?5o���ά���:v���)푆V*4u��p����N����|���f�?c�u�!�_L�[�n����|��"�>� /���]ŏ��VJx�n�\��cǢo�^��r&�9�UeXe�sU�-//��<{s][ɠIFsŊ�駟�裏�_����2��-�S�-��⟩��]x��gT@��&��̊ٵ�̮Z��?���H,���>��I����6��x���r�#����D�Х�2���>���:wB��m�Ӗ���[*J>�9*Q{z���믿�^�)��2�J(2���ч�R�J�H<�!C�v'T�%���'�x����d�k����~����@?���B����3�{5j��4dee��2?E�q80��oUf-�Ox�<�$�*�9
o��ffT�|ſ���Gzo�3�up��8���J�/�_R���>������O���$}�+S%57�F���Ƕ-��f�x��r��0��iذ~=�}�\tᅺ�_�SXO���/�£�<Zl�)��m[6]��������۶n�NjA@�����:lM.��t�t�2[�зO�׉�:�\jf���C����໻����m���WJ�Y��d��bX�w��_�h!��^�����_���*ڋ�	Z�1�w����a�B^���t|߁�'U
�4q�Q��-,���1a�J�=U�9�����NJ��= �r]���1��W0��	�ζʼ�������yx�����K/�Nco��^;i(��?��@���u�ȑ#�h�#!����F����9�[f��zH��������|���ū��s��z�
���zg㪫�
�gYڌ�3K�b�c���+�������Ǚ?⥗�cܸ�������eR:����ǝ�Tk��g��Ѝ�bz͹xť��`Ϟ�^����B�.]t5o(]!OR4��Y:t6o� ��ê ^�~��8ӻw4k�u���UT�h��]z���˖��]	��=gö����Ï�k{�E��T�ק�~��%���#"Ѵi3�B]Su���7';�R��Ҕ�n���VS�JЎ||�ɧ8���|�
_/�]	hLl��h��m�"11QG����uo�;v�;�Yg|�T�H��E_�.�W����=u�4LU%9W{y���D�=M�4Vץ�>o�$��RSS�a�l޴I��[_W�2L�:_r�
��0�L0w]���u�4G����u��n2�Jz��]�V]�dx_�X����(��N8�_�������ȑ��v� ���N��B��I��K�.�3�����Qڵ7oެ۶�'|��C�.Fq6=���=�;�^�I�$��t�2L�<����\ރ|O۴i�{�K�HG�C��r�򹦧�y9w��LӁ��}s���c��A>�G���}��/��\=�7mܨ�[�d��%�ף�t�S�֭[6+��)s���2>�����ak2�H!�ک��H 5��_�|9�?5��`�Db���T%�W^y��#פtu���ԗW��M�:����k�Nx�;�oÓO<�F�h�8Ce�Ru tu�+
�R��ۯ/���J�v�ih�����̈;)q�P�9����oM�R�1�f�Ϟ{n֫���]7�
�u0��3p�:N�޽Ѥq#=��s9���6�k\�����}{���#Ìf��:��^��"�>R�s�v.
�a*A�ޣ7�P���[�j�;W���W�dΤcۤI�����e�	�34t�x̘�طgRS���v":�N9�\}�U�qӦMu	�s]dH�֭��ݷ�����W`���"C�O���}zW����3�ǘ����yp'��o�駝����,���!�1�S��߅�����Y�,2K�s�{]VN����y"����}��ΕΠի� g�u&.��b=�q�ƺ7���zA~>RTfm��%�����H�Qِ�o�}�]�pB=����m곸��{p�-7���]���;u������gj��Q#1��u?�Lɐİ��?��kf@�R�+���D6Х�P������*p_Ub'�|*~�a�q�@Ĩ���'9��x��W�������6g�l��X��mX�z%�W	�۪�Ѩa�J't�P�\��T%���;q뭷��JPQ�L�p))�҅<������>V��t�Q%�����[���x��Gq�E��P��8R"�ݳ�w�'��?��*SeyUR��N�m\�а�8T`�*�G��"�*�ȃ�Եi�Jp�+c�\��-[��u-q�
�R��
�e��B�u��l�kޢ�=4LW97�_��K�jת���ҹ���N�ñ��?��IUb���{�͚4���^֬߀ѣ�ww����'�n��s�mh�2c��:��&������Izʿ8�E/�(ٰr�r�S�O|�Mԫ�P�{]�냅�Q������O�Ї���멈s�m�y2��|�q��aʔ)5r�:�����$C�j�9��nE�Bf��Gq��Յ���2����4��>A�I	��zg�'�q��ϬH�Zž�b���u���1}��qc�}˻C<��&g<�[��c�=�i_M��8B�)�|�ɧx���T�V�6j�Q�G��7�Ꜽ���R%����믿�vxz���T��^��K�DwZ�VaoǑ`0d�`]���۱g�.��lܸIWG׫�$.֊�K|ݺ��8����I����[Ǥ$<���X�n}���H&�ƽ8�{��1ͅ-���?U�1c���nƖ�-�c`��d=#�t���a�ĉX��[�թJ��1b�H]����ɞ�V_]O�II��V�	V��3f`�*9ߦ2��Q��J��u�_��T�3�9?o��!�Ho��]Z��~oSKK��|��:��^��X锸��Zzj|j^�9bz.w��멚�)N:rI��+�['P2�HL%&�6�i�ܵ��.2K5�u7p� =L+�]�#z�����J��t5���H{�|�ǨK/��\gW{�C���]����ݯl'��I�ᤷ�*wk�.=��`^ѡ���:^t�:�D�g=6X�z�J�+��;�w�q��ů"ץW������1F�t}��H�[O<�.8�����{��N��T`�>��C�aݺu8EmW���]���-��V�e��O>����+0��g���L{����t�{�+6��hˬ��z(��g֥〥)�|��a�葅����h*�I��K/�K�,յVs�H��c��	�N���Ց]���g��m�vM_d�p/SfVWs~��ŋ�[0�j��숃���V�ǞxLw[�'�([)�l~��ttx�� u��8��tӍ�ڸ��A�L�������mE��ύ7݄s�����9IIpР���O�x���1t�=iK'��֝�RʖL�ۓ�Fj�>x���J\~�e>k,���*�O�4��C("7JG+����S�#S�Ju�Ν�U���|�M�A�n+̋�Ƌ/�Pw}a����$C}��1�����Nt�p�Zb���W^#�j�G�)S�m�U��y�f�?p $k,��Ͱ�۳�&��KG���l[�V��P�i)��~��7�Y��~i�'�T.��SN�|;�����}�}�a���k�������s7�p�n���qM=%�u�]W���:w�&M���`��G'Z�l��.��2:$�~b}��f���A]�&"#�����)�Oj�V�Z�:�y�xm�>C�u�Ǒ���w�5)P����蒤�NS�*	����2��:wŭ�ݪ�D��.���o���f��.�+K��e:��^�\���0��$��a�k׮���B�{��]��Cꚻ:�ѱbJ��M&a.GMkC�_:Qe����B�+�ۄ�y���$\q���L��OI�.��=��?�:�X�b��5hr�9�<����uĀJ�엨J;�u@_�u�SO;�U��� �p��z���L��U-��V�[a���+���ؼE/S|��s��ǣg��*�JB����m�uQ��^�s��Uj+�2�aa�ͼC��z\�ަuk�{޹z� ��ҿ�.�M���[�5h�Hw@�L�kO@�*yw��	�M�n����̬��б�>k��]/�jb�db��[J�6�`�=D���3�:�[�
h��Kz��w�y�c�UU����0�!�^}UB)=g+P"UF�a��^����r�#��.N����72C��- �>=z�@�J���u��$��ye�лO�J��/���KH��uY�C:�z��(���3o�<����^v��F���,u��x�	i�8p &�5�G��ۇ*�"�Kf�c����(�;YAN'���*s��"1tL�v���u9�����M�>f��ܵL�*�W�L�b���:2ɔ���B�F�4i}�7\�c,XY�K�}9���B:]�t��{��_�׶BSO��1 �Ԇ���qb�>/A+�g��IV�mV�5�ef�U������U+Cw2S׿V-�m��zQ_v�ك��Vx}�k�nh߾j�Hr7M<����J&ϑ9�s�n��^r�ש�������"B���VMcNgH��Ւ����yU��n��sTt�ϭ$G*������٧�`)Î��z�Y���j��ڷw���n٪�l.=����� �+KWT��{�ԓ�4k��e�����H:�1u"ݮ]�J��}]t3���A�?�l��%ǩlgTڶ�ː@���;�`0���I����K[7o�|�y�w53+���m�Fe
7O�d�$3lU�.�Ռot4�_˫r����$ш�Yb1��4W�Ȕ���ɬ�i�u}TsV��]R�����<�b�0��;v�eJ��(qq�t'�ʒ�k�')=���y?�u*�픡��&ޛD\%t9Ve�U��쨌M�7##����=\��[Uj�_��d`�e|v�ڭgᓀ~dLDFE�q��Nz%�*ڼ-��b��/�$t���g���3�I�!���*s�I[]%�Ƃ��͝��Y��4C��I�oU�	��!+�Ig$�6:�t����W+N=j��IЊ�=�Z��k\�V2TU-Zer�t��*S)&	�nݢ�}�H&j��=���_�HaS��L�*�Y��?x�S�W�8��A�@L:TD������YCg&~U���JJ2��M�����۷O�U�w��`���4�eɼ޲�CU/BӴi]��(�8��;��[��.�?G��X�(U:�N�H���Q��H�������܇�}޷G��YO�����Ǐ�믿T�o��ѽ��z�����d�1�F��(8I	�^4o�L��]KJ����MWz]=��i�suj);�7�����/�yJ�99e�2�:Oα2w�T�JG��&�;F5J�$�v42 R"=��M��R�&��x#�k2��q6e�&5��؏�d����j�k�#�\m�5�m�Q�ƈ�]���:�i{�w��`&��[�M�*>
U��1���Idsr+7,�nS�+�����]M��W���e<���X�����z�Uѩ��jH	���n����dLm�zu�o���.;�Ɂ������O���V��G��*@Ib���C���l5s��J.�J�*��<�f"W]HG���e��@u�*��d�;Y����r{��jh@o�X퓒�F�3^�kv$Y6P��7o�3e5o��u�`>?��>�P`��+\��U���Q�*��SNUC�1G9��qk%�Nӽ�0���pk���a��򎥚�gϞ�V�;���˗/׳N�`��ʒ�F^}�5|��7�бz��޽{��%�KOfo3_IU��`)�hf��0HR��g=9�!c��5>�'
��L���C�v�\�3G�f3u���@T1�Yn���5��^*�K`?�a=fu��eض-�:f��#%g�/%EO��c�6����l��ZĐ�3z��K/����)�N�p"	��(�H�`)�W5�s����OT͝Oǎs��
M�?��$&�?f��:U0��8ӟznC�u:N�n[`��(�mHNކ�9�]�]��7�B<�*=Ʒmݬ���ڷo�zi����A�p~PzȘ*�gdT}�_��Z+�و���Ы��`^+�{'O�0J�\h�8��TT�Mu�H�ʽRU}'�zY����?���_�e��]	؇���%����t򓕮�ԫ[O�Ѷ��(��Ν;u�۪v�59���v��1̍f63�٤������Y����mT�:1������]޵Ls������U���v���_�d�R8�rF[�nÌ߫�J�̭>RS�v*���� Q�������*K:ffe!.6�J����]�N�L*Svq9������m�2��Uږ����۷��~�]���R����ft���;�-^��k���Æ�;vbʔ/зO�c6C��gb����|�z���#q֠Az-i�O�^�zhּ6m�^�e�Mz�}\_s-������6��u2;�$x�����BNN�I�d�����K.�Z�%yd^�#��n�Ն^3'��%k�r�U)}���^��u��]vN9i�Q�b��yr2>��s���d6�����mZ���O�܇gq����1��_,�"��u�֣e��
[�n�ƍ��mXY�֭u��(ڨ�^�nv�*��|#d	S�z������H���.���R� 'AIa�������������t�m6\~�e��/�q�:��ٰ=y^z�%t萄���G�)�L@1y��X��?�7��s���0{;�������`�1�Х��Qe
N+LtE�i�쟱{��>���٫�^~��ߊ �y���T@�a񬁕+WaŊ�8픓z\��������s�~��*cQ6@�&MФqc�h���:�����N~3u�	[yU�5��]�}�Νqɥ�`��qz&'+�&M������ȣ�e�i�l���{((��L&�hּ��'A��9���[q۱}�f�*���]wމvm����ٻ3�NG>���ckšO�����}'R �=$�����s����>uON�2����.\�_���Ԕ�أ�d/:��]�>�p�'�se6s����巽BL��:/l�
�W]}��6�[��e����+HHH��s"�ë얔m�*�?�̳ػ�[�z"��.��{�*w�R��ۯ�;��f����0u�T64`S�����|K/���ŤI��úw>ё����3�w��S8�����^ݗ�^���k ��r�ÙY���U0���;��2�UI=�S]�h�����z�I�YN�l2����~�m�a�S��p���؟��}N_��o����W�|�^�/��,^���dNt��7�|�.e�:ݎ^��?�|UZ����&m�'N���N9�J�/9�e+V���^Cf�� ({+JO�s�=͛5�B
$��ڧo�4�GX�1�=9/�8mޜ����W|e�Q���o�nW;g�uV��i��ЭÏ4�y�d����Ə:sJ"\݀7� ��*O��+/��6]���O�^<p?ڵi��	D ����3Ĩ��x��`����E�.]�>�Yg���y�υU_��[6���c�L%rmZ�:���j߇^��*�[�V�hѪ.��|]�
���O��UW_�y��!+Ӻs܌�CR�x��'sd�Lxz��^�cǎՙ~o��N���5ADd�^��j1���<�Kܒ%�ωe@p�v�����ª���n�{�X6d��a�oa��ŸM��SZ������6�I]6mقw�yWW��L���NJ�W_}���
�۞eY
��oT���*�;�����J4�0t�0�ya:�kW�DN��c�.<��p|�ŗ��l�$,,�^{-�w��`NU��s��_���V�z~~�|��G������n|���ҫ�ɧ��?{�j�v��|��hP�~���ccbi�?��}���3rM����t�SB7ٖQ��XRU7��0l�CؽSz�Z}A}����O=���'�����y��'�u�V��c^r9��,lܸ�~����5V�Ҭ����X�W<s }����}���~��3>��S��e%��_���}��GqҀ�^�&��Zi..Z�J*���7��/�p��	'���E�������{J��}��WGw��.:s�����q�
�����"G%_��Q����g��Y::{�ٺ�����w����<k�̾t�����z�T��n_���N�e�U�Zn	ݕ蒇L6q�嗫l�	��jއ��Ds~�	���;Z�j�~���G�����84i�1��:�K)\������{�`ٲ�X�d�.�oS9��Y�|��LO��1ϣm����}݄x�Y�իWc��%�J䤏��ٳ�f�\}�5�����!)Ig ��N:mڼ	ӿ��>�[6m.�WYN�l��?��^�`NUi����{���#��]z���eMM����q���~-[�@���}f��`��ǧ�->��l\���8ѵ{<��Cz\zM����j�ɢ֭�z���];q�}`��i�ԩ���9����ߥ�q�1��+�ak�r���6`�ZD����_�uz���F`�~�+odC��v�����٧vĨĠN|��)�H@�ǲT@Vw�����}�߳|�I'�ŗơO�^���ӫWO�5��s�^��[-Į�;0�����T/5+��e<�L#����g��)Y�p!�'o��᫆����`��0���@T��b-*(�y�ر};�y�/C@��z���xRe�'O���w��4j�	ut'���=m�r����زe�*I�.��{�F���SO���WMIg�}Ʃz+U��s�^�ru2���4���as��2q�i������G��T@/�#�蚢*\����$��z��c\r�˗-��Jg�[��d!�Çӽl��J���0���{�y1�Yt��9 7�9C�F���裏b��M�ԥ��k�v��~�=�UxD�c����<��Ư��M�5�SÇ��T����hеR*0H&2?� ���C�v�m�#遽i�z���˯��uהφ������3#��y�&x��q�X���d������u2
���X|�\������{�a���HP����z�Q^���ß�Rsx��e�^�6mZc��Q�q��ɖ��\+o�:W�L�ÿ��[q��w�I�FKdH��a�����ß��E���^)z����I���ʕ[�ҵ�J܆�63���&%ntlɽ�X}wF??J��ߞ�6�I/k�Mi�W��*�+�[^F���mݦ-�����
�\�����G��X����f
�))ػo��Ŧj�
��k����={b�ĉ��������H�|=�ze��W��SO;��s7�W���$��;g�^Fv�8���-2����U�9�s��:�	���K����ݺu�Čp�3���^��:�=��Ӻ���W^����aZ� X�E�ʻ���=22��q�}�����DU�]N_�#�=���{?v�H��A����HNN>f+\)���ˣ�����?��ުґCf�[�j5������G���!O�[OO[y�5W��s��OH�۽kL��:��x������,l.�H�M���O���O9�]w�^�F&�����^!N����5Z��W�������@�S�Z4���q��^��z�Ksp�	�>����*�e���G~y]lt4n��z=c�dοV���7��~?3��C���
�Q1�ر��Tw���6jРR���Ɏ�{��^�Z���bu<��qD��Is�|��F��}\(oi���9nӦ��=Opv�A�Н�����Ti����õ�K�L���m.���lݲUw�������HH�G�vmq�	'b��A�ӻ7��M�[�*Ty_҃]ޓ�������3�`�?ر}������К�fG�
�mU�\f�2dN:i �={+}��^�[�e�v:�zᜰ��Wmʾ���t�ֽ�LWr��I�V�!5r���֭[�kWu���Ǒ��S�Jur��=�d�%�v��!`��ʔ��{�,�w9���� ̋.׿Es�믎Ӷm�A�Hy�:��2r�sz����9?��ʕ+�����ɽe\
Oa���Eb�D����w.NS%r����Vi�٣�
n9% ��e��/=���tb릮yZڡ��/Sjk���W�\i^�fK��|���i�Oزy3���c��B��Zj3dTP||�����K����]],�J���մNG�s��gC�t�8�3t�;v"y{�^&TƖ������Y���HH�ڵ�PO���5k�\y�W]�fw���[�9��&w���ur�v�Y�F�N�e��Y%#=]�Ws�$*�j��^f��ر:w�W��#d����׫�	Z2���$�뮻���V"""W��+�I���>����QQQ~�ŕ��qϊ]�#>@���S�/�r�p��}e�#������-7�d��|b��+}lԵ�N����6m�ڵk�z��}�����lnn���bս.�=˒��ڵC'��v�{�Z�Z�
��s;��S��w�-kO�\�����S�|��/-�%� _��C�:�����Sqݮ

�����~%'�:u�ѨQC4i�T��1�2�S�
Ԭr�"�W݌�*ˣg����ِ\���5���@$��A)J%J2�Qj�����_��%�o��>�]� C��2w�zߒ ��� ��Ë����}�u�Dӓp�:�ʪ���qU{�o�VD�=��������"�LU}��qq�Q��)�/�I���&=ⳳ���ס�}��$�(:yHf˰�O�H/����r�;P�7��aUu<O�Tc��Q�9��k������΀^)f�K)C�\����b?�w,��#��L�im/��;�hݥ��8��|��8ގ)�ňp�z�����<��58��0K���0�~L��6�@;�\{u�yy�PM����Ni��f7����YB'""
f�S\�[y:�Q�ѝ8�)������^����3�-ӯ6�|v�#""
b���������(�ٝN��ֈ���7=S\�[�,HN�Љ������W~	]�9:����T:v���3M�r'"":�����,�Tn�7+�O"""
�K�ݯ8-%tFt""��d��m�::QPR1����DDDAKW��UBg�8""��e��˝Et""��U�:#:QP���U��8t""�`&U�~lU�?"""
F��ΈNDD�̊��3�)݆ι܉���;��~e/w""�����,�NDD�L��YB'""
jXm�m�DDD��"���������r�z�DDD՞S�r�5""����U*�}�k�r'""
ZR���VN�f,'""
fz�5?7eX'""
V�ߋ�0�'��,�U{�˧2�5?�r�܉�����m�r'""
b��U��DDDA��Nq�����(��~W�Q�b�;Q�Ǚ∈�B g�#""
~�C�˧2�+��^��DDDA���2DDD�ʏ�\�L��NDD���ΨNDD�����*w""���*w""�`�ʝ��(p�8""����kb=S+'�܉��B ;�U\m������K�p.w""�����\�DDD���X�U�DDDA��Q��LqDDD!����,DDD�*�˝m�DDDA�ɉe�������CgX'""
R�
T�Q�͉e���B��m�&�܉������6t"""
F�U��Gk��DDD����܉����
t�#""�`���WЉ����Dh�m��(񃈈���aT$��UBw8�HKK�!�p���� �`PS
Q���c�=�l����j���둓��ז�n��0l�C��Wæ�5�������]8
�������p����*�&6���e��-�8\yS~U��^�t1����h2�g�.��6��sDDDt�I��f4��&��� ""��JJ�:�烈���+UB7��͖n:�� ""��Hfsأ��ege�U;6�-3:::�^�n��������{�g��0=""�I&������K���;w$�Өqӻ<�t^^^/�4cTD��u�ƪ�3*8���c:1ϑ��g�#|���g��OF��x���$�����jժ�y�����W�<l��k�ŧ�O����;v����LP�F��]mn�G���E��l6�&m�v��0�æ�`ap�4�����rd��ϫXf��Ta���
�+����ſ�F�_JoWl����l�	�Q�k1׉x����󇢿B�8*�g�J����b{/���}����(:f��Qxn(���.u��{�`[�~���0T�.b�ҥ�{v�
/���G���NC�&M�T�^n7TWr�֬Y����[f�������=��ILl�o�Nɟ�f��MX�<[Q��}y�~����1�\4%�Y�wϮ�����,�{������vW��3K���yxv�c?%�l�Kb�R��\��W���)|q9��,q%��[����ĮK��}���n�a���{��_�]�r)�'�z_/)���N�l�b+��(�-6-�Y�b����J�-��ڨ�9��G�}{ΧԖ����t��pJ�e���%���-:�b�G�J�JM����.rџ�ݠ��:IϹ��\�������0̘�hg|BvIIs�����Saw���ʇ���G4�΅�Ϡ ?W?j"�gY"P������Ӑ@�p��ÐB�l�S�t8W pr�����T$u:�Õ��p?����w���&���\]$�b��$�o�^ܙ���kѾ����m6�����u�]o�ٽ�ً\t�Ÿ��[Bnn�;z��͸�λt"Q���N���on���'�<�������OOL�<O�EyUw�g��&�%�f�L������õ�Y�I�?\���u����hY<u���	S�,�;u):/��s�]6
ӛb�r�����
_��G���R�����̰�^����kc��4�ͦs�6Wy��-5�0�\�����6�]^cs[�e�._�CA��o��0RB�zHٿo��>�S?�� O�l٪UH��7�

���Vtx�is8t��4��J4�m�j��m�w��/�(5�_�O!_ega2�J%J��#��X�]<�g�إ{�i�'6�^�٧�Lexb�Y��Z�;�'���|��������Jl��2y�.�-�܌Ȉ��Zu#WD ��x���\���j�ژ��~̯s~Y߿}���E���[_a��p�2�mW|�ҥ�R��(�P�F�s+��(��/��(]�*��2�M��x�k�9��?ós�t�<�t�B�{��#�?=�Og^�{Tx6�k��F��'�����ܙ��r����w��=��M\�C���x�y0e[��|�}������vU��2��pU"R��Ɂ�
��c8�Զ��r���گ�S������r�Jt�ܹ�ug����e�,���o��� ����W;����"�#

�eF���e���سgZ6o�/S�T婌���o�c��-]:�mҬ�ks�u���'`��u���+AD,Щ���T<�$$$����J��ʬWr[�l���kt@�`.�;���*CS���f�^��?�>��t��6��{�Q0a@�2ڷh�ǞxR�����v��V&����a�?�`��A�>������_<��sػG��R���Jn߱ø���vh�] "
F�d�q�&�ݧw�_|�^�ڵ����������:��m;����x�駱j�
������f͚���/s�~y��6�w�� "
6�d)-��p|n���V���]*�J[�j5�nۊݺ�:ҝ���1f��y�l�i80ԫW��O>��/��Lꐄ�cǂ�(1���N�#:&f�
�y*�G��¦;�-Y��������λ����(�	N����h׾ݘO?�$%'�0���:Y�6�6m�ʔ���#���5*�M^n6����\s"��Q����{���K���@��0�=�Q��o��}�'�?�fM��;�"�`ŀN�.��b\{��6�#""|Wf��Ȫ/���K����^�jӎ.�bي�1b$��މ��\�����g��w�;��>�Y'>�G<"�`ƀN^����۴9�����U��Uv[�n����t@�$������ѣ�d�b�	�JtTTr��-�L�655/;DD�:y����`r�ڴi�Ff�*;ͫ��b�e8���Q���㭉1��o`5���W��k�.���� �n��O?"�`ǀN^}�~.����j���s�yyQ��q8�p�"���"*22��g��oLx��ٰ*�׊��ѭG��Np�����޻o���:`@'��M�ݺ�@TT�&e~^nS�v�U+Wb_J
Z4k�`�i75r����`��y���ϛ�����C��޻Љ��`@'��z�\vŕ��Ď�QQ۳27-���m۶bÆ�A�u��~w��b�vs�ݞݰA��+W,[8��G�Գ;n��jU��S߾}p�ק�<{�Z〭�%�:tK�.����`$����˒�����|�)�ߓ���mxi� "�N�ɧ����
���e�Ͷ��뻗�t`ѢE��ɑ�AՎ.'+��'�h7���]ٮ}����-c��� "���ɧ_�͚�D�:�W���g��^�j;iG߻oZ�h�`�״����p���n7���hܴ�����)_}��K�aԨ "�n�ɧ��.B�=l˚ի����Xt��۱~���	��SRS1z��^Ǜ6�,����\�պ�k0�|���K "��Щ\	uиq�ݪ�%=-�M�-����y��y�5�fϓv�I����v��:uz��/�ʱ���)�����b@�ru��I��9�U�a�Q�c�t`������Flt�1oG�v�7&L���[��#���7o�r�/?��y���ؽsN?�tUW�T.w�8�{�^�򚣠� �j�U+Wa�޽hӪ��x�#Gc��vsy6���s�͜�����O��3O���:c@�r͚5]��@|B����������e���ؾ�֭?f��<�`�E���_{�����/���w'OQuǀN�:��q�7�t:��/]�+++�n٭����v��:��(���y�EtL̎�mڌ�����0 ��Qv;"����_�z����/��?x�`�mLӡ�S���BlL�QoG�����7����`n���7i������3#����`ND!���Ҹi�rӍ��:���l��]y�e���ػwڴnu��MB�Ju\�j߻w,�����P��'�<��AC�1۶m��oL Q�`@'�<��Ø��iG_�J�9y+�Ihݹs'�o�p��������`���n��]�v�g�������q��_3�QHa@'�HǸ�I���Y����J,�v�e˖��AgU�9I0�/(��＋iS�I�?����#�7i����[2���ѳ[Q#��ÀN~��q=��t"۵�߅�2�3,�V3��ѳ��sƣ�4�g���k��΄U����s/�`J��]�v�Z<x߽ "
5���m����n94��S��`5��X�z��KA�U3�g��u6�y�w��˪vUX��]��Ν;��釙Y���� "
E����Cҹ�ٳW��av�� ?�2��x�M7VY@��JO�ر�������n�ڢeˑsf��)�a��_����Q(b@'�=8t(>��+ԩS{UDDxFA~^�	f��Ұt�2�y��*9��~�?|���0M'���e6���Mz��W�r�x���0⹧AD���o���Z�i���M��ѻ�23�Xm�׽*�G����ܹxy����̀uU���s���Mxz�3�5�[��ND!���ֿ�?^Ƥ����/������m�5�Wc_J
Z6o��K0߲u+F��m[7���m�ڷ����{�r���_���?Q(c@�
9����1))�s�n+m6���Hޖ�M�6,�K0����K/��彩�-�����4m�t��?��9���дi\q� "
u�T!��ɨ];			K#""rsrr"�n�jG_�l�vj@��0M|��g���>���U��a��~�ĩ���K/3���1�Y��Q���N2��3q�"22r}dT�����&V������%K�������J������k>^�"2��[���ۻ��*�<��?�����n4$kBGMk׭�bv�r�s'k7��f�v�Y�j^Rlk�Uh3#l[��dE!0�&"��*'8��e7��s�[�<|?3g8����w��9���L����ܶ�3� ���~�>*J���k������%��8m�F�Y�Dz򃴘מ���5k��\���G�|}[Ǎ�� ���T�|~�3y��' ���~�6�f��ҥm�3�t��_`�Kjj���ٳ
����Z:;e}F��������zWxDĎ�~����
� ?_�n� �pB��oK�zJ[`ƞp�m%��e����A�%-�-RRR"���;�jQ��y_v��]v�����	:���cGW@@���1��v:��Ç%.>ABCCK||}�m6k�����V)*:!]6�x�}:��W���Xa��MY+��f�����	�����Z�N��M*{��:�m������gŠ7T;v��J{{���_�|%M�&�w����74HRR��*+�^Q���ᆌ=|��W^����አc@�B�d��Sr?ʭ���0�Ӹ��*����	z_h1���ƍ�$���<��
�?w�?����/�k� W29�$��ϲ.%��*�~���p3J�su^ZZ*�Ϝ��s�ݷW�l�"6�U<͛�Un���o�ަ��RXX(��� �pE�1 ?��DG��M�'����X-���q6[�?^$֧�b4��禥�Dq�$'�H���t�����=>�Ճ���; �.\���x�ጠc@���f�~��������k�X:�=]Mk����-�q];��,)�k�d�	����N'QQQ{�WO�?c��v����+ �;��������L1u�
�k/{�$?w��������&[�n�?�#�}��Z!�!E3�e���hjn�m��  A� ����c�>bޙ�uZ���{ڨ���(��e2c�t���ҝ��'37HW�7ڢ�r�K�Z~:yrʮ���t�3R[^..  A� DDE�,0��_�Sl��~�����(/���EEb�Q����{W���%yM����Iϭv7��Fo׍��;�צ~x�;��Ȋ�� �_6w�,���Hxxx�ȑ#-�W�~�o�����XZ��亠����F6��Jj�:���/�Ӽ���ZdT�;�ߙ�>����%9�� �w:L�"uz\����-��dn�����R[S��o����)ٻ����i��%A����3��^{�g5���*� �C�1`�G����>Ѿ^��Ω����t��_� {��S�Iz}O���]��.�X����s����s�bc7�d��ߕ�P�1���y� ��:eF|��
h	)3��6���8m]��۷K��Y2g�,�8wN��$u_�WK/��i���_�Т7W�|�.�,~H  �"���ks��y��t����ߔNj��%=-]���$c}�=rD<=��]�GFF��=gv�ƍ�N����
 �cP^߲E��#gΜ)�;엺�����򤪲J*����Ԗ�u?o8j��֙�fnX���g�!�>yR  �t��%�n�Nʻ�|\z��t~�)�'��MR�e���i�L�]���훶lq���ɯ�<)  �:�d2ɒ����������ں��tz�~���w'L�X}Ͻ��ݺu���ݻD�d;A��tZ��J�:m��/>q����ā��%�GZܽ s�����j��u�̝@t�'��˧G���;�x�iʦ���X�V����`0J\|\ުU�v,8䊈���� �aC��?��{\Ǝ���?���b}�.�K��`4��W�Ǜ��j����pF�1$��^��:f츎�G������q���>��K:�n[xT��i�ؤ���[� �Cf�Ν��ޮm�r�������T����C�i�+��<�����-�  ����2˖,��/���s�J�ط���w���-���*<!!��]wߕ|������� }G�1���ِ������l�X��m�I=��������3>m�^9��ŕ���*/���  ���cH͙3Gv��-oeeɁ��"_�$�ݑ�]�Qn���z�;f�y��g�9��ӈ9 Aǐ[�x��d2���D����t:&8�UN���|�����`4�1��Eǋ���ʤ��V  C��8UZ*:�QBCB�'LL375�X::��lA:�����'wtp��u��wZ,�z�j1M�$ ��!���86ih��^��������dn�:V: `�:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
�O��Ր���    IEND�B`�PK
     8p�[��EM  M  /   images/d3694a2e-5bba-40c3-8069-8db85c4c9209.png�PNG

   IHDR   d   d   p�T  TiCCPICC Profile  x�c``RI,(�aa``��+)
rwR���R`����b
����>@%0|����/��:%5�I�^��b��Ջ�D������d ��S��JS�l����):
Ȟb�C�@�$�XMH�3�}�VH�H�����IBOGbC�n��ₜ�J� c���Ԋ�_PY���Q���Tϼd=#CsP�CT�%���X�}�����ߍ�������k'BLÂ�A�����΂ĢD�33��10|Z����� |�'�8��,������z����j��N��������.j���p  !e�2���   	pHYs  %  %IR$�   xeXIfII*            (           J       R   i�    Z       %     %      �    o  �           a���  �zTXtRaw profile type icc  x��S[n�0��)z^�8~$R��b;^eW�J�ё"�@`H�n-|DI�D��@ȴ�v=L�"�	�s,`�ۮ��z����"H����pz����3�ͬ,9&�h'�tN9#���(���d>CQ�h�|q�k��R�R����mOi�q�6�Z�ܶ=���C�>hrK$>���U`�͚t3�s;����%�S�T�c��\���~�y§b�_"%�G"a=}J�H����|)�Ni����2��yl�c���r�E��|�7$��8��s���.PJ����
��wq�8��P'��j����[ܞ�c2����g�+��|����RM�=�c2gҥl��ϞauTh���҈�\�z���줡㜥   %tEXtdate:create 2020-01-31T21:31:09+00:00��y{   %tEXtdate:modify 2020-01-31T21:31:00+00:00	�   tEXtexif:ExifOffset 90Y�ޛ   tEXtexif:PixelXDimension 1391c�   tEXtexif:PixelYDimension 800�요   (tEXticc:copyright Copyright Apple Inc., 2017���   tEXticc:description Display P3�y��  cIDATx��]	xLW~��d�(%�J"��}�%(�Z���B��_[y~R�R[u�E[[����J����ҿZ��j��B)��'s��;��Ĉ����>���=��s�s��-�37:�PTB��A%DaP	QTB��A%DaP	QTB��A%DaP	QTB��A%DaP	QTB��AW÷&��z\I���7�)I*�Ev�Z�:d;iJ�3mtRɲ�������V�$IY6��"a[�d��$}/����~�l���99��t.��$u0Z��d�M��(��5D��a�}0�*�
��?���h��dY~�`ȫq+��L��yY���@���[���������ƍ����0��`�Aк�C��"�|<B&�������r����t�PQ:�;w'N�{˧����a)y���3�t>���ʂ
E@fB\yyP� �f�3b�1�(p�3!�<ÃY=��䫄(�d���?0��&1A3vH�JIi�	�YCd��c,�p?��0���g�Ж���lqtws���%b�G��ɒ�2d'jaxR�v�Zl߈s��S�����_C���2Js;�i���8�f�ɒM>�Q.]�����С�x�g/�5J<����зO̚=�g����f6.:6lX�t]������B��5�D��;ѽ[7���s�p�0g�,�n�=_x��(���E��~/���u{���F�m�6�2�h��!����v����;����dX�i5�7�}�����ٿ�2~޳?��#n������1p�@xV�$��u˖�Ѳe��H�zi��|��u��,�Ν'�����ԩ3�/�5PP��7o���,�_���C�޽ѵK���ǚ5k�t�:>�,^|q 4�XȺ����7!&&�+{�_�~��d��ǎ	SԥkW�o؀������A��n��B�p2�7n����Na��>$3��ARLN�G��&����~�� �����QQ��wq�������Тe+xU�ºu_ lQ������͐�լ�K�.����ԙK�.��9����(�QN4|���X�p&M|�����5�OLLDu��x�"�.Y�9o��&�l7ww7�b�rD�c�)��?��޽E��jO����[���a�0�?B��ۿr6n����o�Y�}��E�E�:uh@lAZZ*�i`5]�ر�u�9Ǻ��<s�4�V���ի۽��1�Q�n�:AƢ����D�?O�F�g:b����a� i4puuÑ�#������W��u� ̜�iL8^<H�Ȏ��ʕ+Bui������®�v�u�zS����u>l�ФΝ�P�U�@.��+��������^M�5c�L�L��S��nW",�Y��e��'""#�|���'B�B�FMТœ8���	�R��ӓC��w��t�b�_G�R׿ƛG߭~=L�6U��?���קў��ݻ[��Z���\�rLd0�q�	��o@Ey.D<kI��
2^U��~�zB�!C^65V�E�6m�W���$!-^�j� ��溃��������͂�٤������m׮j׮����{��l"��e����G�fg�AQ�%{ΫbM�6��F�흚6m"�.\@�ƍD���]P��	��g�ΕG���e?h�V��\��ӊ�����ٳq"m���`1i.�[8c:fd��Y����<P��6���׻�2�sq�{dDG2kd'j	h�͛��)2;U�jW��%�=z|j���)�b~b����!JcӁ�L��+$3�i��ߪ[�Fc�8����2�F����~~���dG��?��%\�9���ɡ���3lw[wGDD���Ç�6�V�Z8AQ?��6U_"���YԢq�0��$��_M�i������W[P��@�nns+�F*Z��@'����!����ǤI��`�<a�CI�>��p������<*T�[�Cɩ�1K�,>�>}�/�h�M�vhD�*��89�-�aq�֭�M0m�t�jQt������5k?C��M�ۻ�Mk5���Z�e����ZSVY'�����L���������'����F����g(4�Ŷ��P�^G�>|<(��p������_�R�VUDK</`9rr��WhI�6��E^��9��~��΁�ʧ(��K�c��K�^���}Ѭis<���b�s���J�efp �e
���,���5��<�5o۶oD��h���%.�sab��F��%a�ȑ4I܍��u�Ȗ-�!00�==̤?�9@���������A��"���K�T����J��2
�������r�̋h���C�Шn+���\�t	�i~`�'t�dA�����Ӄ|�'���GEDCQ��z�5{zP�gA`�@��?�h����\�h*��5���]�r^^^pbb(��1��[ޒbo�ػ^8�s4�叽|�4�@����4}�#0(h�my
?A�#����Mg�<��7��?�il���_ �2Eto�����"����j�37-N^��4g��)�8����&��'�*JBCLQ�JH�C���=d��,���}X5D�2`�����0��g窆(&Q#,���!�.o���e�TF��[���9ʲIQ�[�<l�M�V��|/="D�xOR���vG�_G�3˚��7��aj�gE��s�6��ˋk�Q'I����܊�GBEiB���j���QCG�h4Z�D�$ݢY�-R��By%�V+i�T���I|3����4����ĉؙ}���2r����)���Om�fk\]�zH�|�R�iO�l�Mۗ�I6_dْϜf4G��Fk-匷�ݥe�k�\𛍶���V���_�3���X:�-�b(ڴ#ݾ���KĤ����h$�v!VI~}��+s�^����xg��p�h4"�E@�Ӈ$^N������1���	�����ǁ=j��������o��qbZW�?��i�1��wI�t�G��v��e��^3�x޹���k+�t�w��`-;q<3��rJ�r�##���Κr$55G��޶;�a�±c_�ٿΜ�V�{J9�Ԕd��=�(B���}�\�.1�7����׭w�^v�.\�[��"{x<����̣������{�"o���]�|ҵ�"#��[v��n�ٻoޚ>�Mۢ�̛;[�A���(Ks�#�����@�V�s��I������׸��������gn�fV��8\��@�*e	%F��#�n�����8v� �2�Ǎƙ3�2+yV{<6���ܜ����#d9�¡��ȏ ""�z�ז-_�M���^nzjJ�QNk��i�܇��#��~_�Z(_��?���&��2�G9��ɡ�=�gge|�yx�fY$�Q�/R~�'������ll���<����� ~�N�z�����t
s�PVQ��<^�q�s��mOrrJ@�=�t-���K		粲24x6�;�;�%JHJJ
*�|D��-KKMN!p5�olI�x��ݺ�Ge�F��kǏ�H�"A�ռ!i\�xzz�/_�<�R�u�7�u�����U�F��K0��N�rx����̬L�(B���^b���x:y9��}���E������k��%u����QTB��A%DaP	QTB��A%DaP	QTB��A%DaP	QTB��A%DaP	QTB����Blg���    IEND�B`�PK 
     8p�[_6c�  c�                   cirkitFile.jsonPK 
     8p�[                        ��  jsons/PK 
     8p�[��LQ  Q               ��  jsons/user_defined.jsonPK 
     8p�[                        :�  images/PK 
     8p�[����^� ^� /             _�  images/8a866263-8c14-4821-a3ed-cf7b88c4ff1b.pngPK 
     8p�[����  �  /             
v images/b53b2c7c-bb6b-4047-8ddd-b279832d777a.pngPK 
     8p�[�ة� � /             '� images/8f771a2d-db90-4bfd-8b3e-8d66edcda07a.pngPK 
     8p�[��/F��  ��  /             � images/0c7fd013-2f4e-47d0-a46e-2d19cc1fd6f6.pngPK 
     8p�[�c��f  �f  /             � images/c88b2895-5e8b-4a57-9f9a-b80dd50058b1.pngPK 
     8p�[��EM  M  /             !	 images/d3694a2e-5bba-40c3-8069-8db85c4c9209.pngPK    
 
   �	   