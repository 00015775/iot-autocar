PK
     �k�[�O�k�  k�     cirkitFile.json{"raven_core_version":15,"hardware_version":0,"pin_to_graph":{"pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_0":[],"pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_1":[],"pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_2":[],"pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_3":[],"pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_4":[],"pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_5":[],"pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_6":[],"pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_7":[],"pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_8":[],"pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_10":["pin-type-component_68cda57c-349d-45e9-a6a2-98cf0cbc2416_4"],"pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_11":[],"pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_12":[],"pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_13":[],"pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_14":[],"pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_16":["pin-type-component_68cda57c-349d-45e9-a6a2-98cf0cbc2416_0"],"pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_18":[],"pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_19":[],"pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_20":[],"pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_21":[],"pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_22":[],"pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_23":[],"pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_24":["pin-type-component_68cda57c-349d-45e9-a6a2-98cf0cbc2416_11"],"pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_25":[],"pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_27":["pin-type-component_68cda57c-349d-45e9-a6a2-98cf0cbc2416_1"],"pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_28":["pin-type-component_68cda57c-349d-45e9-a6a2-98cf0cbc2416_5"],"pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_29":[],"pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_30":[],"pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_31":[],"pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_32":[],"pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_33":[],"pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_34":[],"pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_35":[],"pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_36":[],"pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_37":["pin-type-breadboard_ded8e15a-344e-4f93-a7cd-807af81d5cc8_0_0"],"pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_38":[],"pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_39":[],"pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_40":["pin-type-component_68cda57c-349d-45e9-a6a2-98cf0cbc2416_3"],"pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_41":[],"pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_15":[],"pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_17":[],"pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_9":[],"pin-type-component_68cda57c-349d-45e9-a6a2-98cf0cbc2416_0":["pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_16"],"pin-type-component_68cda57c-349d-45e9-a6a2-98cf0cbc2416_1":["pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_27"],"pin-type-component_68cda57c-349d-45e9-a6a2-98cf0cbc2416_2":[],"pin-type-component_68cda57c-349d-45e9-a6a2-98cf0cbc2416_3":["pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_40"],"pin-type-component_68cda57c-349d-45e9-a6a2-98cf0cbc2416_4":["pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_10"],"pin-type-component_68cda57c-349d-45e9-a6a2-98cf0cbc2416_5":["pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_28"],"pin-type-component_68cda57c-349d-45e9-a6a2-98cf0cbc2416_6":["pin-type-component_c3c8c3f0-5cb8-46df-9e8e-6bc9ea246e79_1"],"pin-type-component_68cda57c-349d-45e9-a6a2-98cf0cbc2416_7":["pin-type-component_c3c8c3f0-5cb8-46df-9e8e-6bc9ea246e79_0"],"pin-type-component_68cda57c-349d-45e9-a6a2-98cf0cbc2416_8":["pin-type-component_fc7a62c0-bbca-4c4c-a089-8837f2378795_0"],"pin-type-component_68cda57c-349d-45e9-a6a2-98cf0cbc2416_9":["pin-type-component_fc7a62c0-bbca-4c4c-a089-8837f2378795_1"],"pin-type-component_68cda57c-349d-45e9-a6a2-98cf0cbc2416_10":[],"pin-type-component_68cda57c-349d-45e9-a6a2-98cf0cbc2416_11":["pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_24"],"pin-type-component_68cda57c-349d-45e9-a6a2-98cf0cbc2416_12":[],"pin-type-component_68cda57c-349d-45e9-a6a2-98cf0cbc2416_13":[],"pin-type-component_68cda57c-349d-45e9-a6a2-98cf0cbc2416_14":["pin-type-component_db7d8f7f-8f6f-44a8-be93-8d8d7b68807d_1"],"pin-type-component_68cda57c-349d-45e9-a6a2-98cf0cbc2416_15":["pin-type-component_db7d8f7f-8f6f-44a8-be93-8d8d7b68807d_0","pin-type-breadboard_ded8e15a-344e-4f93-a7cd-807af81d5cc8_0_0"],"pin-type-component_68cda57c-349d-45e9-a6a2-98cf0cbc2416_16":[],"pin-type-component_fc7a62c0-bbca-4c4c-a089-8837f2378795_0":["pin-type-component_68cda57c-349d-45e9-a6a2-98cf0cbc2416_8"],"pin-type-component_fc7a62c0-bbca-4c4c-a089-8837f2378795_1":["pin-type-component_68cda57c-349d-45e9-a6a2-98cf0cbc2416_9"],"pin-type-component_c3c8c3f0-5cb8-46df-9e8e-6bc9ea246e79_0":["pin-type-component_68cda57c-349d-45e9-a6a2-98cf0cbc2416_7"],"pin-type-component_c3c8c3f0-5cb8-46df-9e8e-6bc9ea246e79_1":["pin-type-component_68cda57c-349d-45e9-a6a2-98cf0cbc2416_6"],"pin-type-component_db7d8f7f-8f6f-44a8-be93-8d8d7b68807d_0":["pin-type-component_68cda57c-349d-45e9-a6a2-98cf0cbc2416_15"],"pin-type-component_db7d8f7f-8f6f-44a8-be93-8d8d7b68807d_1":["pin-type-component_68cda57c-349d-45e9-a6a2-98cf0cbc2416_14"],"pin-type-breadboard_ded8e15a-344e-4f93-a7cd-807af81d5cc8_0_0":["pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_37","pin-type-component_68cda57c-349d-45e9-a6a2-98cf0cbc2416_15"],"pin-type-breadboard_ded8e15a-344e-4f93-a7cd-807af81d5cc8_1_0":[],"pin-type-breadboard_ded8e15a-344e-4f93-a7cd-807af81d5cc8_0_1":[],"pin-type-breadboard_ded8e15a-344e-4f93-a7cd-807af81d5cc8_1_1":[],"pin-type-breadboard_ded8e15a-344e-4f93-a7cd-807af81d5cc8_0_2":[],"pin-type-breadboard_ded8e15a-344e-4f93-a7cd-807af81d5cc8_1_2":[],"pin-type-breadboard_ded8e15a-344e-4f93-a7cd-807af81d5cc8_0_3":[],"pin-type-breadboard_ded8e15a-344e-4f93-a7cd-807af81d5cc8_1_3":[],"pin-type-breadboard_ded8e15a-344e-4f93-a7cd-807af81d5cc8_0_4":[],"pin-type-breadboard_ded8e15a-344e-4f93-a7cd-807af81d5cc8_1_4":[],"pin-type-breadboard_ded8e15a-344e-4f93-a7cd-807af81d5cc8_0_5":[],"pin-type-breadboard_ded8e15a-344e-4f93-a7cd-807af81d5cc8_1_5":[],"pin-type-breadboard_ded8e15a-344e-4f93-a7cd-807af81d5cc8_0_6":[],"pin-type-breadboard_ded8e15a-344e-4f93-a7cd-807af81d5cc8_1_6":[],"pin-type-breadboard_ded8e15a-344e-4f93-a7cd-807af81d5cc8_0_7":[],"pin-type-breadboard_ded8e15a-344e-4f93-a7cd-807af81d5cc8_1_7":[],"pin-type-breadboard_ded8e15a-344e-4f93-a7cd-807af81d5cc8_0_8":[],"pin-type-breadboard_ded8e15a-344e-4f93-a7cd-807af81d5cc8_1_8":[],"pin-type-breadboard_ded8e15a-344e-4f93-a7cd-807af81d5cc8_0_9":[],"pin-type-breadboard_ded8e15a-344e-4f93-a7cd-807af81d5cc8_1_9":[],"pin-type-breadboard_ded8e15a-344e-4f93-a7cd-807af81d5cc8_0_10":[],"pin-type-breadboard_ded8e15a-344e-4f93-a7cd-807af81d5cc8_1_10":[],"pin-type-breadboard_ded8e15a-344e-4f93-a7cd-807af81d5cc8_0_11":[],"pin-type-breadboard_ded8e15a-344e-4f93-a7cd-807af81d5cc8_1_11":[],"pin-type-breadboard_ded8e15a-344e-4f93-a7cd-807af81d5cc8_0_12":[],"pin-type-breadboard_ded8e15a-344e-4f93-a7cd-807af81d5cc8_1_12":[],"pin-type-breadboard_ded8e15a-344e-4f93-a7cd-807af81d5cc8_0_13":[],"pin-type-breadboard_ded8e15a-344e-4f93-a7cd-807af81d5cc8_1_13":[],"pin-type-breadboard_ded8e15a-344e-4f93-a7cd-807af81d5cc8_0_14":[],"pin-type-breadboard_ded8e15a-344e-4f93-a7cd-807af81d5cc8_1_14":[],"pin-type-breadboard_ded8e15a-344e-4f93-a7cd-807af81d5cc8_0_15":[],"pin-type-breadboard_ded8e15a-344e-4f93-a7cd-807af81d5cc8_1_15":[],"pin-type-breadboard_ded8e15a-344e-4f93-a7cd-807af81d5cc8_0_16":[],"pin-type-breadboard_ded8e15a-344e-4f93-a7cd-807af81d5cc8_1_16":[]},"pin_to_color":{"pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_0":"#000000","pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_1":"#000000","pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_2":"#000000","pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_3":"#000000","pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_4":"#000000","pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_5":"#000000","pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_6":"#000000","pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_7":"#000000","pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_8":"#000000","pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_10":"#ff2600","pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_11":"#000000","pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_12":"#000000","pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_13":"#000000","pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_14":"#000000","pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_16":"#00f900","pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_18":"#000000","pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_19":"#000000","pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_20":"#000000","pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_21":"#000000","pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_22":"#000000","pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_23":"#000000","pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_24":"#874efe","pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_25":"#000000","pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_27":"#fffb00","pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_28":"#ff9300","pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_29":"#000000","pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_30":"#000000","pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_31":"#000000","pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_32":"#000000","pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_33":"#000000","pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_34":"#000000","pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_35":"#000000","pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_36":"#000000","pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_37":"#000000","pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_38":"#000000","pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_39":"#000000","pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_40":"#aa7942","pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_41":"#000000","pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_15":"#000000","pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_17":"#000000","pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_9":"#000000","pin-type-component_68cda57c-349d-45e9-a6a2-98cf0cbc2416_0":"#00f900","pin-type-component_68cda57c-349d-45e9-a6a2-98cf0cbc2416_1":"#fffb00","pin-type-component_68cda57c-349d-45e9-a6a2-98cf0cbc2416_2":"#000000","pin-type-component_68cda57c-349d-45e9-a6a2-98cf0cbc2416_3":"#aa7942","pin-type-component_68cda57c-349d-45e9-a6a2-98cf0cbc2416_4":"#ff2600","pin-type-component_68cda57c-349d-45e9-a6a2-98cf0cbc2416_5":"#ff9300","pin-type-component_68cda57c-349d-45e9-a6a2-98cf0cbc2416_6":"#000000","pin-type-component_68cda57c-349d-45e9-a6a2-98cf0cbc2416_7":"#ff2600","pin-type-component_68cda57c-349d-45e9-a6a2-98cf0cbc2416_8":"#ff2600","pin-type-component_68cda57c-349d-45e9-a6a2-98cf0cbc2416_9":"#000000","pin-type-component_68cda57c-349d-45e9-a6a2-98cf0cbc2416_10":"#000000","pin-type-component_68cda57c-349d-45e9-a6a2-98cf0cbc2416_11":"#874efe","pin-type-component_68cda57c-349d-45e9-a6a2-98cf0cbc2416_12":"#000000","pin-type-component_68cda57c-349d-45e9-a6a2-98cf0cbc2416_13":"#000000","pin-type-component_68cda57c-349d-45e9-a6a2-98cf0cbc2416_14":"#ff2600","pin-type-component_68cda57c-349d-45e9-a6a2-98cf0cbc2416_15":"#000000","pin-type-component_68cda57c-349d-45e9-a6a2-98cf0cbc2416_16":"#000000","pin-type-component_fc7a62c0-bbca-4c4c-a089-8837f2378795_0":"#ff2600","pin-type-component_fc7a62c0-bbca-4c4c-a089-8837f2378795_1":"#000000","pin-type-component_c3c8c3f0-5cb8-46df-9e8e-6bc9ea246e79_0":"#ff2600","pin-type-component_c3c8c3f0-5cb8-46df-9e8e-6bc9ea246e79_1":"#000000","pin-type-component_db7d8f7f-8f6f-44a8-be93-8d8d7b68807d_0":"#000000","pin-type-component_db7d8f7f-8f6f-44a8-be93-8d8d7b68807d_1":"#ff2600","pin-type-breadboard_ded8e15a-344e-4f93-a7cd-807af81d5cc8_0_0":"#000000","pin-type-breadboard_ded8e15a-344e-4f93-a7cd-807af81d5cc8_1_0":"#000000","pin-type-breadboard_ded8e15a-344e-4f93-a7cd-807af81d5cc8_0_1":"#000000","pin-type-breadboard_ded8e15a-344e-4f93-a7cd-807af81d5cc8_1_1":"#000000","pin-type-breadboard_ded8e15a-344e-4f93-a7cd-807af81d5cc8_0_2":"#000000","pin-type-breadboard_ded8e15a-344e-4f93-a7cd-807af81d5cc8_1_2":"#000000","pin-type-breadboard_ded8e15a-344e-4f93-a7cd-807af81d5cc8_0_3":"#000000","pin-type-breadboard_ded8e15a-344e-4f93-a7cd-807af81d5cc8_1_3":"#000000","pin-type-breadboard_ded8e15a-344e-4f93-a7cd-807af81d5cc8_0_4":"#000000","pin-type-breadboard_ded8e15a-344e-4f93-a7cd-807af81d5cc8_1_4":"#000000","pin-type-breadboard_ded8e15a-344e-4f93-a7cd-807af81d5cc8_0_5":"#000000","pin-type-breadboard_ded8e15a-344e-4f93-a7cd-807af81d5cc8_1_5":"#000000","pin-type-breadboard_ded8e15a-344e-4f93-a7cd-807af81d5cc8_0_6":"#000000","pin-type-breadboard_ded8e15a-344e-4f93-a7cd-807af81d5cc8_1_6":"#000000","pin-type-breadboard_ded8e15a-344e-4f93-a7cd-807af81d5cc8_0_7":"#000000","pin-type-breadboard_ded8e15a-344e-4f93-a7cd-807af81d5cc8_1_7":"#000000","pin-type-breadboard_ded8e15a-344e-4f93-a7cd-807af81d5cc8_0_8":"#000000","pin-type-breadboard_ded8e15a-344e-4f93-a7cd-807af81d5cc8_1_8":"#000000","pin-type-breadboard_ded8e15a-344e-4f93-a7cd-807af81d5cc8_0_9":"#000000","pin-type-breadboard_ded8e15a-344e-4f93-a7cd-807af81d5cc8_1_9":"#000000","pin-type-breadboard_ded8e15a-344e-4f93-a7cd-807af81d5cc8_0_10":"#000000","pin-type-breadboard_ded8e15a-344e-4f93-a7cd-807af81d5cc8_1_10":"#000000","pin-type-breadboard_ded8e15a-344e-4f93-a7cd-807af81d5cc8_0_11":"#000000","pin-type-breadboard_ded8e15a-344e-4f93-a7cd-807af81d5cc8_1_11":"#000000","pin-type-breadboard_ded8e15a-344e-4f93-a7cd-807af81d5cc8_0_12":"#000000","pin-type-breadboard_ded8e15a-344e-4f93-a7cd-807af81d5cc8_1_12":"#000000","pin-type-breadboard_ded8e15a-344e-4f93-a7cd-807af81d5cc8_0_13":"#000000","pin-type-breadboard_ded8e15a-344e-4f93-a7cd-807af81d5cc8_1_13":"#000000","pin-type-breadboard_ded8e15a-344e-4f93-a7cd-807af81d5cc8_0_14":"#000000","pin-type-breadboard_ded8e15a-344e-4f93-a7cd-807af81d5cc8_1_14":"#000000","pin-type-breadboard_ded8e15a-344e-4f93-a7cd-807af81d5cc8_0_15":"#000000","pin-type-breadboard_ded8e15a-344e-4f93-a7cd-807af81d5cc8_1_15":"#000000","pin-type-breadboard_ded8e15a-344e-4f93-a7cd-807af81d5cc8_0_16":"#000000","pin-type-breadboard_ded8e15a-344e-4f93-a7cd-807af81d5cc8_1_16":"#000000"},"pin_to_state":{"pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_0":"neutral","pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_1":"neutral","pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_2":"neutral","pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_3":"neutral","pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_4":"neutral","pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_5":"neutral","pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_6":"neutral","pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_7":"neutral","pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_8":"neutral","pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_10":"neutral","pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_11":"neutral","pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_12":"neutral","pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_13":"neutral","pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_14":"neutral","pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_16":"neutral","pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_18":"neutral","pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_19":"neutral","pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_20":"neutral","pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_21":"neutral","pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_22":"neutral","pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_23":"neutral","pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_24":"neutral","pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_25":"neutral","pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_27":"neutral","pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_28":"neutral","pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_29":"neutral","pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_30":"neutral","pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_31":"neutral","pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_32":"neutral","pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_33":"neutral","pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_34":"neutral","pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_35":"neutral","pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_36":"neutral","pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_37":"neutral","pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_38":"neutral","pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_39":"neutral","pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_40":"neutral","pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_41":"neutral","pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_15":"neutral","pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_17":"neutral","pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_9":"neutral","pin-type-component_68cda57c-349d-45e9-a6a2-98cf0cbc2416_0":"neutral","pin-type-component_68cda57c-349d-45e9-a6a2-98cf0cbc2416_1":"neutral","pin-type-component_68cda57c-349d-45e9-a6a2-98cf0cbc2416_2":"neutral","pin-type-component_68cda57c-349d-45e9-a6a2-98cf0cbc2416_3":"neutral","pin-type-component_68cda57c-349d-45e9-a6a2-98cf0cbc2416_4":"neutral","pin-type-component_68cda57c-349d-45e9-a6a2-98cf0cbc2416_5":"neutral","pin-type-component_68cda57c-349d-45e9-a6a2-98cf0cbc2416_6":"neutral","pin-type-component_68cda57c-349d-45e9-a6a2-98cf0cbc2416_7":"neutral","pin-type-component_68cda57c-349d-45e9-a6a2-98cf0cbc2416_8":"neutral","pin-type-component_68cda57c-349d-45e9-a6a2-98cf0cbc2416_9":"neutral","pin-type-component_68cda57c-349d-45e9-a6a2-98cf0cbc2416_10":"neutral","pin-type-component_68cda57c-349d-45e9-a6a2-98cf0cbc2416_11":"neutral","pin-type-component_68cda57c-349d-45e9-a6a2-98cf0cbc2416_12":"neutral","pin-type-component_68cda57c-349d-45e9-a6a2-98cf0cbc2416_13":"neutral","pin-type-component_68cda57c-349d-45e9-a6a2-98cf0cbc2416_14":"neutral","pin-type-component_68cda57c-349d-45e9-a6a2-98cf0cbc2416_15":"neutral","pin-type-component_68cda57c-349d-45e9-a6a2-98cf0cbc2416_16":"neutral","pin-type-component_fc7a62c0-bbca-4c4c-a089-8837f2378795_0":"neutral","pin-type-component_fc7a62c0-bbca-4c4c-a089-8837f2378795_1":"neutral","pin-type-component_c3c8c3f0-5cb8-46df-9e8e-6bc9ea246e79_0":"neutral","pin-type-component_c3c8c3f0-5cb8-46df-9e8e-6bc9ea246e79_1":"neutral","pin-type-component_db7d8f7f-8f6f-44a8-be93-8d8d7b68807d_0":"neutral","pin-type-component_db7d8f7f-8f6f-44a8-be93-8d8d7b68807d_1":"neutral","pin-type-breadboard_ded8e15a-344e-4f93-a7cd-807af81d5cc8_0_0":"neutral","pin-type-breadboard_ded8e15a-344e-4f93-a7cd-807af81d5cc8_1_0":"neutral","pin-type-breadboard_ded8e15a-344e-4f93-a7cd-807af81d5cc8_0_1":"neutral","pin-type-breadboard_ded8e15a-344e-4f93-a7cd-807af81d5cc8_1_1":"neutral","pin-type-breadboard_ded8e15a-344e-4f93-a7cd-807af81d5cc8_0_2":"neutral","pin-type-breadboard_ded8e15a-344e-4f93-a7cd-807af81d5cc8_1_2":"neutral","pin-type-breadboard_ded8e15a-344e-4f93-a7cd-807af81d5cc8_0_3":"neutral","pin-type-breadboard_ded8e15a-344e-4f93-a7cd-807af81d5cc8_1_3":"neutral","pin-type-breadboard_ded8e15a-344e-4f93-a7cd-807af81d5cc8_0_4":"neutral","pin-type-breadboard_ded8e15a-344e-4f93-a7cd-807af81d5cc8_1_4":"neutral","pin-type-breadboard_ded8e15a-344e-4f93-a7cd-807af81d5cc8_0_5":"neutral","pin-type-breadboard_ded8e15a-344e-4f93-a7cd-807af81d5cc8_1_5":"neutral","pin-type-breadboard_ded8e15a-344e-4f93-a7cd-807af81d5cc8_0_6":"neutral","pin-type-breadboard_ded8e15a-344e-4f93-a7cd-807af81d5cc8_1_6":"neutral","pin-type-breadboard_ded8e15a-344e-4f93-a7cd-807af81d5cc8_0_7":"neutral","pin-type-breadboard_ded8e15a-344e-4f93-a7cd-807af81d5cc8_1_7":"neutral","pin-type-breadboard_ded8e15a-344e-4f93-a7cd-807af81d5cc8_0_8":"neutral","pin-type-breadboard_ded8e15a-344e-4f93-a7cd-807af81d5cc8_1_8":"neutral","pin-type-breadboard_ded8e15a-344e-4f93-a7cd-807af81d5cc8_0_9":"neutral","pin-type-breadboard_ded8e15a-344e-4f93-a7cd-807af81d5cc8_1_9":"neutral","pin-type-breadboard_ded8e15a-344e-4f93-a7cd-807af81d5cc8_0_10":"neutral","pin-type-breadboard_ded8e15a-344e-4f93-a7cd-807af81d5cc8_1_10":"neutral","pin-type-breadboard_ded8e15a-344e-4f93-a7cd-807af81d5cc8_0_11":"neutral","pin-type-breadboard_ded8e15a-344e-4f93-a7cd-807af81d5cc8_1_11":"neutral","pin-type-breadboard_ded8e15a-344e-4f93-a7cd-807af81d5cc8_0_12":"neutral","pin-type-breadboard_ded8e15a-344e-4f93-a7cd-807af81d5cc8_1_12":"neutral","pin-type-breadboard_ded8e15a-344e-4f93-a7cd-807af81d5cc8_0_13":"neutral","pin-type-breadboard_ded8e15a-344e-4f93-a7cd-807af81d5cc8_1_13":"neutral","pin-type-breadboard_ded8e15a-344e-4f93-a7cd-807af81d5cc8_0_14":"neutral","pin-type-breadboard_ded8e15a-344e-4f93-a7cd-807af81d5cc8_1_14":"neutral","pin-type-breadboard_ded8e15a-344e-4f93-a7cd-807af81d5cc8_0_15":"neutral","pin-type-breadboard_ded8e15a-344e-4f93-a7cd-807af81d5cc8_1_15":"neutral","pin-type-breadboard_ded8e15a-344e-4f93-a7cd-807af81d5cc8_0_16":"neutral","pin-type-breadboard_ded8e15a-344e-4f93-a7cd-807af81d5cc8_1_16":"neutral"},"next_color_idx":14,"wires_placed_in_order":[["pin-type-component_db7d8f7f-8f6f-44a8-be93-8d8d7b68807d_1","pin-type-component_68cda57c-349d-45e9-a6a2-98cf0cbc2416_14"],["pin-type-component_db7d8f7f-8f6f-44a8-be93-8d8d7b68807d_0","pin-type-component_68cda57c-349d-45e9-a6a2-98cf0cbc2416_15"],["pin-type-component_fc7a62c0-bbca-4c4c-a089-8837f2378795_0","pin-type-component_68cda57c-349d-45e9-a6a2-98cf0cbc2416_8"],["pin-type-component_fc7a62c0-bbca-4c4c-a089-8837f2378795_0","pin-type-component_68cda57c-349d-45e9-a6a2-98cf0cbc2416_8"],["pin-type-component_fc7a62c0-bbca-4c4c-a089-8837f2378795_1","pin-type-component_68cda57c-349d-45e9-a6a2-98cf0cbc2416_9"],["pin-type-component_c3c8c3f0-5cb8-46df-9e8e-6bc9ea246e79_0","pin-type-component_68cda57c-349d-45e9-a6a2-98cf0cbc2416_7"],["pin-type-component_c3c8c3f0-5cb8-46df-9e8e-6bc9ea246e79_1","pin-type-component_68cda57c-349d-45e9-a6a2-98cf0cbc2416_6"],["pin-type-component_68cda57c-349d-45e9-a6a2-98cf0cbc2416_0","pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_16"],["pin-type-component_68cda57c-349d-45e9-a6a2-98cf0cbc2416_11","pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_24"],["pin-type-component_68cda57c-349d-45e9-a6a2-98cf0cbc2416_1","pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_27"],["pin-type-component_68cda57c-349d-45e9-a6a2-98cf0cbc2416_5","pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_28"],["pin-type-component_68cda57c-349d-45e9-a6a2-98cf0cbc2416_4","pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_10"],["pin-type-component_68cda57c-349d-45e9-a6a2-98cf0cbc2416_3","pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_40"],["pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_37","pin-type-breadboard_ded8e15a-344e-4f93-a7cd-807af81d5cc8_0_0"],["pin-type-breadboard_ded8e15a-344e-4f93-a7cd-807af81d5cc8_0_0","pin-type-component_68cda57c-349d-45e9-a6a2-98cf0cbc2416_15"]],"wires_removed_and_placed_in_order":[[[],[["pin-type-component_db7d8f7f-8f6f-44a8-be93-8d8d7b68807d_1","pin-type-component_68cda57c-349d-45e9-a6a2-98cf0cbc2416_14"]]],[[],[["pin-type-component_db7d8f7f-8f6f-44a8-be93-8d8d7b68807d_0","pin-type-component_68cda57c-349d-45e9-a6a2-98cf0cbc2416_15"]]],[[],[["pin-type-component_fc7a62c0-bbca-4c4c-a089-8837f2378795_0","pin-type-component_68cda57c-349d-45e9-a6a2-98cf0cbc2416_8"]]],[[["pin-type-component_68cda57c-349d-45e9-a6a2-98cf0cbc2416_8","pin-type-component_fc7a62c0-bbca-4c4c-a089-8837f2378795_0"]],[]],[[],[["pin-type-component_fc7a62c0-bbca-4c4c-a089-8837f2378795_0","pin-type-component_68cda57c-349d-45e9-a6a2-98cf0cbc2416_8"]]],[[],[["pin-type-component_fc7a62c0-bbca-4c4c-a089-8837f2378795_1","pin-type-component_68cda57c-349d-45e9-a6a2-98cf0cbc2416_9"]]],[[],[["pin-type-component_c3c8c3f0-5cb8-46df-9e8e-6bc9ea246e79_0","pin-type-component_68cda57c-349d-45e9-a6a2-98cf0cbc2416_7"]]],[[],[["pin-type-component_c3c8c3f0-5cb8-46df-9e8e-6bc9ea246e79_1","pin-type-component_68cda57c-349d-45e9-a6a2-98cf0cbc2416_6"]]],[[],[["pin-type-component_68cda57c-349d-45e9-a6a2-98cf0cbc2416_0","pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_16"]]],[[],[["pin-type-component_68cda57c-349d-45e9-a6a2-98cf0cbc2416_11","pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_24"]]],[[],[["pin-type-component_68cda57c-349d-45e9-a6a2-98cf0cbc2416_1","pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_27"]]],[[],[["pin-type-component_68cda57c-349d-45e9-a6a2-98cf0cbc2416_5","pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_28"]]],[[],[["pin-type-component_68cda57c-349d-45e9-a6a2-98cf0cbc2416_4","pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_10"]]],[[],[["pin-type-component_68cda57c-349d-45e9-a6a2-98cf0cbc2416_3","pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_40"]]],[[],[["pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_37","pin-type-breadboard_ded8e15a-344e-4f93-a7cd-807af81d5cc8_0_0"]]],[[],[["pin-type-breadboard_ded8e15a-344e-4f93-a7cd-807af81d5cc8_0_0","pin-type-component_68cda57c-349d-45e9-a6a2-98cf0cbc2416_15"]]]],"arduino_state":"arduino_off","pin_to_uid":{"pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_0":"_","pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_1":"_","pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_2":"_","pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_3":"_","pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_4":"_","pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_5":"_","pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_6":"_","pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_7":"_","pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_8":"_","pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_10":"0000000000000010","pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_11":"_","pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_12":"_","pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_13":"_","pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_14":"_","pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_16":"0000000000000006","pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_18":"_","pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_19":"_","pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_20":"_","pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_21":"_","pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_22":"_","pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_23":"_","pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_24":"0000000000000007","pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_25":"_","pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_27":"0000000000000008","pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_28":"0000000000000009","pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_29":"_","pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_30":"_","pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_31":"_","pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_32":"_","pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_33":"_","pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_34":"_","pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_35":"_","pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_36":"_","pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_37":"0000000000000001","pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_38":"_","pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_39":"_","pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_40":"0000000000000011","pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_41":"_","pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_15":"_","pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_17":"_","pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_9":"_","pin-type-component_68cda57c-349d-45e9-a6a2-98cf0cbc2416_0":"0000000000000006","pin-type-component_68cda57c-349d-45e9-a6a2-98cf0cbc2416_1":"0000000000000008","pin-type-component_68cda57c-349d-45e9-a6a2-98cf0cbc2416_2":"_","pin-type-component_68cda57c-349d-45e9-a6a2-98cf0cbc2416_3":"0000000000000011","pin-type-component_68cda57c-349d-45e9-a6a2-98cf0cbc2416_4":"0000000000000010","pin-type-component_68cda57c-349d-45e9-a6a2-98cf0cbc2416_5":"0000000000000009","pin-type-component_68cda57c-349d-45e9-a6a2-98cf0cbc2416_6":"0000000000000005","pin-type-component_68cda57c-349d-45e9-a6a2-98cf0cbc2416_7":"0000000000000004","pin-type-component_68cda57c-349d-45e9-a6a2-98cf0cbc2416_8":"0000000000000002","pin-type-component_68cda57c-349d-45e9-a6a2-98cf0cbc2416_9":"0000000000000003","pin-type-component_68cda57c-349d-45e9-a6a2-98cf0cbc2416_10":"_","pin-type-component_68cda57c-349d-45e9-a6a2-98cf0cbc2416_11":"0000000000000007","pin-type-component_68cda57c-349d-45e9-a6a2-98cf0cbc2416_12":"_","pin-type-component_68cda57c-349d-45e9-a6a2-98cf0cbc2416_13":"_","pin-type-component_68cda57c-349d-45e9-a6a2-98cf0cbc2416_14":"0000000000000000","pin-type-component_68cda57c-349d-45e9-a6a2-98cf0cbc2416_15":"0000000000000001","pin-type-component_68cda57c-349d-45e9-a6a2-98cf0cbc2416_16":"_","pin-type-component_fc7a62c0-bbca-4c4c-a089-8837f2378795_0":"0000000000000002","pin-type-component_fc7a62c0-bbca-4c4c-a089-8837f2378795_1":"0000000000000003","pin-type-component_c3c8c3f0-5cb8-46df-9e8e-6bc9ea246e79_0":"0000000000000004","pin-type-component_c3c8c3f0-5cb8-46df-9e8e-6bc9ea246e79_1":"0000000000000005","pin-type-component_db7d8f7f-8f6f-44a8-be93-8d8d7b68807d_0":"0000000000000001","pin-type-component_db7d8f7f-8f6f-44a8-be93-8d8d7b68807d_1":"0000000000000000","pin-type-breadboard_ded8e15a-344e-4f93-a7cd-807af81d5cc8_0_0":"0000000000000001","pin-type-breadboard_ded8e15a-344e-4f93-a7cd-807af81d5cc8_1_0":"_","pin-type-breadboard_ded8e15a-344e-4f93-a7cd-807af81d5cc8_0_1":"_","pin-type-breadboard_ded8e15a-344e-4f93-a7cd-807af81d5cc8_1_1":"_","pin-type-breadboard_ded8e15a-344e-4f93-a7cd-807af81d5cc8_0_2":"_","pin-type-breadboard_ded8e15a-344e-4f93-a7cd-807af81d5cc8_1_2":"_","pin-type-breadboard_ded8e15a-344e-4f93-a7cd-807af81d5cc8_0_3":"_","pin-type-breadboard_ded8e15a-344e-4f93-a7cd-807af81d5cc8_1_3":"_","pin-type-breadboard_ded8e15a-344e-4f93-a7cd-807af81d5cc8_0_4":"_","pin-type-breadboard_ded8e15a-344e-4f93-a7cd-807af81d5cc8_1_4":"_","pin-type-breadboard_ded8e15a-344e-4f93-a7cd-807af81d5cc8_0_5":"_","pin-type-breadboard_ded8e15a-344e-4f93-a7cd-807af81d5cc8_1_5":"_","pin-type-breadboard_ded8e15a-344e-4f93-a7cd-807af81d5cc8_0_6":"_","pin-type-breadboard_ded8e15a-344e-4f93-a7cd-807af81d5cc8_1_6":"_","pin-type-breadboard_ded8e15a-344e-4f93-a7cd-807af81d5cc8_0_7":"_","pin-type-breadboard_ded8e15a-344e-4f93-a7cd-807af81d5cc8_1_7":"_","pin-type-breadboard_ded8e15a-344e-4f93-a7cd-807af81d5cc8_0_8":"_","pin-type-breadboard_ded8e15a-344e-4f93-a7cd-807af81d5cc8_1_8":"_","pin-type-breadboard_ded8e15a-344e-4f93-a7cd-807af81d5cc8_0_9":"_","pin-type-breadboard_ded8e15a-344e-4f93-a7cd-807af81d5cc8_1_9":"_","pin-type-breadboard_ded8e15a-344e-4f93-a7cd-807af81d5cc8_0_10":"_","pin-type-breadboard_ded8e15a-344e-4f93-a7cd-807af81d5cc8_1_10":"_","pin-type-breadboard_ded8e15a-344e-4f93-a7cd-807af81d5cc8_0_11":"_","pin-type-breadboard_ded8e15a-344e-4f93-a7cd-807af81d5cc8_1_11":"_","pin-type-breadboard_ded8e15a-344e-4f93-a7cd-807af81d5cc8_0_12":"_","pin-type-breadboard_ded8e15a-344e-4f93-a7cd-807af81d5cc8_1_12":"_","pin-type-breadboard_ded8e15a-344e-4f93-a7cd-807af81d5cc8_0_13":"_","pin-type-breadboard_ded8e15a-344e-4f93-a7cd-807af81d5cc8_1_13":"_","pin-type-breadboard_ded8e15a-344e-4f93-a7cd-807af81d5cc8_0_14":"_","pin-type-breadboard_ded8e15a-344e-4f93-a7cd-807af81d5cc8_1_14":"_","pin-type-breadboard_ded8e15a-344e-4f93-a7cd-807af81d5cc8_0_15":"_","pin-type-breadboard_ded8e15a-344e-4f93-a7cd-807af81d5cc8_1_15":"_","pin-type-breadboard_ded8e15a-344e-4f93-a7cd-807af81d5cc8_0_16":"_","pin-type-breadboard_ded8e15a-344e-4f93-a7cd-807af81d5cc8_1_16":"_"},"component_id_to_pins":{"d590422c-57c9-4552-b8d5-f912e9490639":["0","1","2","3","4","5","6","7","8","10","11","12","13","14","16","18","19","20","21","22","23","24","25","27","28","29","30","31","32","33","34","35","36","37","38","39","40","41","15","17","9"],"68cda57c-349d-45e9-a6a2-98cf0cbc2416":["0","1","2","3","4","5","6","7","8","9","10","11","12","13","14","15","16"],"fc7a62c0-bbca-4c4c-a089-8837f2378795":["0","1"],"c3c8c3f0-5cb8-46df-9e8e-6bc9ea246e79":["0","1"],"db7d8f7f-8f6f-44a8-be93-8d8d7b68807d":["0","1"],"2dbc197b-6c39-4927-9244-ccf54552ff17":[]},"uid_to_net":{"_":[],"0000000000000000":["pin-type-component_db7d8f7f-8f6f-44a8-be93-8d8d7b68807d_1","pin-type-component_68cda57c-349d-45e9-a6a2-98cf0cbc2416_14"],"0000000000000001":["pin-type-breadboard_ded8e15a-344e-4f93-a7cd-807af81d5cc8_0_0","pin-type-component_68cda57c-349d-45e9-a6a2-98cf0cbc2416_15","pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_37","pin-type-component_db7d8f7f-8f6f-44a8-be93-8d8d7b68807d_0"],"0000000000000002":["pin-type-component_fc7a62c0-bbca-4c4c-a089-8837f2378795_0","pin-type-component_68cda57c-349d-45e9-a6a2-98cf0cbc2416_8"],"0000000000000003":["pin-type-component_fc7a62c0-bbca-4c4c-a089-8837f2378795_1","pin-type-component_68cda57c-349d-45e9-a6a2-98cf0cbc2416_9"],"0000000000000004":["pin-type-component_c3c8c3f0-5cb8-46df-9e8e-6bc9ea246e79_0","pin-type-component_68cda57c-349d-45e9-a6a2-98cf0cbc2416_7"],"0000000000000005":["pin-type-component_c3c8c3f0-5cb8-46df-9e8e-6bc9ea246e79_1","pin-type-component_68cda57c-349d-45e9-a6a2-98cf0cbc2416_6"],"0000000000000006":["pin-type-component_68cda57c-349d-45e9-a6a2-98cf0cbc2416_0","pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_16"],"0000000000000007":["pin-type-component_68cda57c-349d-45e9-a6a2-98cf0cbc2416_11","pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_24"],"0000000000000008":["pin-type-component_68cda57c-349d-45e9-a6a2-98cf0cbc2416_1","pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_27"],"0000000000000009":["pin-type-component_68cda57c-349d-45e9-a6a2-98cf0cbc2416_5","pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_28"],"0000000000000010":["pin-type-component_68cda57c-349d-45e9-a6a2-98cf0cbc2416_4","pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_10"],"0000000000000011":["pin-type-component_68cda57c-349d-45e9-a6a2-98cf0cbc2416_3","pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_40"]},"uid_to_text_label":{"0000000000000000":"Net 0","0000000000000001":"Net 1","0000000000000002":"Net 2","0000000000000003":"Net 3","0000000000000004":"Net 4","0000000000000005":"Net 5","0000000000000006":"Net 6","0000000000000007":"Net 7","0000000000000008":"Net 8","0000000000000009":"Net 9","0000000000000010":"Net 10","0000000000000011":"Net 11"},"all_breadboard_info_list":["44ff7df1-4fd5-4980-a165-c1dce7a13984_17_2_False_99.99999999999999_1210_up","ded8e15a-344e-4f93-a7cd-807af81d5cc8_17_2_False_1375_1105_up"],"breadboard_info_list":["ded8e15a-344e-4f93-a7cd-807af81d5cc8_17_2_False_1375_1105_up"],"componentsData":[{"compProperties":{"mpn":{"version":2,"id":"mpn","label":"mpn","description":"","units":"","type":"string","value":"RPI3-MODB-16GB-NOOBS","displayFormat":"input","showOnComp":false,"isVisibleToUser":false,"name":"mpn","unit":"","userVisible":false,"required":true},"manufacturer":{"version":2,"id":"manufacturer","label":"manufacturer","description":"","units":"","type":"string","value":"Raspberry Pi","displayFormat":"input","showOnComp":false,"isVisibleToUser":false,"name":"manufacturer","unit":"","userVisible":false,"required":true}},"position":[1124.31025,675.44717],"typeId":"9d987227-334c-49a7-9e0b-80422ab638f6","componentVersion":2,"instanceId":"d590422c-57c9-4552-b8d5-f912e9490639","orientation":"up","circleData":[[917.5,530],[932.5,530],[947.5,530],[962.5,530],[977.5,530],[992.5,530],[1007.5,530],[1022.5,530],[1037.5,530],[1067.5,530],[1082.5,530],[1097.5,530],[1112.5,530],[1127.5,530],[1157.5,530],[1187.5,530],[1202.5,530],[1202.5,515],[1187.5,515],[1172.5,515],[1157.5,515],[1142.5,515],[1127.5,515],[1097.5,515],[1082.5,515],[1067.5,515],[1052.5,515],[1037.5,515],[1022.5,515],[1007.5,515],[992.5,515],[977.5,515],[962.5,515],[947.5,515],[932.5,515],[917.5,515],[1052.5,530],[1112.5,515],[1142.5,530],[1172.5,530],[931.6614999999999,831.6770000000001]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[1120.014031,973.1704910000001],"typeId":"8313da4d-6f61-4c01-9e39-e2529c7db0e0","componentVersion":2,"instanceId":"68cda57c-349d-45e9-a6a2-98cf0cbc2416","orientation":"up","circleData":[[1127.4999999999998,1025],[1133.2827054999998,1024.7128805000002],[1126.3984944999997,1018.5881810000002],[1154.3614914999998,1025.138849],[1146.9980364999997,1024.8784955],[1140.3513924999997,1024.8784955],[1169.9854675000001,985.0851395000001],[1170.1263670000003,998.0436395],[1070.3230749999998,987.474722],[1070.0272705,1000.8686270000001],[1162.138144,1018.66511],[1162.0341325,1025.3306315],[1103.3235969999998,998.7550430000001],[1094.5070199999998,998.9065805000001],[1084.6546795,1022.9627015000001],[1098.4100019999998,1022.9627015000001],[1111.3293909999998,1022.9260924999999]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[793.9273495,975.6876065000001],"typeId":"7115dd0c-9076-1603-96e1-f4f66aa483df","componentVersion":7,"instanceId":"fc7a62c0-bbca-4c4c-a089-8837f2378795","orientation":"down","circleData":[[977.5,1025],[977.5,926.162]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"mpn":{"version":2,"id":"mpn","label":"mpn","description":"","units":"","type":"string","value":"3858","displayFormat":"input","showOnComp":false,"isVisibleToUser":false,"name":"mpn","unit":"","userVisible":false,"required":true},"manufacturer":{"version":2,"id":"manufacturer","label":"manufacturer","description":"","units":"","type":"string","value":"Adafruit Industries","displayFormat":"input","showOnComp":false,"isVisibleToUser":false,"name":"manufacturer","unit":"","userVisible":false,"required":true}},"position":[1134.2763234999998,1345.9301645],"typeId":"70e5c902-d992-f164-9b8f-2034db0ec022","componentVersion":1,"instanceId":"db7d8f7f-8f6f-44a8-be93-8d8d7b68807d","orientation":"left","circleData":[[1142.5,1160],[1112.5,1160]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[1431.0726505,969.3123935000006],"typeId":"7115dd0c-9076-1603-96e1-f4f66aa483df","componentVersion":7,"instanceId":"c3c8c3f0-5cb8-46df-9e8e-6bc9ea246e79","orientation":"up","circleData":[[1247.5,920],[1247.5,1018.8379999999999]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"Comment":{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"L298N and DC hobby motor wires and pins:\n\n  Red wires - IN1, IN3\n  Black wires - IN2, IN4\n\n  IN1, IN2 = GPIO7, GPIO8\n  IN3, IN4 = GPIO9, GPIO10\n  ENA, ENB = GPIO13, GPIO12\n\n  12+V (VC) - Connect to Power Supply Battery 2x3.7V\n  GND - GND\n  5+V (VCC) - no need to connect to it \n            since DC motors require 6V each\n  \nNOTE: Both RPi and L298N must have a common ground!\n Connect RPi GND to L298N GND powered from battery","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"backgroundColor":{"version":2,"id":"backgroundColor","label":"Background Color","description":"","units":"","type":"string","value":"#ffffff","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"backgroundOpacity":{"version":2,"id":"backgroundOpacity","label":"Background Opacity","description":"","units":"","type":"decimal","value":"1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"textColor":{"version":2,"id":"textColor","label":"Text Color","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"fontSize":{"version":2,"id":"fontSize","label":"Font Size","description":"","units":"","type":"integer","value":"12","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"font":{"version":2,"id":"font","label":"Font","description":"","units":"","type":"string","value":"Arial","displayFormat":"input","showOnComp":false,"isVisibleToUser":true}},"position":[1595.77707889522,765.953930383508],"typeId":"9a5a4baa-44d4-4aa0-8d82-488487322b20","componentVersion":1,"instanceId":"2dbc197b-6c39-4927-9244-ccf54552ff17","orientation":"up","circleData":[],"cirkitStudioVersion":"1.3.3"}],"bounds":{"top":"494.26042","left":"582.40160","width":"1188.39013","height":"1035.79574","x":"582.40160","y":"494.26042"},"cachedBreadboardPrettyViewWires":["{\"color\":\"#ff2600\",\"startPinId\":\"pin-type-component_68cda57c-349d-45e9-a6a2-98cf0cbc2416_14\",\"endPinId\":\"pin-type-component_db7d8f7f-8f6f-44a8-be93-8d8d7b68807d_1\",\"rawStartPinId\":\"pin-type-component_68cda57c-349d-45e9-a6a2-98cf0cbc2416_14\",\"rawEndPinId\":\"pin-type-component_db7d8f7f-8f6f-44a8-be93-8d8d7b68807d_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1084.6546795000_1022.9627015000\\\",\\\"1084.6546795000_1085.0000000000\\\",\\\"1112.5000000000_1085.0000000000\\\",\\\"1112.5000000000_1160.0000000000\\\"]}\"}","{\"color\":\"#000000\",\"startPinId\":\"pin-type-component_68cda57c-349d-45e9-a6a2-98cf0cbc2416_15\",\"endPinId\":\"pin-type-component_db7d8f7f-8f6f-44a8-be93-8d8d7b68807d_0\",\"rawStartPinId\":\"pin-type-component_68cda57c-349d-45e9-a6a2-98cf0cbc2416_15\",\"rawEndPinId\":\"pin-type-component_db7d8f7f-8f6f-44a8-be93-8d8d7b68807d_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1098.4100020000_1022.9627015000\\\",\\\"1098.4100020000_1070.0000000000\\\",\\\"1210.0000000000_1070.0000000000\\\",\\\"1210.0000000000_1160.0000000000\\\",\\\"1142.5000000000_1160.0000000000\\\"]}\"}","{\"color\":\"#000000\",\"startPinId\":\"pin-type-breadboard_ded8e15a-344e-4f93-a7cd-807af81d5cc8_0_0\",\"endPinId\":\"pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_37\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_ded8e15a-344e-4f93-a7cd-807af81d5cc8_0_0_4\",\"rawEndPinId\":\"pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_37\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1397.5000000000_1115.0000000000\\\",\\\"1397.5000000000_485.0000000000\\\",\\\"947.5000000000_485.0000000000\\\",\\\"947.5000000000_515.0000000000\\\"]}\"}","{\"color\":\"#000000\",\"startPinId\":\"pin-type-breadboard_ded8e15a-344e-4f93-a7cd-807af81d5cc8_0_0\",\"endPinId\":\"pin-type-component_68cda57c-349d-45e9-a6a2-98cf0cbc2416_15\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_ded8e15a-344e-4f93-a7cd-807af81d5cc8_0_0_0\",\"rawEndPinId\":\"pin-type-component_68cda57c-349d-45e9-a6a2-98cf0cbc2416_15\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1337.5000000000_1115.0000000000\\\",\\\"1337.5000000000_1047.5000000000\\\",\\\"1097.5000000000_1047.5000000000\\\",\\\"1097.5000000000_1022.9627015000\\\",\\\"1098.4100020000_1022.9627015000\\\"]}\"}","{\"color\":\"#ff2600\",\"startPinId\":\"pin-type-component_68cda57c-349d-45e9-a6a2-98cf0cbc2416_8\",\"endPinId\":\"pin-type-component_fc7a62c0-bbca-4c4c-a089-8837f2378795_0\",\"rawStartPinId\":\"pin-type-component_68cda57c-349d-45e9-a6a2-98cf0cbc2416_8\",\"rawEndPinId\":\"pin-type-component_fc7a62c0-bbca-4c4c-a089-8837f2378795_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1070.3230750000_987.4747220000\\\",\\\"1022.5000000000_987.4747220000\\\",\\\"1022.5000000000_1025.0000000000\\\",\\\"977.5000000000_1025.0000000000\\\"]}\"}","{\"color\":\"#000000\",\"startPinId\":\"pin-type-component_68cda57c-349d-45e9-a6a2-98cf0cbc2416_9\",\"endPinId\":\"pin-type-component_fc7a62c0-bbca-4c4c-a089-8837f2378795_1\",\"rawStartPinId\":\"pin-type-component_68cda57c-349d-45e9-a6a2-98cf0cbc2416_9\",\"rawEndPinId\":\"pin-type-component_fc7a62c0-bbca-4c4c-a089-8837f2378795_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1070.0272705000_1000.8686270000\\\",\\\"1045.0000000000_1000.8686270000\\\",\\\"1045.0000000000_926.1620000000\\\",\\\"977.5000000000_926.1620000000\\\"]}\"}","{\"color\":\"#ff2600\",\"startPinId\":\"pin-type-component_68cda57c-349d-45e9-a6a2-98cf0cbc2416_7\",\"endPinId\":\"pin-type-component_c3c8c3f0-5cb8-46df-9e8e-6bc9ea246e79_0\",\"rawStartPinId\":\"pin-type-component_68cda57c-349d-45e9-a6a2-98cf0cbc2416_7\",\"rawEndPinId\":\"pin-type-component_c3c8c3f0-5cb8-46df-9e8e-6bc9ea246e79_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1170.1263670000_998.0436395000\\\",\\\"1217.5000000000_998.0436395000\\\",\\\"1217.5000000000_920.0000000000\\\",\\\"1247.5000000000_920.0000000000\\\"]}\"}","{\"color\":\"#000000\",\"startPinId\":\"pin-type-component_68cda57c-349d-45e9-a6a2-98cf0cbc2416_6\",\"endPinId\":\"pin-type-component_c3c8c3f0-5cb8-46df-9e8e-6bc9ea246e79_1\",\"rawStartPinId\":\"pin-type-component_68cda57c-349d-45e9-a6a2-98cf0cbc2416_6\",\"rawEndPinId\":\"pin-type-component_c3c8c3f0-5cb8-46df-9e8e-6bc9ea246e79_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1169.9854675000_985.0851395000\\\",\\\"1169.9854675000_1017.5000000000\\\",\\\"1247.5000000000_1017.5000000000\\\",\\\"1247.5000000000_1018.8380000000\\\"]}\"}","{\"color\":\"#00f900\",\"startPinId\":\"pin-type-component_68cda57c-349d-45e9-a6a2-98cf0cbc2416_0\",\"endPinId\":\"pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_16\",\"rawStartPinId\":\"pin-type-component_68cda57c-349d-45e9-a6a2-98cf0cbc2416_0\",\"rawEndPinId\":\"pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_16\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1127.5000000000_1025.0000000000\\\",\\\"1127.5000000000_1062.5000000000\\\",\\\"850.0000000000_1062.5000000000\\\",\\\"850.0000000000_470.0000000000\\\",\\\"1157.5000000000_470.0000000000\\\",\\\"1157.5000000000_530.0000000000\\\"]}\"}","{\"color\":\"#874efe\",\"startPinId\":\"pin-type-component_68cda57c-349d-45e9-a6a2-98cf0cbc2416_11\",\"endPinId\":\"pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_24\",\"rawStartPinId\":\"pin-type-component_68cda57c-349d-45e9-a6a2-98cf0cbc2416_11\",\"rawEndPinId\":\"pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_24\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1162.0341325000_1025.3306315000\\\",\\\"1162.0341325000_1137.5000000000\\\",\\\"775.0000000000_1137.5000000000\\\",\\\"775.0000000000_395.0000000000\\\",\\\"1142.5000000000_395.0000000000\\\",\\\"1142.5000000000_515.0000000000\\\"]}\"}","{\"color\":\"#fffb00\",\"startPinId\":\"pin-type-component_68cda57c-349d-45e9-a6a2-98cf0cbc2416_1\",\"endPinId\":\"pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_27\",\"rawStartPinId\":\"pin-type-component_68cda57c-349d-45e9-a6a2-98cf0cbc2416_1\",\"rawEndPinId\":\"pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_27\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1133.2827055000_1024.7128805000\\\",\\\"1133.2827055000_1077.5000000000\\\",\\\"835.0000000000_1077.5000000000\\\",\\\"835.0000000000_455.0000000000\\\",\\\"1097.5000000000_455.0000000000\\\",\\\"1097.5000000000_515.0000000000\\\"]}\"}","{\"color\":\"#ff9300\",\"startPinId\":\"pin-type-component_68cda57c-349d-45e9-a6a2-98cf0cbc2416_5\",\"endPinId\":\"pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_28\",\"rawStartPinId\":\"pin-type-component_68cda57c-349d-45e9-a6a2-98cf0cbc2416_5\",\"rawEndPinId\":\"pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_28\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1140.3513925000_1024.8784955000\\\",\\\"1140.3513925000_1092.5000000000\\\",\\\"820.0000000000_1092.5000000000\\\",\\\"820.0000000000_440.0000000000\\\",\\\"1082.5000000000_440.0000000000\\\",\\\"1082.5000000000_515.0000000000\\\"]}\"}","{\"color\":\"#ff2600\",\"startPinId\":\"pin-type-component_68cda57c-349d-45e9-a6a2-98cf0cbc2416_4\",\"endPinId\":\"pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_10\",\"rawStartPinId\":\"pin-type-component_68cda57c-349d-45e9-a6a2-98cf0cbc2416_4\",\"rawEndPinId\":\"pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_10\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1146.9980365000_1024.8784955000\\\",\\\"1146.9980365000_1107.5000000000\\\",\\\"805.0000000000_1107.5000000000\\\",\\\"805.0000000000_425.0000000000\\\",\\\"1067.5000000000_425.0000000000\\\",\\\"1067.5000000000_530.0000000000\\\"]}\"}","{\"color\":\"#aa7942\",\"startPinId\":\"pin-type-component_68cda57c-349d-45e9-a6a2-98cf0cbc2416_3\",\"endPinId\":\"pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_40\",\"rawStartPinId\":\"pin-type-component_68cda57c-349d-45e9-a6a2-98cf0cbc2416_3\",\"rawEndPinId\":\"pin-type-component_d590422c-57c9-4552-b8d5-f912e9490639_40\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1154.3614915000_1025.1388490000\\\",\\\"1154.3614915000_1122.5000000000\\\",\\\"790.0000000000_1122.5000000000\\\",\\\"790.0000000000_410.0000000000\\\",\\\"1052.5000000000_410.0000000000\\\",\\\"1052.5000000000_530.0000000000\\\"]}\"}"],"projectDescription":""}PK
     �k�[               jsons/PK
     �k�[ċ�C+  +     jsons/user_defined.json{"type":"user_defined","version":"0.0.1","subtypes":[{"subtypeName":"Raspberry Pi 3B","category":["User Defined"],"userDefined":true,"id":"9d987227-334c-49a7-9e0b-80422ab638f6","subtypeDescription":"","subtypePic":"67df6019-bb76-4308-bacd-6454b246d44a.png","pinInfo":{"numDisplayCols":"34.16220","numDisplayRows":"22.82490","pins":[{"uniquePinIdString":"0","positionMil":"329.37500,2110.89280","isAnchorPin":true,"label":"1"},{"uniquePinIdString":"1","positionMil":"429.37500,2110.89280","isAnchorPin":false,"label":"3"},{"uniquePinIdString":"2","positionMil":"529.37500,2110.89280","isAnchorPin":false,"label":"5"},{"uniquePinIdString":"3","positionMil":"629.37500,2110.89280","isAnchorPin":false,"label":"7"},{"uniquePinIdString":"4","positionMil":"729.37500,2110.89280","isAnchorPin":false,"label":"9"},{"uniquePinIdString":"5","positionMil":"829.37500,2110.89280","isAnchorPin":false,"label":"11"},{"uniquePinIdString":"6","positionMil":"929.37500,2110.89280","isAnchorPin":false,"label":"13"},{"uniquePinIdString":"7","positionMil":"1029.37500,2110.89280","isAnchorPin":false,"label":"15"},{"uniquePinIdString":"8","positionMil":"1129.37500,2110.89280","isAnchorPin":false,"label":"17"},{"uniquePinIdString":"10","positionMil":"1329.37500,2110.89280","isAnchorPin":false,"label":"21"},{"uniquePinIdString":"11","positionMil":"1429.37500,2110.89280","isAnchorPin":false,"label":"23"},{"uniquePinIdString":"12","positionMil":"1529.37500,2110.89280","isAnchorPin":false,"label":"25"},{"uniquePinIdString":"13","positionMil":"1629.37500,2110.89280","isAnchorPin":false,"label":"27"},{"uniquePinIdString":"14","positionMil":"1729.37500,2110.89280","isAnchorPin":false,"label":"29"},{"uniquePinIdString":"16","positionMil":"1929.37500,2110.89280","isAnchorPin":false,"label":"33"},{"uniquePinIdString":"18","positionMil":"2129.37500,2110.89280","isAnchorPin":false,"label":"37"},{"uniquePinIdString":"19","positionMil":"2229.37500,2110.89280","isAnchorPin":false,"label":"39"},{"uniquePinIdString":"20","positionMil":"2229.37500,2210.89280","isAnchorPin":false,"label":"40"},{"uniquePinIdString":"21","positionMil":"2129.37500,2210.89280","isAnchorPin":false,"label":"38"},{"uniquePinIdString":"22","positionMil":"2029.37500,2210.89280","isAnchorPin":false,"label":"36"},{"uniquePinIdString":"23","positionMil":"1929.37500,2210.89280","isAnchorPin":false,"label":"34"},{"uniquePinIdString":"24","positionMil":"1829.37500,2210.89280","isAnchorPin":false,"label":"32"},{"uniquePinIdString":"25","positionMil":"1729.37500,2210.89280","isAnchorPin":false,"label":"30"},{"uniquePinIdString":"27","positionMil":"1529.37500,2210.89280","isAnchorPin":false,"label":"26"},{"uniquePinIdString":"28","positionMil":"1429.37500,2210.89280","isAnchorPin":false,"label":"24"},{"uniquePinIdString":"29","positionMil":"1329.37500,2210.89280","isAnchorPin":false,"label":"22"},{"uniquePinIdString":"30","positionMil":"1229.37500,2210.89280","isAnchorPin":false,"label":"20"},{"uniquePinIdString":"31","positionMil":"1129.37500,2210.89280","isAnchorPin":false,"label":"18"},{"uniquePinIdString":"32","positionMil":"1029.37500,2210.89280","isAnchorPin":false,"label":"16"},{"uniquePinIdString":"33","positionMil":"929.37500,2210.89280","isAnchorPin":false,"label":"14"},{"uniquePinIdString":"34","positionMil":"829.37500,2210.89280","isAnchorPin":false,"label":"12"},{"uniquePinIdString":"35","positionMil":"729.37500,2210.89280","isAnchorPin":false,"label":"10"},{"uniquePinIdString":"36","positionMil":"629.37500,2210.89280","isAnchorPin":false,"label":"8"},{"uniquePinIdString":"37","positionMil":"529.37500,2210.89280","isAnchorPin":false,"label":"6"},{"uniquePinIdString":"38","positionMil":"429.37500,2210.89280","isAnchorPin":false,"label":"4"},{"uniquePinIdString":"39","positionMil":"329.37500,2210.89280","isAnchorPin":false,"label":"2(5V)"},{"uniquePinIdString":"40","positionMil":"1229.37500,2110.89280","isAnchorPin":false,"label":"19"},{"uniquePinIdString":"41","positionMil":"1629.37500,2210.89280","isAnchorPin":false,"label":"28"},{"uniquePinIdString":"15","positionMil":"1829.37500,2110.89280","isAnchorPin":false,"label":"31"},{"uniquePinIdString":"17","positionMil":"2029.37500,2110.89280","isAnchorPin":false,"label":"35"},{"uniquePinIdString":"9","positionMil":"423.78500,99.71280","isAnchorPin":false,"label":"Power"}],"pinType":"wired"},"properties":[{"type":"string","name":"mpn","value":"RPI3-MODB-16GB-NOOBS","unit":"","showOnComp":false,"userVisible":false,"required":true},{"type":"string","name":"manufacturer","value":"Raspberry Pi","unit":"","showOnComp":false,"userVisible":false,"required":true}],"iconPic":"7de8bea6-aec6-4ad5-83ac-8e47725efc1f.png","componentVersion":2,"imageLocation":"local_cache","hasComponentImageSvg":false,"componentImageSvgUrl":""},{"subtypeName":"ln298","category":["User Defined"],"id":"8313da4d-6f61-4c01-9e39-e2529c7db0e0","componentVersion":2,"userDefined":true,"subtypeDescription":"","subtypePic":"89718c7b-e32a-4492-aa2b-d7960b76d502.png","iconPic":"8883793e-4c9f-4ae6-b420-3a6e91b2597d.png","hasComponentImageSvg":false,"componentImageSvgUrl":"","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"8.07107","numDisplayRows":"8.07107","pins":[{"uniquePinIdString":"0","positionMil":"453.45996,58.02344","isAnchorPin":true,"label":"ena"},{"uniquePinIdString":"1","positionMil":"492.01133,59.93757","isAnchorPin":false,"label":"in1"},{"uniquePinIdString":"2","positionMil":"446.11659,100.76890","isAnchorPin":false,"label":"5v"},{"uniquePinIdString":"3","positionMil":"632.53657,57.09778","isAnchorPin":false,"label":"in4"},{"uniquePinIdString":"4","positionMil":"583.44687,58.83347","isAnchorPin":false,"label":"in3"},{"uniquePinIdString":"5","positionMil":"539.13591,58.83347","isAnchorPin":false,"label":"in2"},{"uniquePinIdString":"6","positionMil":"736.69641,324.12251","isAnchorPin":false,"label":"out4"},{"uniquePinIdString":"7","positionMil":"737.63574,237.73251","isAnchorPin":false,"label":"out3"},{"uniquePinIdString":"8","positionMil":"72.28046,308.19196","isAnchorPin":false,"label":"out1"},{"uniquePinIdString":"9","positionMil":"70.30843,218.89926","isAnchorPin":false,"label":"out2"},{"uniquePinIdString":"10","positionMil":"684.38092,100.25604","isAnchorPin":false,"label":"5v"},{"uniquePinIdString":"11","positionMil":"683.68751,55.81923","isAnchorPin":false,"label":"enb"},{"uniquePinIdString":"12","positionMil":"292.28394,232.98982","isAnchorPin":false,"label":"gnd"},{"uniquePinIdString":"13","positionMil":"233.50676,231.97957","isAnchorPin":false,"label":"12v"},{"uniquePinIdString":"14","positionMil":"167.82449,71.60543","isAnchorPin":false,"label":"12v"},{"uniquePinIdString":"15","positionMil":"259.52664,71.60543","isAnchorPin":false,"label":"gnd"},{"uniquePinIdString":"16","positionMil":"345.65590,71.84949","isAnchorPin":false,"label":"5v"}],"pinType":"wired"},"properties":[],"propertiesV2":[]},{"subtypeName":"DC Gear Motor (3-6V)","category":["User Defined"],"userDefined":true,"id":"7115dd0c-9076-1603-96e1-f4f66aa483df","subtypeDescription":"","subtypePic":"e2e2c934-b375-45fc-834c-534243cbf361.png","iconPic":"6c1978d3-8c4d-4ea9-a1ba-37ab4b096c5d.png","imageLocation":"local_cache","componentVersion":7,"pinInfo":{"numDisplayCols":"26.87010","numDisplayRows":"12.94650","pins":[{"uniquePinIdString":"0","positionMil":"119.68733,976.07429","isAnchorPin":true,"label":"V+"},{"uniquePinIdString":"1","positionMil":"119.68733,317.15429","isAnchorPin":false,"label":"V-"}],"pinType":"wired"},"properties":[],"hasComponentImageSvg":true,"componentImageSvgUrl":"https://abacasstorageaccnt.blob.core.windows.net/cirkit/7f9ce5f4-cc5c-40e6-be98-a947128d0a84.svg","propertiesV2":[]},{"subtypeName":"2 x AA Battery Mount","category":["Power"],"userDefined":false,"id":"70e5c902-d992-f164-9b8f-2034db0ec022","subtypeDescription":"","subtypePic":"f87b1235-301d-4eff-8a86-0c2fbb955692.png","iconPic":"2832311d-4ed1-4369-9d2b-9063d9d0cda0.png","pinInfo":{"numDisplayCols":"23.21680","numDisplayRows":"12.15000","pins":[{"uniquePinIdString":"0","startPositionMil":"2321.68000,552.67549","endPositionMil":"2400.37443,552.67549","isAnchorPin":true,"label":"-"},{"uniquePinIdString":"1","startPositionMil":"2321.68000,742.82175","endPositionMil":"2400.37443,742.82175","isAnchorPin":false,"label":"+"}],"pinType":"movable"},"properties":[{"type":"string","name":"mpn","value":"3858","unit":"","showOnComp":false,"userVisible":false,"required":true},{"type":"string","name":"manufacturer","value":"Adafruit Industries","unit":"","showOnComp":false,"userVisible":false,"required":true}],"componentVersion":1,"imageLocation":"local_cache","hasComponentImageSvg":false,"componentImageSvgUrl":""},{"subtypeName":"DC Gear Motor (3-6V)","category":["User Defined"],"userDefined":true,"id":"7115dd0c-9076-1603-96e1-f4f66aa483df","subtypeDescription":"","subtypePic":"e2e2c934-b375-45fc-834c-534243cbf361.png","iconPic":"6c1978d3-8c4d-4ea9-a1ba-37ab4b096c5d.png","imageLocation":"local_cache","componentVersion":7,"pinInfo":{"numDisplayCols":"26.87010","numDisplayRows":"12.94650","pins":[{"uniquePinIdString":"0","positionMil":"119.68733,976.07429","isAnchorPin":true,"label":"V+"},{"uniquePinIdString":"1","positionMil":"119.68733,317.15429","isAnchorPin":false,"label":"V-"}],"pinType":"wired"},"properties":[],"hasComponentImageSvg":true,"componentImageSvgUrl":"https://abacasstorageaccnt.blob.core.windows.net/cirkit/7f9ce5f4-cc5c-40e6-be98-a947128d0a84.svg","propertiesV2":[]},{"subtypeName":"Comment V2","category":["User Defined"],"componentClass":"textbox","userDefined":true,"id":"9a5a4baa-44d4-4aa0-8d82-488487322b20","subtypeDescription":"","subtypePic":"c88b2895-5e8b-4a57-9f9a-b80dd50058b1.png","pinInfo":{"numPins":"0","polarity":[],"pinType":"movable"},"properties":[{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"text box (click to edit)","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"backgroundColor","label":"Background Color","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"backgroundOpacity","label":"Background Opacity","description":"","units":"","type":"decimal","value":"1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"textColor","label":"Text Color","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"fontSize","label":"Font Size","description":"","units":"","type":"integer","value":"10","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"font","label":"Font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true}],"iconPic":"d3694a2e-5bba-40c3-8069-8db85c4c9209.png","componentVersion":1,"imageLocation":"local_cache","propertiesV2":[],"hasComponentImageSvg":false,"componentImageSvgUrl":""}]}PK
     �k�[               images/PK
     �k�[����^� ^� /   images/67df6019-bb76-4308-bacd-6454b246d44a.png�PNG

   IHDR  �  �   vEj�   	pHYs  �  ���R/   �eXIfII*            (           V       ^   1 
   f   i�    p       �     �     ezgif.com  �       �    �  �    �      �w��  �iTXtXML:com.adobe.xmp     <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="XMP Core 6.0.0">
   <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#">
      <rdf:Description rdf:about=""
            xmlns:tiff="http://ns.adobe.com/tiff/1.0/"
            xmlns:xmp="http://ns.adobe.com/xap/1.0/">
         <tiff:Orientation>1</tiff:Orientation>
         <xmp:CreatorTool>ezgif.com</xmp:CreatorTool>
      </rdf:Description>
   </rdf:RDF>
</x:xmpmeta>
�[n  ��IDATx���	|]gy�����w�ڭ}�-/��@B��B�Z��RJJ��a銁N�$$��t���@[�a�RJ
ek�eŉ�Œ-/�"˖Y�,k�s�׉IKbk��9�����J�%ٺ����<�'Q�z�T����g(K!�ُ���l	έ���                      ��	hI˺��{WԜ�Ҵ�'��mJ�:���gp=�b��L �E�(A��{5�V���˜'�|�v�s��ޞQ��d`��o�                       ���O�?+�m��v���lS7ކt�y{���#Z�Qe�$�2@l�êtv�έM�.����_��Q�ݩ?W�n                       ��fk��g3���=�y�иs�����񧝷���l�Դ DA1�d����Q������p7)�����ʻ�9��                       ���l�v�7�	�m��8��;�>���9�[�� �A1~���T�6;;�;;��5�lR�s�z LH                        �U��v�� ��p^�;�_!�@Yڭ���5#(�OL0L��ԲM�2�0Ζ@                        ��Rg�K!g3f��������?(K�کeX1�b��A�*�W8���l�tv�)7ҵ                        �!K&!�l��5�)=�o+�ojI_ӧ5! 7EP��<�$g��
g��Fgg��#U                       ���V��[��?��9����}UOhP ~A1^�SA��Ev�O;)rn                       �A���*`��k����_VH_�c:  A1n��p���|��ى                       �]�B�����7Bc�=���A1n�*Ի4��wޫ                        ı�1f{H�S@�ղ��'tU@�!(�v*��z�s�g��&g��                       �\�ἾCA}F;�E���Q=% NHK;T��ޭ��yo�                        p+9�����m�~����2�E�Ԭ #(&�g'�s�g�w                        �F�
9ی��C��J�'��N	�!BJ�'��u��sy�s�.                        \r����_�}�y������A1��S�����C��,                        DJ����l�j��NA}J��{|���Hy@I��;5��v�+                        �%�lwk����ۿ���mFPL��tv��S
�:��	                        �Ћ����}S��=��<���py6 fF���                         7y���fc���Փ<���pxX�׌>���                        7{��է����}ZGx A1���c
�.                       �+���6%�MzH�D��ь #(f->�\������^�i	)�IJw�e'�)˹���no'���1R�IJ^�;�;�-jqyɾyiN�PHˡe�.]�3o��hzqV3�Wu�y{i����В                 x��`��q75�ٶ�ݹ���)	I
8/���s�	JM��n����P@���`߿�4�n���U�vnyA�LM����g�׸/��W5��       DT�z�����ǔ�?�N-p!�bVc���������{E%U�����<��>��9��:ϵ'�	1��f�����]�����漽v��m�^ԅ��                �G0TAr֍�v��G�s� T3�4��uq�Θ��g��O_���W/����g�`U      ��Fg�]ֻ��ޯ��o\����ڡm�џ*�������BUg��n%�L+TAr����(=1�ni���&����s::{FG��v�I��Թk�                p���1u�j3K�׹���يRsb6��VR�Ub��<)���|1�dc�\�����gj�Ok����      �RH]
��ڡ�jI֧uQ�Ks+*M	�7�_wދM��G$�Ԙ�Q-���(��0�i��=Y�V��i�}fS���8{����I�|J��㚘;/                @�A;�5�Ru�<�DU�EJ	��5��엥���v�����Ҽ�͞���I�]��Хq;0u9�,      �R��P����W��+\�������в>����������2�fW�-�J���߻Tvb�:sk����5z��/�����I͇                ���d�f���Ը?�e&�)^�:�MY�vS���]]������>f�c����U     ��8ۗ�C����	1��7�a�hAײ~�y/(X����:u�5�#�J����3a:�74�͘_^���I�>�=����S
9/                ��1�N;r�m�{gN��Ӌ�p3&L�-��n�rhYG�L���#�s��_:��e��     <����;�CU�>��Z��g;�j-��P����"m�kҖ�Zu�T+1� �]r0��?���/ץ�Y{B}��1�������                ��JS�%��n]y�JKH����e����e/��Q/�k�������=+      ܐ�l�֌^����N	�2�b��^�(Isn}���6B�$�wmhЋ6�h[^��3���NJ�mv{�B�9���G��s��P               ��K{N�n/hUW^��R��1�Q�����W���)�]8��Oi�ҸB�      �J-iP��)}A@c|@-J�_:�6+%�-�Nw���JO$Q=����r��_�r�ݩ}��~�:%                �UE���SwmV~r��iv{���t��%}����{vPC3�
��     q-W!��v�u��_�검(������{���{¹��8ՒU����e���W�|O�L/�}�/�۳�1�>�O'��mGڔ>˾��hը�3��W�7��D�pk�2/i�jD~t^:F;���,�\(�@݀�R��W�g�Uz�T��sy�tx�a�U�R�:v(�nn)aI���i1qQ~U{�V���'�Nh�pB~�>����mb�ح�'��麧���o5iV�,E�+q���.�\�_���~�^���i�5\;,?�4�I)���R@�ҕ�+��bUNV
�v>�����W�ˉ�tp���[.k�~�'�˯�OW��\�pkE:QxB~�:���C�
���-$.h_�>���cMʾ�-�ڑ�G4���59Wr�x��sO+`�CuC�3�<�v-M��@ ���aͤ�ȯ��;��	֗+1�=�ъQ�Up9��C�J\��r�[����K�omC��
��+n�t�i/9. L8��m���S��w�O��K{�v�ڴ���0�1      ��J��zX��S�w�W�~M�Z��QH�SՐ������[�*g�M��ṡ1/��7N�ѷ���ܒ~�.�G6+�r��2��k_�>_6�L�}��"�ʘ�P�T=����Ƅ�t��V�<E�+�3ԣ=-{4�:+�)�,W�	|W*c"CII��J^LV�@�����������ݾl�3��&D
+�4ޤĥD_[�c�m��l!6n��mܮ��>_6�m:�ɆObe���`�/��6\�`����w%̾!�@��l~R~c֗]]J�F@�Jmڦ�M{5��f���e�8�}���sO���ߘ�s�)e� ���>�C��i.��|u��Tq�BX�5��~*6�ۻ����L��J�6p�v���b�A��:�?M@�J�i���&��T�s9G�#�vm�[{v}���/?��R�l��2[l��b��W�`BbL`5�˕1����d;��o��r����U��VK�/kLi��jae�P3(f�̿A�p���L�DA�^[����
Srn�Ƙa��8�����..�7�     �&jҿ�!���c��A1�f��2�8�LT�&���K�sj�DxWC�F5�߭wռJ�9;������e�s�=�t)�
�T�a�X�f��AM������B*�N�L�-��S3�Tkc�㻆���e�f����G!�ڔ�-����/�4gۨ�D��j�`?6�c��sŢ�zu�N����Ѳ���m;�M��:�a��zzl����b!]=���v�M�h�`R~q#���}%�o����/!]�ud��5�ӅL�4�An��)<_��P�j���g�̱P�b|^�\+��0����~ͦ����ҵ��������g���mUB�sO�a�{�;�˶�ZL�OX!�k���6�cɓ'����M֕�����>�)_���2�24k5lm��M�����F5�7�oX������� S�`֗&H+g������i�����ɿ�T�*'*��3�ъ����h娀H0��͹������f%X�{�h��կ�;�^�����3O�熵��5o     �HV@�j�^�DݯOjZ@�_��C�OK�������EzmI��,�Tf"��~���j/��md愾1ٯ�ݯ�K�B����|cm�֙�3�:�9��i�3�~��G!����-�[|3��Ę���	o,9WbS~h�c����h�k��l����Z���!1kUu��>_.�����+96�4`�RR�;Ыݭ�h�#�t��:��X�Ԙ(�~X�	!m9�"��9Oc&���x�������|#�����`�{�D�jN�E�D\�O3_�b�z	�Y+�.7A�{Z��b�{��fO��\�5�c�mÄ���ٷ��e�n�'z�Z2!���p���Ƌ��u����ٷ��hw�nϯ/m��VN��6j-n©�T���B�>~�C�����eo�^ͤ{����x���B�V&��<_�T����,��x�^S�Mũ�����l��d��s�O������S      V�Z�n=�7�	
���
����^��(���ڲ�tO����k��𿦬r�=P���ٽ�ʉ��5ưvR��)�n=ܪ��M�{���B��0��z�zl��WQH7&�7x���B���C3Ӝ��6�z���L�Ϳ�/��9�������^n�˙��惄Ĭ�	��>�]��vy:,�L͘%�t���5�f��'�U�ѻ�X��>���w�W��vk9��	�����9n�4�I�u����n3_��jUOT��f���T{^���	.mX�ޖ��I�n�	�+:Wĵ�u�C3!�ᑸ������ާ��9yն�mʺ�%�O͉��:VrL^Eix�ϥ{~}ij����c�����H���/©:U��	BH����:�/[���4Ay&��a�lmÁ�׃�3�[�@ix�N��ǔ	֣6�Dw���ś�`?JR���Uw��ʗ���ЗO|_��O
      N4*�j�ީ��agX?���q<�&�2��/-��[�nWuz���S���^������X3
�¯�h�-�8Y��#Ӝ�+�j����f�M棐*�Lv��N�h*�{�|R�������^��τ)���������6���f���q��6`���Ի�z��|��&�B~u'���x�qy��3�x�Q��3���f>BH��<߶��i�vؓ�|'T6Y&��������m��Ya��:}���mګ��/o����/7�B^&x�{����5�콠bBz��p0ǐ�'��}�p�ay!��e֗��oW_G���
*6!���e�B�!]�S�����1�����Bxd�f{v!��e��7�l���A8���W�B����Z`��
��pGA��g�����Ӯ�
�B     �Lg���g���)o]��k���AuiI_sn�ȇL0ȫ���-�/VAr� ���X+
�"��X���AO5�I�f�3�˄��6t�v���L3�-���#�i��P�mИ��NX�T�a��<�4��,<�̷et�m�Bx�f>�}��;�|E��z�U/s?0E�{��xf�;!��a���N�)i9I�7z���|�\�'��2k����e�.�4�Bf��z��6@M�{��τG�)��i���Ҟ�=򊌹gBH	�	+;�}d��5x������b3!��a���D�ͦz#,Ƭ/���~-]�ت<]i���+!������F������m��mv�Wӱ&{]�D�	y�9�d�?!��8ǜ���a}f�a��&�j*�;���FF��u�v��Ƨ�
CP�Bڲ*��z��^���N��7'��|�k     �52��ߧ5�Cz��w��Z���~P�QP_rne�g��m8�ݥە��,��<{2�Е	}�ط�����#:(��</5�1�9�R��ئ�����n
�lHӶ"¬�ڏ�kxiX��r;Ә�?M!U����4��\�Q�H'�:�f���.e�f
�Qx�P���h�+>_��#Ls��`'���k6���|��F^�D��f�2�7�BYII�>�݆������IMG���ɂ�r;,W8U��2B2�2�����>�7�e]ɲ�BH#���v�뉩�7�@��˹Bd�f��7멆��v�6��a����mh�L���LH�Y�ͧ	�Q1Ya�9�T������2�������|��,y)�^kM\�w�[,՝��ǒ^��8ި�g	!��}p����\_�@id���mcm�֙�3r;BH#+o&�s�p]I�D��x��V��'���aT�Q���߭�W�T_8�]���~-��     �c�Ւ~��.}R����W�w����g�ƴ����G��ߡ�D&2c��3J���{u`愾p�;�!�1xS��3H!U4�f>-K����4��H]HU��^WO棐*JBR˱��7Q���﶐j�B�H�B3�)�3����,S����&�ۧ9��1��W3����d>S��0���!����!wO~'�4:�c��t�4Z5*��;^��3Bd���7�B=�l�x�{��i�ax6D�9���f��+96���9��Cm��T�{�b!���K��o�#�4:�mޢ�M{5��ΰBH��t����ʭ!��l�|�;ח�6D�9��A8-G[T4U��2�L`���d�fhہm��;"��Z���s|��m �4:� ��o���@�^Zԡ{+^���<+U���_����G���|RK!ww      �A�����ޠG��"������>����HjB��.ݮ{�oWf"Ӳ�v�Y���z��.����KO]toA��Ls����<S4Q9Yi��G+���g����SH%���4��js��w��oCb(�����&%��4^�f>
�����|Ls�.sh��5��f>;�y�[i�X�F��'�-W�8Ӝ�ń������{5��f>�9G�Ʃ�v�|��ܦ�x��ϔ��l3__{����&��v��V%�����5�X�X�1�!����f���|�l'$&J�y��#�^�d��܆��rs3_��2B��0����lվ�}��鮠bs�<�%/$�a���C����B]&x�\��o��l����Mm�	�'�4z� s�>V6&�!�4�� T��A8��FYHj:�d�%O���B]YW�욾�ٽ�p��������W�,5_�Z���}�w�m�/�O|��     �g����a��>��Xum�T�f���=�`�޸q��)�C�I�¥5�R���s�{qL~������<
�bg�ٍ�He�jDn�r�E������$�����ݮ��G!U���Qh9��%��]��y�B�h��|�=v���f>3͹�H�]���m�Mõ�:�wFn`B*z�z�z-U�.�̷ux��lqOXLթ*�L��e��l�SOi:kZn�4��)�*Qp1���!�E��fO���6��׽�[����MqG3!��a�!�OV+a1A���NHLl���������*�($�k�!s��nCH��6Gi������ذA�#���~�.�#,���)�P���N=���������e�̰�=-{4���e�\�m�7�=昽�t�]_�V�g���0nn��3����m���c�|�x�{�B����@�v7�a1�'��6����*O+.ũ�60�'7ަύKߛ     �e*����O����*k>�]��Ћ���􋵯Ui*�9[r봹�V�?7������3D���m�F�X*�*��kc�B��2�1{�z��uO�'�QH[�ز�d����t�,��|���ʘ��*VL��[��L�w�f!6̾��p��4��f>;�y�G��Ls����l�c��V}�Z��Bl��ͣ��O~ϊm3!��Wt�H	c	�_�?�?��+:Wd��}��o��|��Ɩ9������o���o��2�E9�s��pS3_��"�ib��X����4^�f>c� !���7�/[b��W5Q��S��Ɗ9n0׉�5�;ӟń�vt��g����<N�ds샊��4��!��bY�u"s_�I����bkL)!11�q�A8ձ�c�5�^�b�M�pL�KǡBHc��D��7+9ӟÆ�:ǐi�!�����m�6�j��A8����R���ujϮ)��������	���o8o�3|      LL��!U�q}D�*����#�ӂ������I�j^����`S��Գ�Q_>�}}���4r��D���|��7(�P���v���g $��KAmܦ����5�QH�f2��=������3��=l3��v[P�f��g6��x�{MG�����'b���4����6�
�e�-mXL'�՟�W�$Ӝc�6�n�`���rb��g{Ms)�:��1߆=��T�~��ȟΧ�/����G�{l<�L3_U��LxQ��L!�l3�3a��j�+>_l�{5�kZ�xIl+L��i�KYHb+}.]���}c��gHM)bˬ/���4\;�3ygb�3B��W��ux��l�]X!��Xh���mګ��ج/��di��V֗.Pz�T	K	����`�!e]�b��ў�=�K����`CH�Bk���d��7�j!��r-�FP1a1��!9K�U�L�)ު`�냈��r=���֙}��#���     �+}X;�׏9o��~P��U���sk�<.+1M�U�Lo(���9b"%�t�N�6��c�Կ�yZ�PH��9�O��u�v��Ƨ������.�N~�o�ו�+Q��R��)�2a1fj�Het��(�r���g���wk>1��|&A�=����E����i΄ĸ�	�1Ŗ}m}Q/�4�Q&D
�`���i�nXgr����4g�ɝɍ��wBH�%��|���O�T�m����7vQL��	!�;��&����/��|&��a��}�K��C��:�Ƌv3���߭�EBb�sl���:���nPqÉ�M�	�`��GZ�����~oBH�'{6[]�]�Ӷ'�߻�`��/B�f��	j�׸O2/D�{S��>E�<�@}��B�.f}i���[�5��A8����9��<]i��c���cC�{�<�,�C�|�z�_#�� DNb Aw����/Wz"�u}�9�΢N�8�E_9���     ?��v([Y���ܸ%o�<�
�M疧�ۛPs�˕�HC.b� 9[7�Y�*ڢ�>�w�=+��	��߅�f���G!�;�b�m�io�^ͤG���B*�*=[j�T���c��{�f���6�1�ٽl3�r�o�N3�i3M!fwI�O��^&H*Za1&X�p��F���|�[�P����i�˘Ͱǭ���b&�wu���/j��4m�^���F3_�>]ȊN3_�t�����)<_���v�E��τ��}Qڵ4�]̔�h7�B�^&��K��E��/y)ٮaY_��	�����f���z��%$�uBR��&{,y��dT�%!��9���!g�м��E�!�D�ۘkU�F6i_���̉��2&_��	�q!���|p��jx**�Ϭ/���~�R�yvΞ�=�M����?��H�ܧb�A8U���l�vw1�3�bW�.�b|d��&���u*M�k�	�v(��;�G����     �#�ь��S?�l�d�My�
��~&$�NV�^�4�Q�Y�fSN��p�/�'�M����yN�2SP�4gw3�|�Ѳ��?���4�d\���6���d>
�ܯd��T�F���i���f���u�8���*&��ϲt�<�a1f��9n0žp�ԅԨM�k;�f��9lp)��w�IZ�&
#�4g�3���n���E����@�2�B�V����&�|3!��Wp�@���z���~��t�Af�0�)��|U��T3Q#��9'h�bl3_ed��L����NH�{��Q�@�#�O����2���Y_�Xñ{>r�x<�߇R�K��n}���"T�et�rfrw2�&�g�nPS�S�^�7��P;�/],�RnT�����64�d����ro�^ͤEvN��r[� �*�*��k#�}X_�_�bҍ��ɑ]_"�r�2����΢Nn�1m�>�v��75h��N/\     �Oܫ%�ݧ��/��WJT����s˳#�	zsًt�˔�����W�)�C/.h���[�>"x�)�"$���dEt2�-�`��ܘ�����RyG��u�uh���|}�9{G4���~���n渮r��[�V�F�{�i�[��*!DH��Ec2���<�4g/hoRR(I�E�i�c��w��x���B�H5�uw��N��]_�f��AM�E��τ�6�7�7��f>s|j֗�Lsv�h4�U��V��j��Jϖ��U"��S�Sm�!��gB��8���]k�k9ܢ��E
XS�]͉�o8Vr,"_�R�0��IEj}�5ܥ�YBH�Μ�nk�p��䝉��0��G[��� B:Э�BH���ު���t�tD�G�D�jNB�f�@{�=b�p���k���#�n�w�;ԫ=�{4�٠bD�mzo����.���}uKn�����7&�
�     ��(K�ک�9[d'
ó�w��C*ג�)�ĴfW��oTez� �(K��'�ΞD�ӣ����k�7�B�#Ry����s �a1���43��;�d���L棐�{�/�G���i[�c��)������|�Y�SLs���g7�f����N~ϸ�4g���d>Bb���x���o�c�����ys��B:ح�9BH��<nۏ�k�y	w3!��c��Lד-a^_.%�I�IKI�7���-�[��i�f2»��?^��3��zI�T�		w3_�|�%2�3�	K	�ZB[؛�:v(�R>�<�C�Я��.?֯�3���	��ԅT��jw��wu����oh=ܪ��M�O��k�/V�f�;� ��k�km!��c���s����©>U��j�;� ���N=��tX�.!��\
j��6���Gl¯85W﫿[�r9���LL��ۗvء�'��	     �ެ��s���:[d���Ӽ�������?9�<�՜���wU�J�/��d&����K�y�o��V}
�F!�w���ۆn�S;���G!�wݘ�W7�3��i�3ET��
�c���C!�w���p7�iQ�9�9{Q�T�m����c��w�c���iߣ�Ĺ�|�m�۔5�%xˍf��.O3Ӝ����6�/�wi1��f>c֗��R�	)��|��zW�l�=n0���`BHͤwBb��N~��f���Fj	�1�|c�_�?,_/c.î)��s��k�K{Z����φ�^"��k���r�Ҟs���4!��:��� s��I�j���B�C�]#�ԋ��6�cɓ'�����c�x�2AO�C��ݾ[�a�O5!���C.��\W�<ة��M�gNÉ�Mzv�`\˛�km�]_1���r�K�����~Ep/s�����ʗ+5�CxӦ����_��:�/��S?T�\     ��ӌ�[����+�P�s���V�<�1�Lnz����x]aJ�>�v���������4��i���g6��x��])�Rl�-�ZGXӜ���d���7�QH�}&,�6i��Y��1��=�=4�xX8�����}�
�>�n�o�#�r�:G:)��0d���[�5���f>S��y5S�&��w��珕���kB�}II�>�݆�����4��&�����L3_�b�N�X��!���LP��i޽���6�t���������r�EESE�/=,�b~X����d����z�9o�=�m�3i�*�2�E939�w� �x�Y��!������;�k��^'`�1�X�Rok8֠�bP�K���딟-W�x��]���~g}ٶ�چgBH�ynxTHj;�f�L�o}ij�L����v֗-�[_�@�m��2�3�ý�{5��A8���L�h|���x�	:zO�k՛ߤGG��s�.	     ��ީ�4���~�፫��U��Oέ-�Ӕ�ƍ����W)1@�4��΢N5dn�'G�����B��(�,W�	
�� u!U��{mA�Z�����#��O棐�?2�2�=ح���55�1��?LsƦ����n�.�-,�i��Qp�@���z���5�}s?0�A��x߳���:��Ls��R��t��*&+lc�Z�����&,�6���|���lH��n�,�u'���Z��!��}p�������g�mH�2�?</�|�:�?M��f�u���\���̈́��@`9�-�[��i�f2����5ܥ�YBH��t�Ԯk���	!�s�����iߣ�Ĺ��}�~�3أ��d���N�)i9I�7^�߯:U�����L��m�iW�.-W_�@��s��G�5�4�ɂ�5}s�P|����dϮo�K���pl�SOi:kZp����w+;�k���9���-������3�_      ����C��>*���yPi
��έnyLQJ�>��S�ȩ�W���������_���B��1U}�Z�'��0a/�agW��&�SH�Of2��������QH�?&�e-�|�L��shӚ��LQ]��\�?�f����W0]���v�?L�	�Y�d>c� ����(9[b�/TX��c����f���1d{ߪ������3У�E��N�ʘ���6��B�YBb��<�Ǹ	�Z���Y�nڪ���b=�|6�t�R?1a1��r_kߪ�^�L������#��od��5�Ӆ����P���?
��}�]u��{���GB�f}i�!���k6e�A�f}i�\,2��O*&*�s�X�ت�^��jUOT�a��{���z!�>�Z���k�>�r�E��m��ɹ��ΑN�!}�/l�|}}���A8��`��U�J���W�_e&��ךߪ�3���c_�ե��      p���C����� �?(&����y{�<掂6���ne&�X�K$�ʗ�=�J����]�$�F�ZUNT
�c�%{��ڂ���[_�����jN���c%�V��R��m��^l��f>�m��)�k;ܦUV���u�K�W���G���B�7�����4�#-���v2���luRR	*9Wb��+k�c������4��Rs�IH�?����R�J]HU�@�v�����4�o&�ԗ���G����j��LXP��v��|��lҾ�}��s�f>B�/Ӯq�܏
.�s�SO7>���'�Կ�uHT��e�fSW���!1K����y�8]a�9�V����ԟ�W�d��?�nח�5�x��BH���X�*/Z� BH�k��p6\ڠ�C�/}��N7�n�`���rV7�ӘY�7�Ee�����E�jˮ�#��WC�V7�     �UzD��煸����z�y�3��@�~��.��x��x�9�V����_G���W7)
�W�^�g(��3���;ԫ=�{4���ŖR��)��>Y���.���w
��/u~e�|Ls�?�oXi3Ӝ�/�J�����7o�+�*V�f���d��������̱f�@����*���f>�9��J��̱�i'�ԿV��G���� Ӱ��m�Mח�����g�'�O���!�?s��w���A�E��z�U�/��wh��5����|�ܔY_�@{�W�L��}��ɛ~^�D�jNB�g��]_�m٫����<������_�nT`9��ꑛ~^�x��\�W�R��lW_{���^��!�5�kZ�x��~��g�8k$u����l�d�l�OvΡ6��L�!��\�"���UJ����R���G:ީ?=�O��S�.      �2�X�L�׷����
���n��CR����l~���j@��NJ�i�_y�;���u�\����ͶɗF�.�mp�N~��*~�#���J[P�B�|R���7�]�Z����i���f�|v��`�����qAρ�n���a1Ls�����`���w2_�R�-�M\t�i"�ϭ��N4�l�L�?���=�m���̗>�n������l3��|1R���|;��ɢ� i1I���B�'������BGHL|�;Qg�/��g�G2f	!����g���b����!���6�i�vXg�~��φ�:���yBH�A��lmv֗-Ͽ�$�4~����T�S�Κ��?7�Q&Ԛ��Pz��>�>`�©Bj‹Vս�[�m��;���a�!�N�)i)I�˞Ζ�-ʹ�#�_�����eˑ��̾��p��4�aB����d}��'����Ub A�}���������y     xP���>���q˝@;�Z���M95���{��DA,u_��T��Q�����8'D��8^t�H� �3��N~�Rs���_��q
���5�m�b��?��nT=���i���������ү�붡�l��s���NW��$Ӝ�JHv2�iИ��QXL�b����Wďj�k<ި�g��O̔�-�[��i�f2~�1�L)!1q�t��>��f>Bz��xb���z��}���nBH;uBG^�����d�b칧��Z���Ϝ�lo`�G�C3_������i7�Lď��l{�`�K?!��ǜ�6�����Bօ���!�\ě��jk�����v�M��	��'��6�i٣����B�*NW�cɱ������.e�f
���ܮ]m�q!�q($5i����B�b"ic��v�Ϩ:�X ��t�.�T��+�Ϟ     ��kI��u�>�3B\r_��U���$Ot(�`�7����5�VB���z74��7��>1�W::��L$ܘ�L�L�1Ŕ�l��潚I���*��f>3���z3�T��4unڮ��>��G!U���̷���_o��V�B�R���(�4a1f�����c��G�5�4�ɂI��i�9/1�9�f>ۤѶǾ�4��e'��l��̗u%˾��2>��f>BH�Y_�����M�%�4�=�����f����0R��W~�\���B|j:�d�%O���0=�=J\��%~��	*�a1ͻM�!�q̬#;v���TΔ2�f�뙄�ħ�����SO��m�4!���ww���'5�6Ci3�s��4�F*��1�(���O���c��q$�S�x��BI/¯'�Qjz�29�<WEZ�>��}��W�o�     �A�
��S/u�Y!R�*Ѳ����Dgszb�nx�^��" ϯ,5_Ot�[��k}ojPST�{)W�_����V�m�a R�73}�m�M��(��4��f��q��!�UNT*�T�b%-$	�+e>�[��=���Ls�k!�e�E�K��:Ue���2�2m!���*�. $&��f�M7]__��#$&Ιf>���<��̫�8U���߇�t���jN����f>s�(�P`�B������^;�b�B�o��}�|��6�"~��&�|&s��x����h�QU��f}�L=����x2�2!��,�Ж�-:Vv��%Tz��ֻ�pbBH�۳�pN����j��(����Bx�c�wT�\?]�;��3� ����������}�Y҆     �1ݺ��:o��{��P���E�'FK�'g����.�T n.-!E��t��"�_���o�AHS\Y}� \W8](�0�[����`��)U���f��)ְ�m�1����0�Z	�aח�4��:���Y�x��4�K\g���H\LT�$!����t���Sv��I��f��i@��;U���	�a=������(:_����Sv���
\?�<SAPL�$�������v�9����⥪I/�'G��k�     �ޮ�էO��B\qO�V�s^�DP�QlCb
S�v��)���e*N����[-��               `����Ѷ��-�R V�E�-�d�;���ԅ��     �Ճګ'�!n�#(�a�ݹ�W�-�^���6�'��꽲x�Y��_���9               X��i��U��/ �לU�'6�[�=�y�Ϟ     ��$*�/�C��#:!ą��<�MZ�g�뽶x�~��J`�6��걎_�o}^g�]               ��k˪�G[߮�tX���<=�����/h��     xH���e�W/�gtM���|DyZ�W���J��w׼Zo.{� �GUF�>��n}t�/t��)               X�;�:�`�O*1�  뗙����v��8�����}     �^%�q���۠�y�����A{���E� �6$g�ю��ǆ�J{/�	               ���Uڣ_�}��� �OR0Ql�)�&g�'�M      ��zH������k��١��o���d��4�U��
@d�&$����w|I�~��                ��{����W�R "�0=P��&e��g     xF@����1��b��ן�����h�G���Y����6}r�+��Ԡ                ���*_f7 �gB��b     ���*���z���%�������3��s+K.�����-o���Z���@�~�����ϓ{               �@ �j^�7m�M �ǄŤ'��ƾ���     �zݡJ}ع���/E?(fF�p^o�Ke&��m��%�B �+���Tz0E3�C               ���ؾ��n��x� D�]�=6,汃�OK�e     x�������EӾE7(惺C��k�2!1���N�g�
@l�i�}�M[�ۉ]               �U�y���&�Y�) ���g���~�ֺ     �\���>�-zD3��D/(�C�Ғ>��J������^Bb 0a1�T�:-,/���               ⍩��պ��\�,���ġ�V(DX     p�:-���/	����E����%�����Ԟ���K���{�ߠ����׳�               ēwU�R�/� �xU�]]��?�{     x�/�a}Y�ҷ߈NP��ڮ�;S�	�͖��3�F �%���7kni^?<?"                �l՝zK���>o,����9}��U     ��
鏴S��6'�B�bv*Y3�3�V�\ƄP|��ԓ�( �t=������T߅��w%%%(3=:�d�0���W����JVB0 ��8}�9�E$��$*=�u��?�ڵ%��-
�����v��ny9��y!��R����}��좮-,	���ٻ��������Y4�mɖ,۲%y���ر�A�
Jp����H�r�5���+p�
d����@[�VRL�=�eK^d���K�e�w�Q&�JB4�<#�z͜$h�F����|���S~n���7�9��1�ɖ���P�_�u��sv�gS]0���)b1��?��D5:��2�r���e�����HDQ�߲)/
(+��kO�Ȭ3��2��r������3��!g߀�
��1f*�/g��eTH���t�.�0q�)�Re|96>��Y��g��|V��)|�)fg���8��d��
)-h���1�'f`&U��m�����$�_&[^n�l��`Ɨã��5$U��/'����4מ���p˟�8S�c�`�w�<O�s3�A��     �\���)g�)aQH��ڣ�+�y�,�s�n��3��d� ���b�j�;�W���#�-BjZ�$[�R��I�c�jn�ؤ�dg���వ�͒���^��I�̟I��U�*�KS�⹖�Ój���̤;��5�v�o4�ɦ>�����I�u�
��2��<Nݽ�j�V��S�E�L��{�j����o銝���Zz5<&$���kr|B᰽�s�0�p�d��ڶq�fg�e�A���VS۠F'�$�{F�����e��}CCK��&��$�(���di��~{C�#Sja|����Q_��҂v�̐����9��$�XU�#�
[|���Sg'�K7���"~��o�J߹����44*$���+559��Ǘ�]#��6�!����u�ie�LMă�6���U�3���]k���������MLJ���N��e9Z�2W���F�"jn�8s���=k��?h���\ih�u�>�|�f2UU,QV��9N��^0�'��9�?Iv�Yk��7h�M�f��e�3�f|��.[�K��D ����hbnZ?�|R      V��ݤ�z^Hy�]��q�w�o��>��B�n�6H�@H�6�[7�K��}Bjڽ�BO<�`��(�����w{Y,
��li���h�nBU<��'��މ��Og��#��+�f�ߟ����XU�D��4uv�*�l��B$&�w��bb~�{wU��ǎ)la,��o�9w`e�[6o\�õ�233USk��~��a�Qz(����g땑n߂���!�=1��ې�H��O[�'�mTlξ�S��w8g��ܐ�VYi���6[�1:�#���=g�գO�+-h�ߟ����c�;���+;+]�-=
�:���Ęq/�K7��>���Z�y��3���`��kllL1�!]Q]Y���>��Y���/�s��n�ڳ�R�=y��XLG��"�ξAp�i�����+c1&���'?�W���5�kt����XLSۀb1���,V{w�ӣO�[�1����Aq��eKrT�����+�6�H����p��1��ǜ�eȾ������X�fi<��3`],&U�&�/S���j]E$H)׬�Tӣz��V      ʧ��
���ćL).����Ƿ�G�,sq���l� ���`��zӕ���]�RS<��I)f�-'&g��=��}���⥹2���׷Y3�*�i�%�2�߯��\�G?�P��14<��As�a�E��ķ6�b��)s�-"1�2v��c_,�DbF���o��fb15�Q���[���܉���W�`Ls�:�&+3�3v��.c��9==);W��a_,f22������r֞a�WT��MW�pm�U��ZM�7����r��u��bFF#�5Q{ޞ���e��M��<��p�&��o8wo�u��ށq����SHw�X�Q�q`��XL�N�-��˨=��E/==��<���7�s����TdBp�|,�Y�){��SSsj�싏/�\�vM^^��o�/��6���q���b��M��H�Kw-/ɋom���#1�Db�_��C�w�v�3&342�����X�9g��7hM,Ɯ7�l�V0S��eʪ�)�_T_!��?j ����[�/�-5��m     ��N�*]�l�,���bnҕ���΂J]��M��J���w듇����R�����'����[&���O$�#��r��2kb1�-}���H��XL�5���b"�Gl���/��q�����m���q���̖�e��m�"�ĘǜCz"�y��z+��#1Db<2�iPln���HL�K��X�捫���4��H�7l�ŘHLO���bS,&���Db��z�,�;kO�~��2Bޏ/M$fd�H�W�W���q;b1�����">���b�<�ʚX���LN���i�VY�1����^�=y��b�lZ��#�V�/���xj~|yB>''�%�b1�HL�����9�b�Ɨި^W����GbZz`|���cÁ� ���?M���n�p��     ��b��>���U������F���oe�ՙ�t��+���4sǄ[��Ч뾯h���8���ٵ��X��Č:���x͖XL��İ��S�X�Ï�P������I���X<����ϳX��>U��">��X�Y�_X�����?F$�6�b^��;琞2���-�Ŵu)2=I$�c�vTx�!c[b1&���S�-�����z�Y��5��9��s7e�b1&s����ǂ΁��3���c�=���N�������i�\����^_���K&���J=��	�=����=�����X̳�5�n�?5=���>�=y�� ˊXLs� ���]�/�+���=61���A�=y��b�9\cs����fLA$��X�o����X���$���1���fs��=���@X�6�[�lH]�i����?�M����      ,����9۫����PL�nu�W�"E����+����]�����tW�/���e,&��!c��XL���hW(��	U&Ý���O�}��c��}+��'c���K�[/b1�HLS��,L��y�1���1"1���b��il��X�܋��� �9m��~�'����a"1���4*6���)���H�=�c1�:\���b��V"1��:���2��DyiA|�E,&�����E|�0����x�����(�Kl�Z����$c�/�c|i��p�v��],��H�Uvl�.1���~"1��:��6��hD�����9��
z0��Db:{��
�+��[/b1f|�����&s������KKx�17�;��痩.��mxg��� R�ʌ%�?ߥ[[3Q�     K��!}\w�zVHI��E������@(�Y��' ���{�95��v>%��x,����[�?19�&RY�xYn|�v,���_Db�b&^�����X��Ȕ����ƋX̋�?��x������l��~,�H�����=�Ŵu�H����ڱFO>۠؜{��im'c����x,�H]���˦��bDbl�R,�Ғ����F�#�/
,�b,���9�s��">;�X��{���cǔ�b,�pB�Db�����܋Ř;��$c�b1�=#�$c�c1�S�M}���Us<þ�&/�bL�Խ�xs�����p��;k�����Ϗ���ɋXL||��+�K���y��H����Db��c�"^�b⑘&�琩��ʷh{~� ,�sW��uo���H      ��+��s�gk~9R��O����S�,a��Y%��\]q��'zT3�$��=�+]��LEf��5�">K��i�GbX�g��b1G]�x;2Qo������f,f>�K$�Rn�bz�ǉ�X��XL<����\�������^�g6(��ݝ;�G4==I$�R�vT�����Sk'�[�X̦+]�ŘHL�E|V���T��1���^"1���b�1���$=cF���H����9{���c�v!3�!c����b�#1�,�T<s�:=�L�2\��v��jbr�kO�r3�Ĵ�)�b�/�|,f�j����Us����_�ʌ/qƗA>G���Qg7sleb1�XLM-]��b[��sƗ6��b�V�7f|��q�H���g���?��X�U64��(�ې��Z�G�/�& ��뜿���N�s�c     ��O{�q]�/�B�Y�i&�p�Q�U�|�^��d� ,N�_Y�v]w�N�GF��eb1�>Y��N�7�e22���~&RY��b����Ov(-��I4�}��`�x,fO�~��q�Cɛ@c"1=}�Db,gb1f�eW<�����K�&Y���b��]�7�H�b�ށq����P�r&s�H�Ɠ��5���^��X-''����ك�I�Ř;�Oq�w�X��4H���bL$����7pi5�b1�Db����<�x��^H�1}t,��>"1�+_Y�&3��4����Ŝ�B,�Db�F�����b�E522��XL<��C$�r!�ޙ�X�|$f�kO�s#c"1Mm�Db,WX��J,��cXss�ng�Ǘǝ�D��&����ە��#ٱ��an��ⱘ�܆��b�Ĥ�����Z�����8����H�"�1�\�_}� ,^X}�N�upCT     `�/j�~�<X(�bv�IT_�d��P����}�_/ �[A([�Z�}�з4c�}*ۻk]�b1����*��ŷɊ�4��HLj��PU��;��$�bF�"��'�*֮Y�&#c&R�$�2�BA缡2i����q���I[7�&-c"1�&�"������B,�))�;L$f�k��b��
=�L�bI��D"DbR���l\�R�G��i"�2L,�3�%-36Qw� מR�����ͩ���ǗfyNc3��T��X�Y�g"1�/S���:\מ�X����7�@��RA"��3�ξa���}cDbR�|,�I�ӑ�33���p�)%$;��9���)!5�1s��WZ�DbR�K����HM$���!�I�܆��)"1)��b�)9������Y
���}��,qC��ܩ�in�
     ��R#�J&���p���t��K�X����f.�X�6�ԇ�\�;~.�6s���'Z���u�0�*ŘXL��؂�+�)��_,��1���ێ����-���9ŘX�Y��Г���'YėbL,f�����nx����XǾ!��X��#-
�vR���/wzO-&�bE��#�����S��];+t��y��oGO����([EK�KB�enn��)��b�o]������&D�4��Y�T��S��baǗ�3�~��e*1����R.���o�e|�bL,���vu��I1&���X�c��O0�L9;��VMm�s�_�}������bb1˖�k.	�˩�)�)Č/w�f��:�{�t�^H1&38<�'vn�ܜ9$�J�܆�ե��X��}���HL�1��������?0����e�3q�Omx�
C9���o�������D9�     ��V}Rw�sR�B�b|�קe�40^Y�K��SǛW�V�x��~^               �M���D�rW	��c}�J}d����ɟ
     �BK�u��o���0����6�y�,quť��)�S�ukߨ��5�w               ��닷����S��ۯmՃ=     `��>��Н������C1W( ���{�6�Ғ�pjJ������wj::#               �K�Å���p�~�tt�M��     �L�f�1g�OH	�>S�w9�e���\}��28��g.Շ�\��N�L               �W>�n�~�2�p�
B���+t���4�     �Ub����m��z뽺P�
8��[�9_��|�r���7���g����1               ^����j}N� �2{��]~�����      ,���nr��
�{u���z��Nx[�^mϯ >�O7V�EW=w�g�               �iS�*���l@�;W���:8�(      �\�[�}VÂ�^](Ƨe������U� ~[^Z�n�z�>U�]�b1               n�
��ɪ���� 	>��ξ���n���      ,��Y}��~A�ڟ��Q�:ϻ䱐/�H� �kG�:]�|�~��                7\��*� ~גP�>��2���     �27h���<�k���>.�o�Z��L ��|`�zz�:&               $��K6�K�
 ���0����     �"e�۝�����B1�T���y�*�To^�K ��	��t㺷蓇�Q,               �Y���Zs� ���f���P��f'     `�>�<�y�0�RZ(fVw~�~y(���c�.���� El�[���F��~N               @2|��b��
 ����l}h�E�҉     �E��f����W��^y(�z-�OW�co/;[k�� ^.���3C�ꏌ               XH[���ol /��g����C'     `��;B1�z塘4��y�C�E���
 ^��@XW��Ds�               Jȟ�ֽY>�O �r�}���]����MSs�     �BL�Z��+�z�����R=�s�n�|�B�W����K6iO�=�_'               `!\Y�Z��( �R%��{�y���~     X§���l��`�WV[�Y�)���%�wjs�*���ڊ7���M�E               �k�J���=�?�ه��=���]     ���a�?��f���PLT�O��f��� ^���\�s�9���               ��U�*�� �Tfrͺ7��Cw+�	     �˕�K��	Vy���[U�i�U���󔛖) x�./ݣ���S�T�               �?��K6iK�j���)�\gm��}G     `�>$B1�y���]�<�呕K���g B����\����G               �T��W_$ X(^s��8�HtF      �D��\�U�`������Ї+.�� `��-ڨ���깡�               ^�����8�/ X(K�����=�~�o     `��f�g�ׂ5^^(�fmUL����tzA� `�}d�%���횋E               ��l]Qz� `��s�9�U��F�     �9��%B1Vyy����!�|~}pՅ�dX��L����;����?�����y������RC,��䴢��ߘBi!M�L�c`h")��¼l
�cffN��Yg�����/�@ �����!yF���o��������:��#���1��}3�a����L)�cMO/��!;+C�SB��O�q"?7[ݑ	gl!�3����8�z�?�����ch(Iמ�s��N��:fg�455������
�4;7#����7��1�?�LLN;��3�iaǗ��i����e��e*�t�I_fgjrr\HC�S����������1I0S�9V�sɅ���tdJH���I�ې��~��dn.��g�נR,SZ0M3��/S���d�ƗY�ؕ�e*�L�*b�=-��5ם���3�dn�->��Be� -ݟ�����ϟ�g     X`�n�V}^�+��P�t�<ri��� $��,�~�sP�sD#���?�ёq-_��������;�Ť 3����v/�J��/��С#M�fBUJhm�?6��}�������c1_*0����:T�,9����t�kQtnV�߉�=��('k��%K�u�h��GG��HLsK���$���d�t����|)�p]����D̅����(Sj[59I,&��k�$i�ˌp��Z;�!J�m~|��N�¼��5kf��J���k��]�$m|y�ɯΞ^�~ѹ�j�v����!��7�8��9Ɨ)���O!���%g|Yw¯�!Bũ`*2����X���eXG�[_���c]��	ɗZ��]�4Kk�4>>&�oxxB]]�Z^������[:D,&5�i���|�%�:Xע��I�~]�#�D��6�L���-��\{:��K�&��S~�3��m&�"�Z�
Ē�o�_����`?sC��':U�,9琹�!9�B,�k�Jt~�6@���l����q��     ��bz��L(�<s�v:ϕ�@��;V�- H���,]�|�~�����Q8��6�^���|RK��������� /���0��V���E3�,�Yk��f"�
�I{���e�����Y"�����0�d�kce��7k�	UV3��P0������ח��Q��\"�������
3U��:N,�z&�����D �����:X۪	��n��"1��@�^��$W1竹��X���B��#���2y�fQ�vg|y��E���`/���PZZ�ƗkW/�-b1V3���um�O��2;3�-��Us��X��L$Ƨ9���_n�,Q퉨����L$���[�9�_����u��S�s&ɵ'��HLfدd}��w��e�bR���tv*3#-i�aƗ���L,�v���e~�f��mC�iRd���L$flt\�P�=U�*t�1�w���'wnCf8M[̵��&��2�������f$s|�\u'D,�r&s�DG�F5ɒ��ƪr���ܕ�ΗO�C�<fnԕ�Ӿ��	     ��t����W���~Uo\q���r �vE���Y�������?��HLª����Zkg�X�g���&��̤�-��������������6z��XivvNuGە�¾�,�P��X�Œ�IH�bj�I##�bl�F$&aI���J?٪h�X���Mn$&�L�޶q�ԶhrrB���Ф����N�"��������������d� L,f��U:X۬ib1V��N~$&��b朝BOo�`7"1	�Y��X��c-,�TCs��I��$������;���0��l�F$&!��,��m�b,��HLB"s�H��&���ȍHL���gdM�H�5�I�{!��dƗ-�D��`����Gb֔ŷ�b��F$&���nXM,�bɎ�$��qƗC��}�p��I�!Sw�_z�*�T�
� ɶ��Z�s�tt�M      ���u���g���4>��6y �ҳ n�����������L$�`ؕHLByY�b>���X�M�'R%�N���XL�۴u��I�Z��9����@�����ֹ�I0̈́�#�}�:��Db��l�.U�Qid�X�M&&���ܣ�l��L,f.Z��ƶ�y�q�ΝHL���}���s�&�&{O��gЕHLB��<g�Us[�k�'�qnFb���F,�J&3>6�PZ��%T�Yjވ��#Fj���ms�ړ��l�Z�/�Y�g�x$&��HLB|1_�r՞0a;b16�GbN��I(*�T��2�'c��㝮DbL,f�ƕ:Xצ��1��#��EbJK��[b1�1A����!��e��rb1r3�`b1ј���I|nÑvW"1	��W�o�3;����Gbf�3�a>S��'b�g|i�9zܝHL��Ŭ_�RG�[��x�=���! ����u��#�     ���<�X�_Es�v9ϫ�7/ߥ�P� �-o-ۣ�|R��,�s����U��HL{'�x�I����m����=���L)to�eB����>�o�X����$�p��Zb1�0���@���V�X�zb161����nW#1	�K�䋕�DSv,�v$&��b�m*ס�V�=9!x�Db��ݍ�$�;�Ks�hn�`B��#1�FbL,f�Fg�Pע�ib16�"�PU�,>���'c/"1	9١����E��ؠ��O>g���?��XY��Gc��b$&۽HL����X�U⑘t����&X�mC�s٦1b1V0����ee�?�4�����/��d�#1	�X̆r�kU$�����Gb<_�]U��[Gw��#1\{��4��rgL��[��I0���+���OC������$�ehC%sܶ)�\;��	 ܲ�`���V�p�      <�v�q��`b�����4>�I�������ى������\djrnz"���b�O�f���~�?�y�gu��遴��@zFV0������/"���a]^�W�6�JH>/#1	��
�F���ݷ��e$&a>�J�ꚸ���^��ܟd��~]���4����x�,�=��I$&!�X�5���$���idtT������eKMԶ�X���&�����~�U�S�b�d"1].���w��ȗ��ss{'���q�w��αu�ty�I�^�,~.��G,�K�Q!����S�s��i=��H���D ���ҧ��W��!FꥩȬ�뻔��ݾ��b|&�Ъh4*x���.O"1	&c�=�uƗ�H=�e$&aEIn|&U���n�$B�
�u}��5kfzZ�Noߨ�UzȻk���ķ�b��e$&��b6U�T�_�1��RKۀ3���V�s꺡�Du'D,�c^Fb�܆��V�h}�K��g�����h$6<3931;��NOL�͌�Ţ��ٹ�I_@�����>(H����23��������?��{]Y�Z}��     xl�n�V}QO��O�/��l���f
����:'&��G�Gf�k�g�L�f�O�<�����{5���_�`{8<=ݟ��y��(HϮ(N�/*
�R�9Žy�n�K�������HL�"�b>utw�!�`�nݰ�X���:�<��$T�-����o�X�L$�p������f�%�/�7�*�y��޼���R�m��ww����{<��$�XL�W��Fb1^1���L��f��M�b�44<�y$&��� �%�x$�_�[0�|1s�I����&3�q$&��bY||��O,��HLm��K�ټ�\5�Z�q/מ�����i$&!>�\_��GE,�#��s����4�PT��j�$�!��H�y~pƗ�7��`m�&&����cS���/��ZiIn|K,�;&��a�4!�_n߰�X��z��448�]x��bb򩳛�x��HLBvV��8��������hm��̴g���D,��DT�CÂ�l��$�gh��r�ou��mH��yښ�F8�E�s����tod�{02~lln���\�@dr��o�?N���}�W/\�!ߙ���ف�k
ҳ�������>o�=����}Ё�     x�o������-w���e�����L��3<3m����yzxv���YS?��}����Z����gs�w��{?������,
�_���aUVqN��꧔�>hř���WBr�#1�vDb*V�狩��	Un�_��aE$&�,.ݲ~u��[��L�t�|$fҊHL���Dc�� �7��Ix��[��b\6����l�sl�XF,�&��ح�l�g$/ɖ/V��Mmο�`�M�G;��a�x"�ٸR��h�9��{�#1�VDbL,&�3w���cS$&!�ٸ�9o �6�"1	�k�ŷ�b�eS$&�D�T��Y�G,�U&��z�IH�bj�I##�b�d"1�OtX�I0��*��q��#㦣'����$�}�_�q��Ĵ��[�I0�������!���a��=�!��C�-��D��#1��������UE�B�:{z���I0��MU�t�x3���H�L$�`Ў9��Tvc�
՞����I��b*˜�N��$zW��©'27�����������O�L��7ox0)w'����7:������W�qᲜhڕy��K���m]�Y�$�g�w�}ЁB1     �s&��SxU�_��|\vQ�e3������y�g�y������w��M}o����~r}���u6���|�u��|Y+�(|ce���L;>�ER�a���A�C��#��l��$�)/�!����~��D*��%�I���[&#���m탚�O��g����ֺb՝�jl|PH��٨jN�� 7,��ehCe��~0�&T���HLB"SSצ�a���HL²�ي�LG�}�q�x��2��ٵk�O�f��^g�,�s�|$f��HLª����剦.�5G:���$��Amް�9o`|�x$ft\��]�K��b��q�OH���>R�a�"��YoƗǛ���M-vEb�9��R���GY���HL��,�7,)�t��C����ĄdM$&!�9P�C*v��XĺHLBYI^||y��]p�m����x�t�֚sHƗn�������s֮^ߞl�F8n0�K�"1	�s��U�:���'7��h&2mM$&!��;���s�`"1�'����$d�z]���d|���+�5o�pj�͜����xd�{o�?����ݫ�7'�_x�w������%iyo��.�Rηo`�g�AU9�:>ʵ     �3u���Y1��C��l_��㪀ϯ���-,n&�8����ɑ���c�?&��}��Y67��{�9/�5������[�WV�Ȱk� LN0C��w<!,�����M��]�%~[Z0��4'���`M�rsB����rs���/&$��ЄN6�*��������|f�������g�8�{�a�,�L���a�ͤ5{w�q"G�N3!���������
��58l���p���霰SBCs���œ����媵üW�x�L�ȬԴ8�K�>�B!�fag���͇ FF�=N��嫥ݜ�F����X}�,���p8]��Y<b��u�x깦x\��kO����Y;���oD�4�94[+7;K~�����2�}Ҍ/}�xߐ���<��3�ZچT�4��KO�9�3�l7�W1�L��9=�7����o�^8=�y���X�
��V�/���%�_&��Ĵ׵[�miii�mp�3����f��27O�`|�l�jl��&�-+;��.y����/�G����a>���{�ŭozd��X����_���������>�sw�Ͼ�Ї�zѻJ��W��\ʵ�x����=����     �4�����G�g~�E�+dn��z��%U.�ɹH��H�Ѷ��O����t����O���M��(ܷ6{�{�rJm��^���أ�v>��x��Є�x�IJ�w��[���3 Ƴ�:M���0;;����.H�w�d�����϶	0�e�u�����|M� ��}$� ������������.���^P{�W�108�Ǚۀ<�%�h��? ��/OMKB��y�X|���N�v���vgo�/��w_J��q�/�����y��V/��pYF�u��Vo�ӄ�圢M�v�W�bn     �O�P��~(�\g:υr�	3`q���n��eb������Es{�*�7����KW�|~[ޚ!?�Ţ8��=E�p�              �����=
���1:3=8��h���5w���Z$���?�_���������7.�(�}{~�ٹ�L��(�}~]�b����     x��\�<���>���_���U��)�Ɖ����/��}�\p�"�͏=�sg�ss1}E�;v�=;3�	)��ҽ�b               NQY��..�!,��#�����eb��t��瞏>X�lλ��gf~�5k�X�宨���ŧ�{-����      <R��k���Z���B_Lg��s�m�{���>�7up����7u��Q�B^��~����e�ܻ�ȯ��`Lj[�S�Xi               N-���Tf0]Hm�3��GN��k��]�޸H���8���7}0ky�K��}���<�1),#��KKN�?�=,      ��d!�b<�_/��s�ۨ�p�X.Ю�j!u�O��>=x����n�ʾ�D���T���e�������p}E���_������-+�$              p�1�/[��z,���t��ct����T���o��Ʉ���{�t�-˳��㮢���tn���.[�K?lT��)uo_     `�X<s������V�9�����k��(27�'��G�������{��G�ͦ�v�۶��FUvi��rvU� ����1              �԰#�����'������Ǉ;����/z!�s�{�t��ʼ�tZ~E���Z�T�$���*���1     x�,�3�5��n� �_�FH=�c���|��>������k������Go{��^��c9i~!e}�~�v����               pj��d��zz"C3O���ۯ���?腀N�շ_z��U_^�^�.���Kv�     ^Z��\_V�����og���*�VQ(GH�sS�G�j��׵����wgTxY�r�On���77���ּ5+��a.�������               ���e��*!uDcQ=6p�ѮK�q����q������?�e���̢�{̍���(�����     �'��<�Pp����u���x��:ǻF�8�>��o�^�{>�`��)��mo���6ߐ��	�+iK�jn               ��OS�RC����#�u7�q�Ͼ*�b/�u�^u�%�?3Ý���4�z&�sA�k�	     �#{D(��9�q�r���z��y�Q�N��\,������Co�o��«�kr���"��3�O�d��ֻ�d�              �E�����ӄ���PCS�T�Y߹�?څW�Ϋ�;"��.�5���]T�C?h}X1�     �{O��P�O��y}���������LF�_s��W��s������gzYg����,ٸ[���%�s2C���              ��-o�����o�:p����}�
�;Wǃ;kn���}���[�<��Z.ж�5:0�       l�>�Ǭ����i�[/�s�.,��n�����'�����k|ZXp��o���9󆯿���-����?M�S���mӏ;�               ���wv������5w^��I����˕c�E9w���B���b��      �֐*�m�����i�b���r-K��U3���\�a�����'$՗?�㫦�~�­w凲��n�s�l&              �H��Ӵ��Z�W�d���CG^��kŤ�$3!��;��ڕ����̥���,\�p ���i     �ί�"����i�[/|��͂��8v�׭�;���?+��Ϋ񭙯�՟U���႐`�9+�,=_=�!              `q�]T.�N�F��5m���_�
����_=��rl�x�����K���Uz��      \������^
�ܬ,�T�Ƌ����E��b1��?���~����}��MU��TZ�U�-X�����%����G              ���%��V��[���߳��	�U߼���+�]Q6����5���9�+s��̈́b     �7b�*��PLT[�ߍݚ�ZE��.&�`ϡ��U?�\��w���1x�6F;�6�$W��9�b               ��@H�T
�y~��阚6ܻo�������7�}Wl���fG��*�*�V)3���و      \F(�/�b�ڢ�;/zv�&�.&��|�y��{���u�U�b���W�	֨�.UI�@]S�              �Ⱛ�Z!�`�g����e��}�gO�X̦}�6<;^���j�`��/�]��u�!     ��\7(__֐���B1Qm�/�/���u�B1�y���?���w���g���?�k�W�V��|:g�f�S��              ��p��-�]�l$c�}��E���+�j��ѝ���k��d3�     �����l\��^��n�[���,�����g?|��u����C���&�4t�,sIX��9K	�               ,��t�(�ya�������Db�s���˺�-��i'��^!X��òa��M	     �U1U�P��^
���	��)� ����}����Q�ַ?�'}_
�y���O�r����e-ײ�<�D�              �Զ3�R!�tmqr�s��`��{o�O��R��o����:�Tf�(<��jg�:����      \�j�U�}5{�/h.����-ݵ�3g
ֻ�����%%;�%+�	�ۑ�N��~V               Hm�0��=�����N����C���v�X�ߥ��	f.	�ϙ�:�b     �����ܨB�97�/V.Ҋ�B�{��=OO�o�o��i!%|�_�8����Pr���}~�[�V�              Hq>�O;
�	������?rѽ7�TH	�~�����K�w>������YXߧ�b1     ��G(�m��;��wRZ��������K���>!��v�����od�{��-
�zM~����fcs              @j��*Qa(G�V����{��|��_�ZH)w_�����C������pCTo�e��i'�:     �"B1.��u'SH(�k����j�����������.9jjޚ��L�LF ]rW�f�I               HM�s3T+<�w���]���R�m���y�Ⱥ蜥�_+xjg~%�     ඕڧ��\1��i�|�}��?M��V�z���on���������}�m�Y�Qذ$�<c>$              ��v����Ѷ���MJ�	�뱎���ۺ�s�
Ϝ^X��q_a     ઠ�T�l�W$"��~��y��x�y�g��}�R!��s����ۃ׿��;�>����ේ               ROf0]�s���LFk�.�{�7�BJۿo���;��_�Y�lN03ɷ2��!g���a��N	     �5i�fI����P�OE�~���LE#�g����}L�����΢o�����g	�X�Y��P���G              ��򚼵
��w�?�������¢`~��wf|�ŧ�"x"��k{~��     �k��,�K�/l�$������H_�������@�-K�3�f���|ڔ�J�               R���Ղw�l���?�UXT�z�O�����wlϯX-xbs�*B1     �mIo��%��b�Vg�h�}�s�Jaѹ�}��B__]�Qt���ܷ)��P              @
ڐ�R����D��H��E�v����쒺�`&��=�1�\      ���qS"S��Y�]� O�Dg�l��w�߷VX��qݿ{�7o�]�~��:.�              ��t�*�Ko<�[{�=}�VX��s݃ǋ���͋���a�uk���o�<57-      �	���ٻ8��:���S����s�ؓ�a$��we�^W���껫��k���꾬CXT\��ADǰ
�����9����sj�0��z����OS�a�j��~�<O=�wfC1�*��0!�B����_�w��	J����%��3=��J�L[j�
�Ob,�              �5��1���L��v������{݊��}`yh^��Q���WW-��&�     �!�xd�x��*�O���PL!L$#����傒��u?�o�;�����Wub}��8q\               P�U�ǽL�k�D�Mw���
J����/���!��Y��[	�      �R/p�G��?�U7{AoM�B��?���^��^AYx~`��5U×/6VuJ�bB1               Ed]�PL!<?q���7=�5AY���ǿ���[��,_.pԺ�E  ��ʷJj<5bx�>��HjDF
 ��4㱾C*�`i�YB��Y�����A��Ӷ'����?,6�?G��^,�-               (��P�r1Tǥ�i9�BPV�c��1��k��#pκ���2\�5�  ��㱎��W�>Yg�#kHee�TUUI1x~�yB1 P����>�dů�	ְ�^/L��������?z뺇Z?�,�8����4               z[l�JO��Y�O{遛v?-(+�����߼ok����=��X�   ��U�U�����1D8� �Cm���#.��@��P��Y=ё��S���}���.�|^���; M�j�O               ��4�"pV"��c�W�RWr�������\�s�Yc�  �Ҳ5�U.�\,�  �b�q�G�����N�7�y���=iAY�u�_�����.�T
�4�L(              �,��b�N{i��ޯ~�ɗe����B�[�Y�j��1K�?   J�ߚ�S  ��y�����0�5�"��ƒәh������]l�E����yj�               @oK���L�3:���2����+wb��4��<   �"`����� ����1�X���ٚ��R�	���T�c��=�������O����
��(              @QXʾOG�����'����n��Ě��n����:  ��qA�� @[�����
������d6%}�ɛe�ᶇ���|wScͥGP[              П}!�_X��㑁�%��xl��խ�$pD��Z�<2��	   ��z�z @s�b��x�T��KC����o����>��] KWb���l�R��J�Tԋ��H�L               �d�q7C����d�i���D`��⟇���
�$�,{';   ��g��Ϲ�  ���o{�UQ�����ݪ|I�Y�����?�[���WN{pY��%ʹ�,
5ʱ�~              ������Qf�~��mg�<�gV��?kj��@���B1   ��c}B� �=C�r߄b�Q���F�3��{n|t� ���oC���
�ZA(              @g���������*���Ϙb^�����     �ң4��8�h��i�@r���Ls�o+���;�9P+               ��=�s,20��-O�(��<x�Ϝ�Ъ��y�����     Pj��b�ޠT��gD'n����H����#[jV�(���               Z#��������	����C�.(G     ��(�Lp�`b"y��������׶�ȭ�|p              �+�0�����KN�� �`l������Z�1��L�      �e�J��9>=�O��0����$o�}����               tU�	������y�cO�O��ǟ|�܇�F[CMA�R>k̳Ǿ�Ԍ      �4(Ŵ&8e$5�-^��?�éӿ�`xmxq�@�&���d̬               @/��qwLOl�Y^Gw|���Pӹ�챏P     @�P�i���KdRID��u�����/�\���i��e0>!               �{ܝ3���� �c49��uC(�-�ye�[      Pԅb��;�#28��-{�R�u��f�n��q@���P              ��Z���x6i���ud��_M4�����      J��PL��Z��prr� o`�g�D�"f�<�@�FX               ��y:�+2<��U{���{��n������jJq~     @iQ���ꍧ"��~���9�];�6��Q�T�7$               ��<�1��+�ILL�_Y��\�Ra��     ()JB1�aH��B��i��F�M��0��ڻV�<�R,�              ���w'L$�?�$L&�OZ7�bc�;     @iQ�	���1��FS���o�I� 'a:���Q.��               Z����%\��pf��Ǭ��(U�%     `�ַ���Y(v�\�K.�d*��$SEm����NR,��m�����|�              ��0���Q����� 'ၛv?}ٷO7C�!P��     ����W�t��=�����x %���1���$-9��y	3�򳈮P�[!               �O�<��OL0���y�e8�     ��l62���������h:v@����֖����/6�	�BaoH               ��
�O|����x��Td@�9�^3����<����$     ���Q��i�z�b�	�8"�I�`�R�q�P�Ba�               ��b�Έ�����L:�cݬ(e��C(     �;�4C�a���ń\�z�L�Y�`*�n�����              �M��=�N�e���h*��9O�c      ��a�|z�C1^���ū��W8�� sM';��-e��� 욘               @^�W�^�L�`���'P��f     0��� �C1n�Z3�x����������(eGb�⒴d               z`��3R��1� �J�����      ��B=�a��bX@Rn&O0Gi3K(�����               ]����h�� s�N�f�      ��f��Q����)	�x��+����Q*��(�5<��               @"	�eͬtF��WƜDf���b�!;A�,x9�     @ØW���f�v�$�u)yX�J2��B�9��@9bY               za�z�l��Ӷ'-�<��p�C�^-�O�c      (w�����LӬ,��\.�C1�֕�f�,�c�2����              ����PUKg�� oBZ2�k�(�     �]6�]n�[�r�\�z,%+=B1�e�$�9˘��r��               z��ߩZ��������	Ũ��b�      ��ܑ;v�����)�43̑�4#�.j�               :q�K�VV��b�d�Lֺ�T!��    �rgƊ>}G>L�JOVX�UΠ���s�@���               �=�`�;���v�d�V1  �`^�<�w뽂�c�f�\:�R�l�e (Iy� �;�cǎ�I�w��p:��`JB1)3-P�-�1w�[B�RY�@               ���$(�7��)��kG��� @9�z��o��-   �����iI$o%�v����|0%��4Hʹ\�b0w.�T
�K�A"              �V�㮞��"��7��kG9bY  �'��#�P�@  (	>�O����b���\|���=ǺY+��f��M{>SIl$�M��n� s�1�j�r|�              �����sy�}�M�<�vc�;  ����JUU�   �����\ozz�����|�;�n�l}��z�z1M���3����}�;�N�nS�T��)�PH�U�|̑+�Y,P�1              @/)"	�y]��]ۛ�v��!N�w���c��st0Ĳ  (/.�K*++  �T�Q�`0(�h�O��=����x<�J$����4�і�2zQ�:6�^y�?�ꪫ���JB13+P+��{�#�˽H���               zI�q�')+�B18i��{�@9.�
 @y�O�6C   JY �x<.v���^i��H$.�d2[��%�h�%��|�ֱY^K4JB1Dԫ�T��Ɯ�ܞ�r\q              @/D��s��Y7��$.��r�q �|؁��'   ����K$���b��oё��}<ߏ�&��r^�G���+���#�$�˻H�T�̊)yz              �-J���>�g� s�s�qc   ���Qr�0  ��t?��#~.������*��$��]�����*O�P�b�L\               ��H�=�N���0!O`�@9�@  ʇ��  �r���O ��꫻���JB1S��@=�ۻɺyH���V���N�               za��3��R� ��/(� @�0MS   ʅ��>>��V�K(��Uxk��:oe�@��4�              �nf�qɚYqz_a��U�+�0Uފ�R��5��  (�tZ   ʅ��>�@`�ꫯ�G�c�	�JpD�7�F����/m_Z�r��$�              ��\(!��7(P��W� �4�k�JM�c�P  (�l6w´ǣ��a   �$�Iё��2}>��T=��P�G4�����U���	�c�              ��d:J(F��@���9����?9(���{.�W��f��� @���bRUU%   �,�J�y:
����k~���,�ٵa�4�0�:��5;�v�m{�U;��Jw���XD              ��T�}��֗���aݽO�7P�q�睨�w  ʏ}Ҵ����  �R��f%��n쵮����_s�5��|%���i��f�R�� R%��#��ԟYw�!����6���D               -KpF�Sq���I�t��c� �<١�4%
  @)I��233������񘕕���ꪫ����R��S���zB�B18	*Z�M�              ��g4��[8	��3�M�c  �S<�d2)�@@�^��\.1C   ����d2�H$r�7���������\q�?q����b�R�2��N�VC |� o���_���
�O�               �3����0X�@���(P?O��x�� �rf�T��  P����̟?�=]tQĩ�U�����p�@�E�����JO�JJ����               �3���W�{��u�Y����x����Y�r����     @�؁�P(t�����|�?w����b�,�;��W����;�q�#���@��#�               @O�q�y:%쪺޺!��T�����q     ���cVTT�X]]�\~��{
��P���q��Ni�U�w�P^��P�
�r���2I              �~���y��x�����L0�     �Y^�����]��WZ[[?��w�k�п'e��j�Y�;W�װs����������wd              �k81)Y3+.�%PkE�y;�v�m{$*������W�k(gZ_C�I     �s����xb����������Vcc�#�\rIB4�,Aq�9�+��]���k���W���ڛ� �              �������4��jU����9�	����:��S��(7��ʍ}      ��0�t(z޺�{����v'��;b�f��r�X�������D^���R�9e�{1)cf�Mm]9�ϸ�*�����e���� ���淄e���T��}_�d�r�}D���.zo��*.I�˥�g|�S��5-i>Sj�z���J �]��9�1*���m;g��٤=1]u�IgOLLS���u-�����#	9r|L�f�u|>�l��"n��?t�+��cD���
����-�;#^��s���H��H�j��qd��>��1C����PR��=�4���[��e�дtt�H"�q�JK�Is�_뵧d*-��cȑ1旪��V3-��"��c����R�u��$\钀���h,%G�Ge|�cH�����������@��O](~���ˉɸ���ǐ*���~u�����!ۿ�#�G�o��'��9c�5�����C#3r�{Z�q��ί�-A��i{o�56�0�T��g�{����̞�	9�ɭIB�5+����e���/c��u�0*cz�{JAQ�/���e/���3'���z{;�����	a�y      ��0��Ν;�JQ��#1v,�9P#Poq�����]�߻���/p�`bB�����q�j���i��ʎ���,;g���A��c266�e,Ǝ�$�Q�z�G���R���-c1v$��XL��r������>I&bZ�b�HL6���N�d��fٻ�S�X��LBF���'�{�*�ϧk����cH��.9��&$�M�r�X��'�ّ���)�u��B9�=�\e�/k����Ǻ���268a��ZI��284�e,Ǝ�Dcɚ��y���s�Z�O�r�Ɏ�t�Z����v�|���h$�e,Ǝ�d2���M����R�ɖM����ů��|v$�w`�z������N_&O?�n��yB��k6�������.���G{��_ڑ���	֥`/C�����_�2c���uq��-5�r��?0�e,fp$"3�1���VK��ކ_��4�_ڑ���!��Zp��-�?8.3�-c1����L�~��kB%��-gnY.�<w���_ڑ����9㴥�܋bf��_�w��z��t2��tb�:�p��n�8����pJ�ߺ�m5�*,8��       ��<�&���@EY(��!��y���u�������V����鋎
^����23�q{��v�`;fͪ9xؔ�I�b1}�Db�V���3V����*3����[*[Nm��^��.�I$�qu�!�pJ�v�;38<n��c,&����c2B
�9�sKrG�����ĸ���p�1\.-c1v$�h�u�)�NZ��)w�[,f6chxQ��YǍ:�bf#1�)	�S6��H^�߭],��w<��s��*d����k����0�t��y�����b�HP8������B�b1����qY�:�b�����a�}"k;�lIc�V�X���L.���9�ކ�k��#1ǻ���i�-��z�����"1Q"1
}rƖ��bf#1�/��uˉ���:��n�'�7�~O��������u�o�����o��kC��<     P��<�ȳ�"��{ll̓�dr�UVVf���S'q�b�;�L4�4�>3([jV�s.ir�}κ{� �+�8%���cڣ��7�[,Ǝ��7Ry�4SkW͓��E��'ť�����)�'��BE�/�y�٣��P��KDb
K�X����)�b1��W�+eI�X̫#1p޼����%cGb&����n��WGb�<�b1��3Db
D�X̫#1p��y��N����_��MJ&C.��U�b1Db
K�X��.�$N�+�b1Db
G�X��"1�=�n�;35C$�t���.S�q���b��g���`Gb����t���)��[�j�ig~9'��tֲ����P^eYռ+�i�     @��?-���2����Dno��{ �����I}}�=f�hLi(�#�"���U/ڶ�m�gO�>遄�U�����#`��&�e2�]b1l�҃.�;��)$;s�酏��у.�"1��K,�H�t������N"1�f�b�Y����޳7����"1��/]b1Db��K,fpdFf���WH��bR�,�l�تE,Ǝ�$�1A����DS�7H$��r��g�����X�D$F�`M��%31��s��wʖ.��\$�c�z�`~YH��bG��%�����6���˧�4��=���韐D2F$��t���у.�;c2���	�Z^�x�����ͻ%({���U����!�     ��������v@&�L���b�4�>�"���՞�͡O��UP���Z�8���9+t,��H��F*m:�78%��:�H����H�&
����,�-:3!��B�bf#1�A$F���n��#1c������X��~uX��ؑ�c���/5Q�XL.�$>:cGb�{X{�E�c1�}�J��W�XL.3D$Fg�����"1�(t,&�%����b�������W$�E$F����ч����b~�kk~p�@�H�^
�!��B�b���б��n"1o�PbR"�����z��� T�9���e�����.���DӉܘ     P����������������QNY\�q!S�v����5����oN�b1٬�F**C$F?���ؑ��^����B�b���P��H4)��l��L!b1�HLǈ."1:)T,�H�~�X�;���ĸ9��J�b1���2�06h�P�"1z*T,�H�~
��ƒҗ{oh�P�"1�)T,�H�~N�bV:�!��B�b�F#Db4c�b�~�*�c1Db�T�XLO�$���b1�-�g�?�h,�H��
���6�&��7�4M��)�V�3N�Yv·������w	����ְ�f��Ǵ�sc     @9z�u�b_3Q�Ie����P����뮽�����ǿ!([K-�gS���#��7��X��9�9�F*M9��'�-�c1Db��t,��w�H������D���I|�r2���t�єӱ;3:a�
4�t,&kf�X��M9�!�/�c1v$��{X<�9�����Lq��fc1Ͽ�n7��HL� R]ٱ�_=}�:�wf�G$F_N�b&��22F$FGN�b�����X��xD�g��_j��XL�H���X̾}25=��ކށ)旚
����b����D,渘g�|\ �k'�Jw��lT}ɺ�A�Z`��S�	rP���     �$��[{t�P�Ö[�޺!S��j��-k��8�#��
�b1'��N$Fw�X�!��	��;#�5�b1�TZ�zFģ��o�S�;��$�r*C$�88���H�A$Fgv,&wտ���"1�s*���t؛�9�OgN�b���ϩX�l$�M$FkN�b��'%ɕ޵f�bN۴Ty,&�HI��'�i+�Ŵ�ўS�;3<6A$FcN�b���b1�c��&�3;�6{]��#P8�$S֯�/���XL���$��mЙS�"1�a�e��b���tކ���]�����W���ζ�M5K�#pTG�=�      �H}(&2(�7���zɒ��_t��ѣ���<������NʘY��ձ���A��^$֮V����h<�&�"0�y��c�l�#1��#�&ST�b:{�%�%ST�b��������Î]Uo����[U�"1��b1�yX�����).�c1C#3Db���X���:s"%ST�b�HLw�('�	ձ;c�)
�c1�3q�c��T�bNDb���	ձ"1����X�˕�b1���6ձ;�8EAu,&�$SLT�b:���M��5j���5wXw�����]��jv�9�xd@      Pz�/���8�e�dyx�.�n���\�낳6W/?E�(���T6-x��X�9g����u�������HUd�X��/�%���|�4%#SL�X̺5��;��3z�F��;��s�bJ~ǆH4A$��ر��E-242����� Sd�X�S����xot4B$��ر���D"��8?<6%6`;��sV�s/��c��M�)2v,fz&&�T�7�O�̈�ㆢa�b6m\"G���s�ޞ1"1EƎ�<�B�d�O���&F$��ر��K��0���ށaN�+2v,�ik~i�{~9%Sd�X��d�LLM�����'����K���|��^.֞�����IJ"��cONN�*"v,f˩K��ូ?vW�8{���yd��=��f�Db���Y�r������{���\,���b��<az���@$&_�E$mf��3:���u���>���{fecgێ��e���Q�EP�      �&�ž2ݓ[`��%p���%�w~�ݗ���������_�8��i����c�b���_��3�������d�l�$S�<^5c����ɽ_�S*E�����M���Wܮ�n�wO�j(F�IA���旼��Ϛ_zU�x=���%~ǎ�\��A6����Q26�&��(������i>+/Fn����؟3�Q{���ؐ��8��uY�
����Q����P�|^���>f&C����n�!�_��y���DH�)�I��YU�@��z_س�]{�u�hH	��h�W���aǣ��p�4     �R�|��^Xj����y��׆�%�Xw	Ŕ������͵�V	��S               P<Lw�)�3�V�;���7����k�8�ukݪ��w     ���H�y�t��XY9��cw���ۯ�ӂ��!��n������S              {��{�-pV�7�Zh�w���(��*o��`�d�      �49�90�%U��kW~��۶�Ӄ������~�m+*��7���}              �x�CEa�Y��o�p��?��nAɺ��^rz��͂����     @ir,��h��xV�<j�=WP���s���jWTP��               ��hbJ��~k��<�[N�]���m�ַ��e%��{u���?d�]�y��6��      �&GB1C�I�����]��k�|����oJ��ݵ�*V��P              @q���65�)���j��=��u�
Aəny顳*7�

�=�      �͑P�m�t�l�o8�m������v|�޶G���qÝ�~bK��5��90�":              @1�c
�j�((�s������_z��'�����ؾ�܆����`�      �6�B1/N�m�b
�5��^8�ۺ�6AI���Z�mX���a
c2��3              �����1A������'"muM�=��mm�<����0h��

�q�6     �R�X(�ٱ#b���(�s�ם{�]�ܲ���n�U��?��U9�3�?���Q1�/               ��ب���d^�NP+*�W����u�RA�;{~�VU.��@|\z�     ���Xdb$9%�!Yj�a}�[w��f�H<�՛�<,(Z����=��z�bAA=;~D               P��?"UP8okXw�G��껯��Ek��\{nú���8��      �:�B16;�@(���}U�ӫW<k�ky��ᤠ�\��K��ָ�C��2��&�	               �׳c�b
�c��u�5~[��oy�EAѹ���ok<�n�����C     (u��b�����&(�U�j�N�̺{���\���k�Ѵ�_�.Gt�'�TD               P�^�l�������B��U��4,��<����U{₢q���z����WE%��Rٴ�<�!      (m��f��H&.!w@PX�֭=�{�{�m�}�:AQ��m5g4�x��f]v�
               �-�Mɾ�N9�f���VVί���h�]#(���YY��FPp{�:%�I
      J��������&������2C�oܴ3qg�Ȯ��@kmmm.M��C-a��%              P�}��b�pz���}��?���_&����w�cg֮� �{�     ʃ����c��h�c������Kޑ>r�M?��@[��C��\�v�@����               ?{��Υ��a[��Kw'��_>������]v�;��_,��o�      J�㡘�=(]�#)A�<ƅM��C���q��O<&�Χ���'ή_{�@��/Y3+               (~��Q9�e�A���M�o���N��_�ܸ�O_ؼ����`�a=�     @�s<3��ɋ���ڕ=T{��w�l�~���/���_
��{��[�lZ�@+?�'               (?�G(F#��i/j��?�wH�Λ~�wm�p祟�������?��g��q     (Y���	���v��r�O�;�w��O

�w��7�k�x�@+��?�%               (?�+��|1C�;��e�K2w������.����S?�#��_��     (Y����A���BAZ/����¦�v�w~���+(�����Ƕ�o�X�;t�5�              ������~YY9_���+�l�{�.W�n����Mw^ֶ���������^鋍	      �CAV�f�qy~�l�[-�K�7�:��w�������Q�ڶy�-���Y�k������              ��c_P�P�~<�[.j��)�=��ۮ��u��r�{�9�q�N�����({�     �I�R��":�=U{��w���U�.��;n��g�����7����Z�l�@K#�)90�%P+�HI4�����^I&E&�LK&���C�1\.1�YA�'�JƆ��_b񔠸$�3���̚.럆�m
�GR��೎ҩ��x��I���B~�=���`24���Z���^�d�7Uǐ�O�񨠸$)I���zp�ݒ����j%��旑(�O��~=�{��^�2��H��Ȣ�L�Y�������x�fV���/����5.���G2�T��d�/��/�I*��^)�������׋Q�z=$����!k��q�N<�n�ɾ��=��f����n��PL������+�$���w������/֞����^���B���%�7��W�j_�����x�tȧ�~��׸�}�\��~_���     @�(خ��FI�L��`㋎n�\�r������~n翿O���r�Ƴ��ri��J������Ǖ��R��9,-���Qhn���G\261.(�_���
%��-�W�vI�XLQ�����䌒����R^>�+3�iAqػ�GZ�J��vI{W��)�SbfRJƆ������SIb1���d���Z���cۯ/��-���b�DG稄*������
�����d���Lf���~%��c�r�%#cc���ʑA����a���v����.b1Ebz&!#���֞���#S��/������\R��~�K�t�p�N���T"�dlh�Y��.�ŉ�{~��^%�K�^_^�[:{�9ɬHt��Y�!!cCM�B^>�e�[X{*v$�C}2�I����1��^4*(G�Im�W��/�����W�$�%Pf�	S6���������8�;�'Muj�6�=9t���Ebd,"�XL���XW)/�h,"�߉�������'��%���=)4���C3���j�@?���;ֿ�yϱ�W޶��o�3!P��3�YU���i5˗�e�Y�q~   �B�d�=�G���C��1���:����}��+*Ԭ# �W�*-�L\~5zP�5l�ɾ"�y���[�@�c_��̯]�{H�w�����/����&i�ɡ�ؑ�c�����:���z��9xD��;ST7,��TȚ����n1���tfGbF%X�U��.kpظn��t�G"����HLu���	ۂ�p�X���H��tD|>��Ƿ� �Ni�Ɔ.I$�j��Nl�������?k��Z1�Y�"�9;cf��v�9�2�ʆ���� ��ّ��G�$\�W�kV4ˡc����btgGb*|���p@֭ZL,�ؑ���a	խ=�_�@^>�#3�/�gGb��Ԭ5ؚr����b������_�Z���t�by9w2_T���HLm��c�����F,Fv$&�L�ǣf��s6��Ɔ��d~���HLuX�ذzyS�Xrh�X���H��c*�Õ~9e�bb1E IHWװT��/�, S$�HL8�noC}]PV�"b1E��Č���K5ǐ�g��-"Sf#1��*�6T�a}�w����Џ�^$�9;\���������v�\�wW�y�[���di�YAY����   �0����������~/3��o����G  ����)��PL�T���>Z��C�s�M���E[[�+:�7��p��=����?�gz�Xd@���H̬�X́#Y�����+}RY��%�Y�P^9�C,FS'"1c�"1��X̦u��hNu$f����/�w�ѕ�H̬\,f�bb1s"3k��z���詣Km$f�}\b�b^>�!�4'��Ȏ�:��$�Y��5K&+26N,FW�H��P���Y�r��r�;we�Gu$f��e�Ƶ�ek~9e~�+Ց�Yv,�4��vb1��(��̲c1���wK,N,FG���~g�v,ƚ^JW�]�􍟈ĸծ=�b1�X��bt�D$f֪eM�@��(�]���̲c1��,����$�a�IGv$�Sa$f���:3ˎŬ�Er�X��TGbf��b^<�%1b�Zr"3k~K8����X�2?zY�]�]n��x�+j��?��~���'A�ܸ�ҿ�ְ�﫼.��ٔ��+    �w����7�yR{����������햚��\8f���A���	 �+h(楩v鍏ʂ@�@o����;������M�\���k��zV��AQ�a��5r����rf�bo�Z�r�<l���@/�K��#N폯�����Qb1��]$ƙ���X����e&�շt���^��rnak~s8������U�q*3�w��nI$b}8�����.wK,F?�HLF}$f��ٸv	�9���b�+������M0�ԍ�	8��U[]!kV�ёS��Y�X�:b1��kCV���_67T�a.�#�btcGbF�&�Gbfٱ���|��$��R+��f.vn~ٺ�6wK,F?v$&��+���
<�~m��=�%�tR��t:#_�מV/o���яS��YU�~ٰ�X������"�7�"1���?��cݒ5���dԡH�,���S�-&�!'#1��b1�t�b1�<�d���ra�f����e-g�c��5<{��?�C�ނ�m;�*{{�)�4���b���}�1   ��&&&����v^��{GGGs�JEE��c^����  �SAC1�ƻ</W/�P�?��+�7o|_������=x�Gsv���Ϸ7���xC֋D,��=#��O8���;�o�<9`�b�̧�W�K0��禹U�b�29���	�"1��XL���{$�d>]��Ĩ���Z�R��%���!g#1�r�����@,F���̲c1�aJ���@NGbfٱ�k���W�$��|Z�Eb�8����_��'��%�}8��e�b֮\l����h��H̬\,攅��@�L3�Ԇӑ�YM��bʉXg����H�,����)�]�k>{4��c1��R:{�����H̬��r�bb1�#1:��e�b�a�X�6���̲c1�����N�d�_� KJGװT����@,F?�_q63��ې�.���=��JPx�1������g��O!"1��T���/����R���%S$���ֺ՛��*�������	��;��8�f���8����    �{��G%�H8�\�X,�����G���zsјW�c����v�3p �s
��=1�\�z�x�l����%���5�S��/\��Nʇ��}�P�׬X�r��g�{%�q栽�ؑ��G���̲׭l�}��2���w'�q�g���*�lm�e��歽t�$!�sg��d2� 	�;���\Ba0!��Y +�,$���ֱ,��h�w��U�JK-���9B-�ݒU�9U��>o�Jǖ���S�=�}��2��MCb\i���肪���UѤ!1S����h�b�����D�Bb,��q�L�-���)Z!1����+�v�loQ�M�YND���r��P��C��4a1�v?$f[����Ú��a1U����NHLvdCb,�� K�����NH�%/'݄�t����E��Č��IVFt�=i鹆
��9!�k+��VH���8+�_�b� Z!1�����t���a1�d����F�RUU�K AJ�qh��h��Xv�b����m��͐˙S%~��/�+Z!1���4�?s��А���i�VXL[��2k�NCb�3��䲴(St~IXL�-��eff1�!1������0���h��X*���<wd�0�P�Z���9�Y"p���bW���e�Ͽ>�q��_�'P�s���|"��S�^^�C��I��    �������;��ޖ��i3��r�v�ctX�2��Œ��-  ����ŭUi^�'
Α��Jx]ɥ7���m�c��o����
���w�3q���_�����s�3�S��#��4I����o:[&��	�^q����d�G/$�RX�!g����(�vH��t~�+�;]c��N��h�vH���X��LXL��ĤD7\4-5I.֟��]#��D�?��D���r�D�$H@&�g�����4�UJ[����y���ݐ����c�����%At���Ԅ�/��S)]}c��D����ep_<�PNXL��uD7$Ƣa1-�#,&j��c1a1���D���'���g�b�'�!1����.�b��!1���J�1an���h��nH�E�b�TIa�Q��lG5$Ƣ�⹳��D[�Cb,�(7a�ܿ�����^H�E�b.4����D�Bb,U:��a��M
a1������5?(pm^�=E���X��y_����}�O/���C�ו���/wF�b�K�Z9'   ���ݻ�9�x<fLNN>�mw����������: �\��\�^��IP�C��T�f�?s�Ew�7f����"�w��?����$w��_�u�h=�^���qA��%$�b�b�4,& �TE����D�˼Q�b�H��qv	��h����J��9&a1�v�cL���@�b��0a1g��KZZ2a1Qb�">K͉��!A��g�e��KVF����������Ґ�����Xt^SW{\��daiQYv	���纤�T�t0��4��~H��
���9.kk���2!16���iX��\F&�Ϙ_F�	���~H�E�b��Wʝ����D�����&��qh�0���X2ҿ�9"��mA��)$�Rw�T��	���II
�f~���n�b:	��8��AH�e',�[d��g��K��/*����H�KH�%Y�6v
��T���221|f�s�X����'_/�	�y���������I퇏�������_���;��篽z6���sO�$P��Hހ/x��#    "ohhHb��Bd���$''g'D&//o'D���HRS�s] �-�Z�\�Iς��
Σ����pv�b�诲?5���3O�җ�zE�[��?P�y��.䜬�⹳}~� t�cїiS]��w'8nAd�-$�RT��o��h��-#���UH�E��/6T���QY][D��Bb,��r�g�Ad�-$�b����g��c��ԉB���Ԭ 2F����6��$+3̈́Ŵ�豁 �H�[H�E�7��Ǥ�Odj�b�H����T��/�3��t�t�뱁�e$�-$Ƣa1*�Ŭ�"�n!1�������(��H�[H�E�O����旑�����"�|��'����%[��X�Ŝ�����3��"���tO�*$Ƣa1="���_F��Bb,y��bD#��
��ל����Y���!R�c)-ʒ�@��� +R4$��6Xa1w;�dy��a�_޳UH��*8�$�=5旡�����g������Ԑ]Uz:�칲�.�1�1��?��_�8��?{�jWɇ��~<5�^�i8��϶�{��~    ���%��|>Y\\4cpp���YYY;!2V���X� ��w0��OO>/�x�Ε����ڒ?>����U��G�����o.�Z����^��S�eu1���{������WgnBû퓶�	�t���=� VW�{E�:�qn�sR��&k{-��������b��`'�<�208m���zl8u�T�n]\�!����&L̮�Bn�K

dd|F^K��woIRS�dk۞��k���삆��s����ֈdf���PZ�++k[2A�N��̮JR��$��2p!!QNT��Y��������i�cCUy�,�n��nã�R\��=痩��R~�4�>1!z%᳹�ޞ)I��SU%����uAxu����4������HƧ�qh�յM�3��U�^{:&�}GB�zi�����,Y]͗��9Ax-,��+5A���~�=_{'+��̼�/������r뎽����Ž��Aqݫ'"�&��0C��9�LNN���R�7��2�4���k\2l|]ڬmXfmC$��kD�m����49V\,SB������HZ�}�'�J��K�6D­;㶞_��k�/C�S����J.
�#�+51Y�Ya��K��.z~la�?|�W��8�~��OU�<y%���i����i>5�m   y[[[��rwuuՌ����%''Kvv�NxL^^�N�Lqq���\
 �`�����[������f'���қ����]��K�9�8��X���s��w2��o�ϭ�I" &f|~�l��y3׉��Ve�q���x�ƈ jxt�@=��� ��g�@��p�m"mȢ{C��-�����1������w�P=��f �k�@�n�dum��%v4�0.��7�b��y���o`x�@1��?�k���Ҁ\�?-p6Hyea�y[�����k�3��~����e�a?�ǯ{eEF��_̯y<#)����Ǥ�5�  �h���<��,..�18��kiě���"c�X���� p0�	���o���OV�J�R3����U�}�?P�1�1���~��?&1��������,��S��r1Eb4(               ��S�&(&��'�������y��T�d�����_ṱ���w>-�_��W'7�d�JuF��r��i�{>=�    �YZZ2ch���.��E�1yyy;�2�X�f  ��&(F��T��h���`�?�H�ׯ�i�*g>z�����[������o~��)��w�3�^�-O/�ņܪ�L��c��ӷŽ�&               �_�܃2�vOj2�	bGbB��˭.����������|{z������,��?�K��Ն��W��P���֦���    ��J����199�����$���1�1��1V�LQQ����
 �[] \�Z�g����,�M'2J2�����s�çF=3_����ч����bSo�����3�XZ�O�f�^zE�+�1-���$I�               �N�]z�y���-�M�����W�����W��g=�kSߚ�v����+������gAr�/�d��*W�K�>5�msL   �D�����E3��r�v�cth���X���kl��"�J��4��LvyAp�)��M��T����읅��/������ۿ2�?������yNZֿ=����S���3���!�������               ��L��T��0-G�*]E��x}���_��󾡵��٭�/��?��_x�V4�lo���]�J�xsqj���,�-L͡j��\6�"    ��<����lKNN���l��1cʔ���� �4�;r�������gu��Q�Q��>��o=�T�ƽͅ�����+��oz�/|��	��}�;_�\S����I�o�Jr]-J�n��()�Nq%
��'ƾ)               ��|�����N�� ~hKpha�����O\�ύ/m�u�z=�^���ғ��Wo��g�彯���������ߓ���X�^TY��k��D���X    8��+���f>���r���a�ʤ�� ؑ-/���3򊂳��@�����4���������ѻ����_�z�6�����z�|	�Y����߿��$JRVR�d$$$&$&%O$�$&��&��RRJ��\�rS�r�Rs�Rm�2@��X��1               ,�{�E~��	)L�ħ�Ԝ��>��C���ɫ���Ս孵�U�gzÿ=���No������>�V�7��N�%���yRrbqb �8-1�XJbrizb��dWiNJF~aZvzfR:��1��b�A    �+8����c�����v������32�c�	 �b˄���{�N�ޢF,y�����%�|zB��g               �m˿-������	`�@�LW�K\E��Ӳ�$@�}<x��c   ��"$�<,D&))IrrrLh���hp�(STT$��� �bˠ�����Da�$&$
 D�w��wuB               ���x�U~��	)M� ���M�|y��     ����������lw�\;�1:4HFe��8
��Lx�幹v���� ��#��
               �o�'������ ����>'�~�     ����199�����d���6�1��1V�LII�� c��GF��W5IRB� @8}c�C��	               �R�2}K~��{�xz� @8Mo,�Wgn    {HII �^�,..�188��m������cdtX2V�Lzz� ���b&=���myC�c ���婱g               xo�'{N�s� 'm���    ����l�b�����/KKKf��Q.�k'<F���X�2�8!!A �>[Ũ�F������DR� �������
               �r�6sG~��{�:�T  ��g�ٻ   �^���eaaA�h�x<fLNN>�MÌv���Bdt�v �����M���ķ单� 5�oS>4�5               ���_~I�}�- ����/�/x�   `/�������^���Κ���������� }���  ���A1�cߔח\���\�P����eakE               ������,t�?+� �����R�    ��'Nȝ;wp"��c�����RSSMh��Ck�����D`����o˓�_�_9�c �2��(���.               �a���/ɕ�Ӓ��e� �����"    쩡�A���/��֖ �D��{����l)..�	��&���. "�1W���k�:~UsN ��ޜ��{ũ6S6%m;M�����)Y*`õ!�[ɒ�s�)�%Aĝ���|IHHķ���Y͑� ɽ�Ο��ՌU�Y�`)gI
�o�O�;_�O�S�%}���r��h�H O���-S|)�8<UX�^��bV]�������~�3ݒ��/�r���/�KB��e��%�d3mS2<赧�E�s�I�A�l3�����/�����5�$� ��������sq*mZ�����c� ��L|G&6�   �=i ���祵�U�x���b�����222vd������=�T���/ʟ^�y�� �m��|g�[���|�\m�*�-� ~��蕩�)Y�^����k-}MZ�Z$5�*�گI��1�y1]Hu��]Y�]�ӣ��b�B����Ι;���)��.K��b�x�O�Kk}�Yx{�����k�hҜG�~p���Y�7�+7�n�V�\�*��LA�(��ccR�Yn�#96�/�iil����^{J�T�4���d����ɩ�SR9S)�_Z��B����n�(�_Bz��-Y�\���z)],įقY�^���+{.�4����E6�7�J��Z�į��2X6(��R7T��2�m�l�kO���%m��e�
zN��T�TOUK�d� ~�\�f�MI��ʵ�6�3�������]?\/%s%
�1���K'{j������ 5[ �(�����c�    ���׾V:::��� ���u3���ؖ��$999;�1&c�Ijj� 8<G�e�_���g���K.
 <*_�/9�%q:���r�E��_��M:�ŝ���.�.�6O�K���ڱZ[ơ5ך�4���[����S��v/�R�U��k�ŧ��9i?�nk�ԍ�r��$���7���f�MYO[7�k�A
݅��������M�Z�]��go˅�& �E�9774�7�k���䕮+��N1_<�;�'E��D�	��/>����F�ѷ�������r��e��B�*ė죘/NY!�j#mÄI��a1�&��[u�dŵb�w�tI`( ����!�ׂo��tKk]�\�,���fw��}A���V��E�=��R5]0m��0ܠg�R1W����ҵI#�x��=o�ɛ1χ��7�K#�8e��*=w�s�ħ�!�������,�-ğ{E�������)�oS><������R �(>8�UY�m    {s�\��?����O~Rn����dqqь���m�5G���&@�
���d�sF���Kq���}Y���Jn
�<��L|G�צ%h��.���yE�<�ŋ�ݜw�,�4;�ŗ��,���b���w!��b��dus�M��4,�b������nm�����Ǝ��nλ���r�����	�ij6獻�ַʥ�K���+���9�F1_|ZM_�ֆ�}M���M�N�f� >�!�P��v��Z6R7̹�^{J��y���z�����}�[��~)���/�����@�������f�j/w]�D?a1�bo�E�i����w� ~�qA�[�6S0c4�����cw�E�6�s�Ϋ��a�W�0kNw�\��6X�pΌ�ď��%�]{�E_�J�N<�Bj��5sϊ�
A��*������x���1� ���^��L�    ����(KKK���O<"}�,//�1<<�����������͕�D֨ ~9.(fy{]�z�+�k�� �aMo,�Sc�J��"�˝�%ۓ-�q	"�\He�)�jľ�Bb,�ŗ�ZHe�b>-�;9qR�vwsދb��b�97�S7���?�vs��t~��n�w��b���h����y�[gnQ�'L7�]2�?��v����rFp~Y����
*��qU\t~�u/Bj��/����JGMǾ�t�a��ۘ_��;�l�)���n��5מʧ��M�!un�s������k׺�I���e��J�2�{CH-wO�5�Bw� ��T?BjY�]��3����DPq�/�t�����uE��i������CH-4/���Zh�_^*���_�/��T߫�6}�?6.�K���}���=�6IMp�} Q����>k�%    ��'�0a����essS �����ݻg�^III������� +P&55U�X�ȫ�_��%�.>'���Z	�p�����ےX�])�m/��y/����|޼��j{诡�/>��B*�ȱ�%���(�бl�x�tZ{��O������� ^���^�3_�_*f������ךkMn��4����b�Fچ)�|���)��;'����*��YCH���봘����r��"�|1�a!�����Y�v]��u:�Ǫ�!�P�Bj���VPq�67�c�^O���V����U��vҶTOVb��C���c�;��t�?I�^.���v�M��d�D8o�E&���CH-���r�lp~���2�d~���֥�K���+�M���v�mqg������
Į���Zh�^.�Ԣ��g�F8��a!�N7������5 ��ѯ����    p���&�����^:;;eaaA ����3�7��^o���|Qx��XGvv6��x��
԰�����Jb�)��ѐ��K�˴������rݜ��b��ڶ�a1,��9s�s�^�.A1_l;�B*�x�l'lK��|���9��|��]��/F�n�7^6$��_�o�ҙ/6=���^��{���I1_,�ߖ��� �|�b���rݜ�҂��b��w��9���ȕ�+��F��Xs�R����a�A{Bjѹ�����x�㒶E��X���D���1||�NNR���*�d�d�@�VCD��5˵��c�ACb,]'�L�o�\)��s�R�;�-�u�r����XtА˭3�X����!�8���_j�����z`A�9H��F8�MCH[�Zd#y�@�~�lD|)4Ez��t}C,���7�E�R�Q" pc25�-   �\�׽Ό��UY\\���%q��|��:�: G���f����Mw�������yyyf;`w��K�7��#���Ϟ|� ��Y�^������ij��bAl8h7�r�����b�Xr��t��>�/�v!�e�h��ә/v���^Z�g[�_��m��b�au,t�A�ӿΓ�/��y/����<o�"�~�^6�8y����)�~��S�+�XoBb�c1�|��r��b�Xr��ݴ�S���V�����6ܔ�����Xf
fL��	*&�4&���1�8\7g�h ��/]���
����ACH-#�GėL1_��ꑩ⃅�Z�>�t�;Bj��6�3��`BHO痹��_�e��sO3��3���!��'�hH�^����ah#�h�[Bj�Nl:l�E��>Q;Z˵�2P1 ����������?#�	��x8�c�Q�ge��k�    �+++ˌ���}�{<&���"&@F�e��}��������Y3��r�^ ��1V��>fm=���+�>3�yUQ���. x�?�������:NvHCB��s��p��漗;�-/�}A�y�U1@���GE1_�xԅT�̧A3MMt�CC2Zz�n�{iXL��f��vU\[�9�'�c>c�3_�0ݜ�s x&p��:�ǈ�vsޫ��w��f)�s��vs�k�u�����$)�$p.����Z���n��M1_�x�R��նQ�#4�TC$�)�k
�/;�J��b>��L�4ř�:��b>��h1.xh��Å�X�������&,&u;U�l:'hihy���_�/�$�TMU	��QCH-8t��\�&�>�f��QCH-R?X/���g{�R���B�I�N��!���'v<j�E���U�Pa11��Dp~Y�h�K'�Y��߻!���+ ����c���~   p&��Q\\,555l� �����P�X�F�~�crr�m��ɒ��mBc4<F_�:�ynn�$&r����j�/�����Ʌ�()���_F�Y薯ϵI���3Ig�l�L�LG]HeY�\�ֆV:�9�.�?6.�G�^�9�QRY�r��w�����蓉��#}-�k9�"WگH�f������^t�s>S�s��ݜ���-�� �4o����r��v��#���~�oU�T
��Q�9�e�o[L@�����W|�,�?*��w��P�LG!�P����ر�#��uE��)�s�ʹMinx���D�9�P��\G!�hP���\m�/��_:�QCH-�e���R=Q-p&Bz����xi&,�j�K�2!����}��CH-]5]
H�|)�pJ��Z�Z9�Ԣ�p���1�O#u���c�=��h��|�)�f.�s���F8:?in��C鿟�3h�y�yr�i��V��� �gjc1x���    �nB��:����|����&c���ssss��u�5a ^��9Y�����IJJ����������׳>OOO T��2�6-O�|M~�� �Z�^�?���W������|�\�,G�漗�ַ�"�b�G�tˏ���B1�s���^���,�|����n[��鶥� �H�J���P��4�������Gg>�2!1�we1�h!1]��AR�:�I��ߝFC��O?z7�*ė���j��������~�R�����(�s��<Pq�RK��6�������Fu4�!����-!���u�K=�$w5W�,�u�QwCBu�H��t~�4�D1����:̼"t~�|�ل���\gY�^2�p�2|lX�	^9=~Z�,�Āܪ�%+����X6R7��\�	�J��%T!����&l�b�B�,&���!�w���).w�ǉBBj��s���6�	�چ���>�k]��,&����!�N��m��v���ᅟ��� x1_�/�����bS    �04�";;ی���}����	�X]]}Q���ll��f��i��K��(�˵�C�d4@�z�Z\��bԧ'���y5r5�V ������Y�Z�x�W�'ۉ�R=U-p�Pus�K�u���CKh@L(RYL1�P���S������|Σ��9�7�����*��.K�z��B��y/:�9O��9屢����.�گI�&��N����:C�}���}�b>��'��f�MYOMH���5Q��$���RKWu�	$*�-8�	�	�����y/S���9�|����ܔb>g	uH�E�FK1���:�ԢA�Fz���dlf�a>o^�N��������kg���A�MhpC�BH-z?��_�doL,a�y:�?6n� B���_h�� ��ۦ�E�BH-k�5||�38�0�t�P��Zh��<6��tJ�&��bk���/O痹��_:M��||��� �����K��    @8h���
��z�;�1���d��t�s��Z�crr�m���cBc4<F�c�@���"IM��/^,&VY���}V����%'�Ee ����w�e�W 2\6ln���<)��Pws����w��ŖN�]�u�t�t��2})泿p�X����ۖvs�_�-]xK1�3�+$�Bg>�u7�t!�.���A����N�{�C��y/���c��sjhCH-V1��6�b�N�!�ˇe��H�~FoU�96T�����B��y���53���y�b>�3!�'�d&?�!�-�c~�8y��fؾ?�|��ҝ������Ody��6�?'�5�a���%��K�I�PמlN�!o6�>�Բ���T����6�W��4�Iږ��j��m�l�kO�Z۠�K�4�p�O�I�#��B#�Р�����}w�[n��M#W�Si�cy��!�J @i@�     Z���w(jjjؾ;HfuuU���Mx������n����Y��+��g^_:�'��O��V��h����'f*��V��?'�^�� #k3�����d���Ylyz���v�n�{i1�.��3���n�E�[He����vR�������X�c�`��i��3�YHE1������^Z��~�]���XliS������	~hgث�W%ӓ)����Is~����|�>���Ϯ���y/-�k>�L1��U�hI���W��k����d�97�/$Ƣ�%��[$BH-:������R�=�;��B1�������������*�;/K�'[`O���I������i��0� �'m8���"�a�9&�T�!ۯJ�v��~���1n�Ǉ�ϣ�}m�l��l��v���"W:�H���vdBHk�BjѰS�(�+%,Ʀ�Bj�i��u��b�
w��~���O��.�M2�9��Ƿ%����96    �]��y)�g'�B��h�����9��
O�C ^�kN������5���m^�%%%RTT�"���+��\O�E1u���.���M���� ~m���޿�-����Ƌ��"����^���y/:�ٗ�Fu��t�t�~&�|���T�̧�-5�b>{1ݶ4$&+rݶ���q�Q����n�{�g�S�gS��漟����}E����n'z9~l\�"�3��j��.���pws�K�כ����K�����G���Bj.6�'�(�3߫�E�u5�k�k�M$CH-Z4
H�<�|v����3w"��(泯H���v�ᦹ֐��'�=���H�)�o�W�������迋Ah������R�H5,Ƶ�؋�����?$�B#��z���H�m0k)��`~iC�!�tWw��'��O�BH-�N�p�(��[u�	!u�{��/�/��k��t��2�1/    �t.�ˌ���}�[A2������l�dv��v ���zw^[���/ږ��$999&4F�c���v��
%-���NswO�j�Kr.�T��@|z��?��Z��f�x�,����]D:$�Bg>�1�j:L @�i1�$�TOT�!��,�a��|�b�m�B���/��8�!	R<WL1�MD���^����U.wS�g����(泗��c2X6(����u_lhғY�@��9�?O!(泑�[Ou�LD.$�2R6b���)泋H��Z��X�ITL1�=D#���}��|��مs���\��b>�1!�����ȅ�X4��|�y)p�/!����i�m�CP�-�s��ȅ�Z����f��yM263��s"8�,���R�l'lK�k�"�!�=&i#��mW%���;0!��������/i�c?K9Kr��v�.�p�'!�N���m��W+�.>' ��3�w噙ȅw   @4YA2/E�-VVVL���	������y �e�|>�K��(}�Z�1:4HFe��ԓ�W̭���m�;;?*r�?JF27��x��l�|~�Y�p��G�RYv:�]��|�d
uNEg!�e�ذx���@��9�eu��B�_� z4$F:�2֢�g��3Ig�l�L]��漗�Z8f:��	���Hws��|��|c�"��y���9Sp������n�{��u]�����Iu�j�d&o&j���q�/֎�rl��h��Z��(泋h��Z����5�ʙJAt�̚p�h���>�Bj��D�P�/�K疃�!�,�,��3��B�I�=E�vʶ�����"�ϯ?�J���d	�(8�����5�1?;�O���k5}UZ[������r�E�u\�ԭTA�D3��B#��{�#Bj������e4E3��i���sr2�TNd���2晓?��     �KNN�	����y`��hX����������Y3���c������uj���WUUIZkB�-�bԸgN�����ku?AJG�צ��?'8S�w����|�D�vNmih����邪+�W��%f!U�]m��/�/�c�EK��9��zl�b>�b��,���i�n[�����P1M��h�f7罴��F����(Zݜ�c�A��Bw� :�N��D�D������R�M�!ݡ�|��E��7t��0�}�m�x�����=Z���L�u�Y�|F��͍�h�C�e�r@|�>���D�Tє���^��b��C�E����d����Q���R�;�-w���Ş��`_�$��E+�t�ֆV��sIrWs�g����\~��4�h��Zt~�a��گI�f� �L��[���R�p�O��;OuF��a�_���i�Ev!u�oK~��c�'���d&�~��oS~;��_�n
    �`4����Ȍ�hH���	���c��h��G�����3vKJJ�ӧO�k^�9v� :b2(F=?�%��x^~��	�V��[��_��:�B���|�XlivYHeѰ:�E��RY&K&M��|��n�{i�����t���~�����X�+����jAdE���^�EOԻ9��t���[2O1_D����w�pJ�b��v7��P�Z�g�9� �Ԣ�|��jjDV��9��/f~I1_��)��2||���E�X�TD?��B1_�������!����.s�*�-D�4D�.ܙni�o��ݗ%��4����7�o��2`�����R�.DP�H�){��ZL#��N��um��C�6]��	$��Y{��Zh�=z��:�!��D��BH�7ZQ�  ��IDATdbc^~����u?�=V yO�gdt}V     ����(yyyf���������������IOO����ʫ_�j����>�uFA�Ũ�����*��y,4b�^@�þ�ȤgApx�l���N1_�إ��~���r�e��d�ORݪ�%+.���X(�<�ts��t�k�.�:)��;��pC�R�j�l�NN�����9�E1_�٩��^]'�L�@��"C��w>�?#vC1_�٭Pg7��"+��۵��u��)�1���)��ts�k'����dlf�ώ!������A��9��BH-�E�	�	���Bj��5�ފ�
Ad��"���Z�\k&�L�Y%�_F����Ե�*$Ƣ� �/#G�wk�BjY�Y0k.�\�6�Yc�|޼��j�����G�yU2=���c��F8�7Y4)�'z�nv�_��m�D�CH���|�|b�����' b��ǿ!ߚ��}    ����f����]�b������b��?�N����g�5����DVL��~��ݟ�?���R��' b�Gǿ.��w	�N1_�-�ͮ�v��[��.v�םRY(��us�K�W:�E�v�47�{!�Hو�R|rz�@�p������X(�;vs���%��b�b�p�_��9�>ݜ���/r�c��/2��kBH3�{Cr!wA�ϴKS_A�af�n�{��t^�,O� |4�Ou�Bj��/2�r�|XF���]Q�9v!��W����jA�]U]2]4-v���v��t�UI�'	�g%sEn��;��e�P�/���/��2��]���r���p"`.N�k���ZZ�JWp~���2�LHL�=CH-4�;?6.��]�`�4]��;���4A��9��I>4�59�u\���
��t{iP�v�Y    �Szz�����n�z�;�1V��5� ��'@�{����@^��W
"'��bԲw]~���������&���.wZ��##\@S��pS�|L�,�',��P�^NXHe�b��ڶ�a1,�9;wsދ�|᧡Z��u@����q�OԎ�R�&=U=2Ul�n�{Q�~v��W�w���UBO�g7�L1_�=M�(��ŜE�S{G��b��rB�e>{�t~��/|���y?��&T,ۓ-=�W�{��3�N��T�P� <4�t�dT�b��sBH�e�l�́NN���	!=�a�[ٝ�-�-r��$�Y�N!��~[�(�/����H�!u�7$Ʋ����$�p�ԁ�ݓ����/赆�U�ȅ�BH-4�	���c2X怵�9O�fᄑ��v�����Q�5��$���;��    �L���RXXh�K�x<����3VWWM��>������M��3�<#���/��Ћ��4�+��=��w��87�2�6#������2����bK��B�I�,�.�jij���q�������	ݜ�Cg���H�0�q���j�x����b�漗�Yݝ)�-'ts�K��	������,���X6�(�'��Z(�B�pS���c�b�ξ ��<��2����y?��R�zN
!�hX�v�6�|a��R�|�c���;#��2R6"���=-3�<�_�:h~�E��nȵ�k��e~JK9Kr���8I��n�'��l�L:N
!��F8�7M eb�Aop��z�$z/�F8��R�p�C�=i�m��4�	��s��!1!�Q��o����d%s=���M�����k    �\.�ee���\[[���%Y^^��md��>֡A3@,������O���FAd��*�o̵K�H�������-l���c�^�-8�|��n�{i1_CB��S�ڽJ靴��B1_�9���~t���K���+8�ʹM�.��b>]�0� d����9�a1󅖓�9�E1_h����9gؿ��^�V ���iǅ�Z(�-�_�6�:*�ԢAh��r�����n����/�6S7���ّ�K��B,�W�S�#S�	��P�z:��Bz'/7�D�h-AR!`Bbj��b�sBb,z_����r��y	*���9i?�RKoe�ٟ˧�G��R��i��pBé!�m���Bw���Bj�N�T�x�8�pBˉ!�N1�>+���1yW�%%�{j��y>�����s�D    �'33ӌ����oz�^YYY12���j�>�Bet1�}}}2;;+��ł�����������& ���ے_����l��a�i�o�/E�h�����Y�)g�H�,�|G��T��B�iݜ�s��-��B`ݵ.7�n8z!�L��)T�����:Nu�\��Bb,����Y�u]�����sb7�(���YwS�2�ĩ(��{���焳�9�E1_h��g��Z�����U�t^�D��O��̉ݜ���|�C�R������R=�;���)�;s[.�\N�96<*=6t�t�Lތ8�|���R�d���|R7T���L��[�:�SiPq˹s�2m���Q���JGM�8Y_E�l'nK�T����񵥩ő!�ᄎ�-u��dm�ۤ~�^J�Kh�sN!��'t���T���6�'4t.���>m�ayO�g�W���c��i���}Nn-9{�0     r���%??ߌ����k����	�q��f�c�n��|��ݻw嵯}� ����_~I��
�r]�'���{=���Ug߀v-6�[�x	�yN��WoU�YT1]!8���M�z�E�NG1�9���~Lg��sR�Lg�GaBbnH,���Z�w���|���ݜ|k�`4}���P��(4,���3�9�E1�јn��7e=�yݜ�����u\�ԭT���J���%mK�d��𶓷M���CH-��χ�v���Q9���^';�>�^J�(�{�Bjqg��N�:�?"=o�8����L1_�%�]���Q,e/��5�`�`���������UwKV\�������|�\k�&����Bo���Z�ˆ͵Փ�'�gBH��Bj����J���d�96�Ε2�|�Bj��_>�';e&��!��M,��:�s�mR�Q,o�|� p��ƞ�����59    �=h�LAA�/��������������|aaA66��8�344$�����|��u}B�s��R�yL 8��=}g�[[I[�|��b�C���T���~� ��|�c&6ވ��T��M�tsޫ��M��d�b��X�X��ck!�;�-��ަ��b���~t�-�|�����:%�P��h�I~��pӜw�
�K\?w�b�Gݜ�>>l���Vʖ���BH�E��ֵ�do�ݮ8�X��WWu�	J+�-\,��X��;�|���w��H�.:g����b)��2S0cB���#���ބ�.�B����p�G��p	NC}�9D,9>"�d���Y�al�l� �X�_����R����ۜ7T���0bq~i�υ�t]a~y&��d����F��F8�&�BH��#��Jij����� p����LP     ��r��(+������,--�����l=֡A3@�LMM��瓤���;��"��\y��m�ot>%��R��# ���ǿ%�0�,�,S��x�,�H�J<��$�������H;�颠ʩJ���y���5�RY��O[>���$�b�=��S���Y�Y�X�8ڙ�x�X�򖳖�N��EZ�����|�yI���/�L7�3�d͵&�H��.�^��5���o���y/��´��:��@tn�ߌ�n�{Y�|W:���M���*�Bj�b�@R@NL��<����X
!���NV5�����s}�E�p9x������V3W͜"i1��i)�|/O�m��̼<Y�|y�y���Ŝ��r��L�4Fz&���M�H���`:�l�o�+=W�9�����!������S�$���r�R��y���5V#����MX�A��藩��
!��W��cC�a��!17�nJ,�����V��}��� �~�]sc+�Ԣ�pt>AX���~�^[!�N����9)Jϑ��5�n/��|�y)    ��222�x� ��++++���(���j�>֯i�s^��Ĭ��IN��k�����o.����M�����\x��d	 {���-����
�C���`P�ǆ� 6�7������Ov�~ +�+���@�9��H8���9�֥o	`�b�_�ђQ3 ��ι��z+{� 4,���_�>-��|��|��7А���V�D��i��t] 5P9`�������<�)��y>�����w��,M9�v׽2.���1��    �����%??ߌ��Ë5�cyy�Ƹ��>��_X���	�����Q������)�I� ����yo�gM�                Vm��MX̻ϽEj���=�M˯u��x|�    @�JJJ�	�y)�G�X]]���������!�1� 6�A1jxmڄ��Ϧ����t`/��w�{�>CH               �oC�{Ǉ�νU�2���Lx��u|HV�     ޹\.3���=�z�;�1���d��t��@�:r�0�>(F�Nɯw~D���fIOJ ���Ҁ�n�ߋ/�                ^,o�˯�P~��OK��H ��̦[����,n�
     xy��ɒ��oFMM��wɬ�����	��P������Zs`7�b��syT~��c�o���Z�h���o_��~�                �F�(���!y���JIZ� ����e����1a1      4v���������N�����:���dkkK�xB"�.����������� ,����!��Ώʆ�7e               į�M����'��M?%%i� :4�mOʽ�E     ����$���f�����k<�	�Y]]���e$c��,,,��Ɔ ��4�=n,��o���V�ŕ�& "�e�O~�����                �Mz�����Hyz� �,�yG��2EH     ��r��x)^�WVVVv�c4HF�[_��@@ � (fm�a�ն'�w��,��.�z�]]����W                �7��_������ ՙ� 2F�g����e     Δ��,���f����|��_�����KFF��5>�O�~�lnn��ښ	�� ��m��A1/�wuB�k����7KnJ� �gg���~Z|�$              ���V���F~������
^�kS���?$���     b�ì�������B���0�2��鲽�-�G���eiiɄ�蘛����-"����X�2���nz�������T������@�               ��V��o���jz�4fW	���X�_�xJ�|     ���5cIMM���"3TBB�$%%Ibb�x����h���������"@��2�<s�_�5u��r<�@ ��'ƿ)O�<MH               p \�?�?,���'�r�iZ-�}�;ݟ���    ��c�И��,3��ʤ��фɨ��M����۽&��5�Ff��"(� &=���_��?)M9'��g�>࣪����{$��&M�M������Dľ�UWwuWײ�������
� "�TtA��&@$��>ɼ��?�H�B&	�7��r�̝�D'w�������ޅ�"a�                �/�0_�m���Z����@�����zy��r�
     PLL����W�V�J\����Wa!�G�=�bܔ���#����vWiH��p�����>GkRv
               @ř7����I��/����Ԙ/l}p`�f�-      P�����"���s��$��C���3��-3�;+A                N��������ڏ���� T������kI�F      ���
2�hS�N�K�=mG���G ܳ?��:SG���               P9�'mQb^���t�����{2�9zr�ڜ+  �������
]&�-   �P�)����r�g��\�P�@(�j��c�\��	               @�ڞq@l|KOt�^͂��lqىzb���q  ��5Mk����+t���p   �bN�O)�t�7�X�k�*�� ���r��C+���o�:�               ��8���{��G��R�:@�V%o׿v�SVa�      ���P�i2�����G�������d;����y�!y�                �y9�y���9�"��nmu�|���E�"������)*      P����.��߮O�-��js�|�|���d�߶�RBn�                T�����d%��sƩ����]zA����֥�      PS��D�(6;Q�0N��������Q/�Z���               ��Mi�u��7����!����ծ�x=�m���
     ��	WJJ� w��d[�cu��7�P�1��F��$�0_�ٻH���                �K�O����-�/Ѩ�}���%�l�r�4?a��ٿXEN     TG����b�6B1g�#?C�n��+�Ӕ�����Ì�o��c��ڟ}T                ��|�S���R������c�&��K-��;?՚��     �΂������b���?j]����5j�@@md^�^�7�~-��P                ���S��u���vW�_�s�VkSv����R�)     ��.  @��Ŝa�YGu���hJ�5�a_yyy	�-̇��o秊I�%                �_ZA�����.j�Mw��\�>�j�|�S��[�	��NQ     �چPL04��g�~N٣߷�Bu�C�t˓��ݟ)Ù#                5˷G�kWf�n�ڄ4P���J�s;�*.;Q      @mE(�
�v�Э?���[^�z���K@M�R����|iC1                j�ج��w�ը�nj1L�>�j����9�B�,��U(      �6#S�2��zi�gZ��Q����AQj�˥�{ݾ�w�2�9               P���4?�G�cT��{���j��鱚�k��$	      8��Mi�u׺�uC�!�d�|��TW	����3�O�+                ���f��-�5�~W���R�����N|����Ykw�
      �-�xP~Q��ٿX˓����T������P\�Yq�+��               ���7�=�^�R��wm.���T7˒6������)      �lC(�ؕ��׽�a�ꖖ�(�/D���Kݣ7�-Rl�Q               8{$�g�m��-���h5B-C�9I��w�~J�%      �lE(��p�������t��j�_~�<=�z�r������&e�   J��u
���|k��$�           @M�>u�~��u]Ҡ�&��:�����qK�y�j��      ��(�T3��\����>��njy�FuP2�9�sp���ANW�   ��>�=��M�           ��L�c��-KڢqM/И&����G��f�k���:�����      �PL�u(7Y�l�H��ӭ�.U��hg���|����D�N><               p2�cJ�S��7趖��gݶΔ5);��ޯt 'I       ��PL5�S�.Ť��Q�tS���$(R@ep�Y��U��.V|�C                P�ج�����\7��P��PY�d�i���1m�       ��PL`�˓�ب�	�Ln1\���	8Ł���� uu                �`kz����=uo��ZӹuZ
8U��4#�Z��W       JG(�)����]C꟫�U�����r��&e�f�~�=Y�                �kKz���G����}h�ڞqP�|�U�      P>B15��U�o��ײ��uq���|5�'�$��"-Kڬ���^1                ΀u�{�~�^��w��i2@��[(�ƴ}���J���)       �#S�廜�"a��L�I}�����
;`��뛣?듃?�h^�                �Lr�\Z��ݎ�!�tU��5$�\�xyp�Y�ةY�i{�      �8B1����t�c��B�����0�,�R�i�A��W)ә#  ����v���M�-L^���            ��;+A����ޏ���j�_���@��cv��$q�>9�R�r�      ����eve���?8�DW4�a�]�$�~�2苄5�>q���B  xRN�:�=�\E           @����=53v�F6�{�a`]����qhё-:�Lg�       �>B1���@�|��־oԯ�9ٰ���i-///��0�/Kڬ/�hO�a               @u����G�i�����Z�女Q����'�EN�r����1Z��W.�K       *��Z�|Ⱥ<i�M#uI���AE��5׮�x[U����                jױ�u�{�x}�B��э��eH��:����G���#?+� K       �B1g�C��zg�b͈���E�����w�v�k��9IZ��Y�&�W|�C                P�e:s��p�Y��a�ua��� �������/%?S+����n�8        g�����U�I[�0���50��.�� �1��ѼT��خe�[�%=V                P۸\.mN���=_�cX3���Q�*�/D�>2�9Z�ة�I����~?      @�!s��/*�*�;^���GuР�.��F�^>B�;����ɛ�}�f�ʌ                �-�\Ev'�f���k�m��ƽ_d��
U��a~Hަe���>m�
�=G       <�P��*�շG����N���=���GvT��(��0�o�<���;�.u�vg%�">                �͜�B�I�i��no�	i���α�mH#yyy	gF\v�V9�k]�^mJ�o�       �G(%�+*��3�ٿX��{D��z��m���K�t�M������Mݭlg�                 %+riWf�3㖨�_�Ϋ�R��uP�z��$��tg�6��۸�v�Pr~�       T?�>����%���c#��O�Ú�Kxu
k�����(��u�'6;Q[�b�%#N[��l(                pj�
��<i��^�j�@��6�����؈Jw4/U���5�l���YG��      �zN�S��Š��
�)m��ױ����T��:�5WǰfjXW^^^:��iwf�0̶c���\  �j����I�&j�\M�4Uh@�|���c�]�S����tJ;���x�Oٯ¢B�f0���Md5�h� � ��ٹ��ed�@��IڣC��r��
           @mW�*��;$������������)�������Gg#��P����(�֌8�I�K      ����l�"��f�����ڱ0�'{�� �Ip�څ6V�h�����MT�?T��#?C�2��=v��r��HI  �
������jH�!�Ӭ��5�&�/���Ӷ��s F��.Ӓ�Kt0�����v�V]w=���;󕖛fGjN�����7y�bSbu&<4�!E�D�8��w�#q��B���{�Xl=PZPx�{{{2�ӊ}+�����O�'y�            pv8����&��ў���V���۷�mݏ6��U;I5۸o�n�s�:jG���R     TW�E(g�)���kQ���C���u� 0�À_�����1��H^����pn��Ä<���ˋ
  ��g6��v��<�N��0BA~A�|]��ָ����E.�K?�Y�n�T3bf�@�J�ݣ:����ʖ��nc(���Fo�X�3W�����v��lS�Yߙ����������R�f�O�:���e/��#��Uq����W5{�l
            g�BW��mܗk����|��2��ݦݎ s�ǎG���K�+"St�~$�g�Hn��m�S�?6b��(ә+      �,����E(U*)?ݎ����xL���+�7�~�^��a��_N�������K7���/�z~�/a�g����������,9�3����r�  @�1���z��'չa�3r�&BӳiO;�z���_����Y��*<0\�w�܎����n��g�{F�6��1��Ğ��%O�E��z��[��㉋�У��Q            ���6�����[�^>vǨ�#��p������m�Ͷ����c���������ۭu��������3
����:v��m�������Yv'��yi�r      �=�����P��wq���������z���"���"�\.eRD  �:6��Ƽ�!m�T�:}�}tY���X�o���a����3s��wo�:/-�Q�y�	L�qo�v�����j�9����O�PBz�            ��2A�C��vT�����}�� o_��R������e��       N	��
��Lg�=^|  ��cr��z������pA����z��7t׼�T��z�������k��������lX�a�h�G����u��<Z������c�*v�            ��R�*��6�      ��A(   @�e��3�����{*t���tmHؠ����K�SF^��yv.�/PQ!QjZ��ZG�V��]����zyyix��I����n�N�_���UG7��Qo�{��m�q4�V�[��;��S��5�yl^��:��Z^����r��qxc-�s�ƿ?^�,                    ��    Ւ������&�����1b4w�\}��sm?����~>~�ٴ�.l{��>�juo�]����/�m/O��"�"t^��4�� �b(�6:W3����߹\.�K��=o�;�ޱ�wYLfF����m��)�~��O�f}4���
�,u� � ͹q���~�[�                    �@(   @��ҕ/��1a�g�}F��V��z

�*v�����P���p�&���ЀPU���jڪi����\��b=<�a�)�Ȏ#uc�5=f�����]dc@�EbL ��E��P�!��ۄd�k�-���y�?5�ۄR���񷱘��֚�5j3��֢nPrd;t0�}/,�yo1���<߆�2�2���:��4O�7�WZn�P�� ����j`��j�F�"��9���M���u�h��/W7���7T�_�]&>=^�E�                 �g�   P��?�~�u�]e.c�!S�L��;���uo?�]wz���1=2��s�=6�P����f����/(�7����6�o��n����i�#[k�����.�KM�⦏n�'?9�uť��ڙ���m_j����T�r�y�d�'�=��gP��	���/�[W�w��5�vyOؔ�I�w.�g[>ӏ�?�e��z{��'E�L8�YD3��<Z��\���}���Em9�E�3�~˼���6���z7�}Ҽy���/}ZZ�'���k
�Օ]�ԥ.�sM�4=�2�}���yk�[�j�W              ��쐼*v�z��   �   P�to�]���e.�|�r]=�j�<z�nGJN���a���U�>�u��0Bՙ���y<�L�c�%1_�{�X��$o/o͸v�"�#K]&13Q#���1��ޙkg*��ϧ|n�%1�Ѵk�i�;���zM�!�z�%�q���_=����O�I��v+:4��'�L��־��>����7W�)�c?��H�Z�Sӈ�v����g>\��?���S�(���������n�`�`���ϱO���_-߻\��֔>SU����ꕫ^ѝ��T��V���Z��1c鞥�q֍:�z@              �b���"5  ��|||�t:���,�á���FQߵ���    �6L��D�|�J]f��%��(e�gU�m�M��ȷFjr��z�ʗT���8W�^�o=0��R��u��C1w���P�|vA�}�+3S�82�𖅥��Fu�	�&h���jt�n�:��`/&���v�p�a���\���Qm+���Sj=Ȏ�4k�+�\i��#[u�����o��	��#>��<h<�V?��}���˜��;Wh�!m�h�����~s���g�Y�ھ�                �V���6cFaa���󕓓���,����0̑#G�q��%�2�   Pm���vuiإ��]I�4f��*���ڻ?�k�����ϩ:{�����~�*, ��y����QaQ�<�nP]=}��e.s����c}��@�>��^���R�y~��y�r���+�yv䳺���
�PMЩA'-�}�>�����ߕ������լN3�)(,�χ~��Û=�>�)���߲��G4��s
r��=,�y���15��DՉ	M�bj��v둅�ؐ                 5I@@�BBB���`(;;[������PZZ������A�"   �Z՟����yg�S�̸F�9��G����Ru����y��iR�I%Λ�L��m����"�"J���~�f��y�o��+_��.����K�71.zqy�1����ײ�-�9��&2�3Jc��^]���.������Чy��ϼ'y{y�6i�V������I=��                �:���1���@��������UVV��<xP111�`P��   P-L�=Y��:o��7��

T�}��RC1���'B1&t���:����?{�Jn��`����j����W�2}؆*L��j��W�^jQ�������3�2l8eJ�)56㎨�(���jr�ɚ��D-ۻL��������0��.�[�4����U'����srV��d���۵��z��                �ʖ��c�/fdff*##CyyyJHH���q��    �Z���m�Ι0�߿����M	�ʜoR��<a\�q
/u��/و@U1a��b�ӭ}o-q�qxc��0B�o�\@Uh�\S�N�=nP����/����kҬI��~�j� � ͙8G�w�\g���u���=���oi��5"�                �~�1#55��`�HJJR~>;6E�A(   ���m�W]v)u�|iܑ�ܓ��T�|��<��7�:�_��WV�����e��-}n���W��7���Pθ��=w�s���������u�\.{X�k�$��Z{p������������Y�f�������uq��=��]I��cڢn�
]μf*�z��@�@]r�%vH=��?�_�l�D                ��[aa���ӕ��i�C0��OKKSQQ����    7�Ө2����=�}&�P??U���hh9���/�~���xU�mG�i����zP��&X����g�9����[�T��6U�^���|���Y��m�q^�����]�e����+q����0��u�|���%s�f\;C���Z�e�j*�xͺa�G"1?��A�/}^���>az�˛X��{�ײ��l���Q�+�?DU�YD3ͽq�^^�~���*r�=                �VN�S6�b�/&cFq�Da�w��P   �j�N��:���VmL�(��^p�2�==1Q��o�X�2gÜRC1&c�����<���ܹD��yd���{9�6�aDE��WhR�I6Sҿٛ�ܬ�������_=�W�zE�v���u,ݳT���:�ѹ�}{Md壉�����̣����������_���c���j�=��̵�s̹ctU��*m��[�s��w_�2��v�w�~g�3�-m��[Iv&�Ԍ�34k�,�M�k��~�L^`���=�c#5��                j���~111��1Üg�� �#   ����U�F]K��v׷B�4
+;:a�UmX�a���_�Sn[(��m��텄bpZ�F�U�f}�>����y�Y�{��J��ħ�ku�juj�Im"�ظJY���){��⧕����1��hQ��n�}�u��˯M�b��o��=�{4���m��}ſ�0��I�߳iO5y�������|�N����8�o=<�aM�h�b����cnn������L��q����͸vF��&��ܒ��̷��P���������s9����������N��H$�P�!m?�]u��G��,w�����+�?؞����mG�i������                �sL�8�R�)>m�0���Py�    �nM���˫�����
3�Հ2��PU�ޤ{�s6�@���s�����jZ�i��=�V^� go/oM�5I~@]v���6o����;}����Թag���|�k�Ͼ7����˘X����Z�e���bSb��7O��_������N`;g���a�1f����;��?�%�\r�u�(���O|�B͛4��8���%�f�a����?���A/�xI�bn���h`���u=G3��~h��L ��yw���o�ߟ�Z:i�3}��Zw��Z���C��H����\��v'�>�:�E4����I�I�Q�c��?�Yi�i6~4󺙪l&4T��d�'z�gl8                P�
m�%--M���6�b��6�f����Q-�R5F(   �G�1�ǯ*fD�e�o>�YU���_�t*u�����i?���PL���TDdp�>��������	h<��Q
1�Օ�ڹ���5��H��8RC�����=��ן�)�����?e/����m�&!#A����\rv�.{�2�y��GN���ﳱU���kj/���k��u���m{{��)�os��|Q}��є9S���SU2���RC8�Z�w��.��y7�;i��t��~�V�_iO{�1��_�f�7�n�u�9��5qkԢn��w���O
����Σ~����rۗZ�m�VŭRaщ�_��R}t�G��u}�k������ݯ�x]                 �9�N�1���L���� ���8�)**����`�^^^պ~D(   �G��l[�\V~�bSb��o�_�Z*u~o�^�J�굲���l=�U����]���B�l�����[A~AZ|��r#X�S�c_��|y{y��dh@h�����?i���Z�}�	��L�i���S����6^�u���E�b�?��ɚ3݆_�EΓ�1�?/��6&l��	���M	�l��X|z���>T����������;�^%f%�˞;!6S&�0���L���tUs_>��q��Ky>��&̜Pb�k�c���1�3���~zOw��=��m0��b�-�O���^o��F��3���;4w�\}��m;���e�7֬�g���/�WZN���O��z
���2���Ƽf�ӴU�                �Enn���������Ogee	�>>>
	9��T�b    ��"��:g"1�K�pO�o��^1��e�����Zӈ�e��s쓧�J�U漹�b���^��J�Ę���ݬU��t4��I�u��MT�k�O}��U���6��-Y1�߆b~-)+I��|�w-ݳ��e>Z���d�G?�mso;)H����U�]uR,�8���留�i����n����]<��3��y���8׆ON�y�n���	�?��]R$��c_=f�2�����[�\��HHOp��6�����ֲ�1��8�<��2���q��0A.*���u�Ѥ��y�?էy���|�F�Jz�                �6���QJJ�233���n�/�v U�Q�F6SK�T��   �QM�4)u�|��1��wƿS��g��PU+�96RsR�i���~�5��T�7(�	^�s�=�r]���������֒�N)9)�9c�++_��5o��;]n�&������)&(���66�R��X̷w|�-��~�z��7lx�ّϞ�m0�/�|�K�]��l�	��Xs&�9�H�	��8�F�1�R�ϙ�ʅo\Xj��D������q��Ӂ���̳��,��ۍ	ݺ���m"ۨw�ާ};L0��A����	             Ps���m�  ��\.��������94!�_a�N���E�B�    ��L�4���(_ۨ��q��oѿ������\��V7�n��i�i򴣙G˜�\�} 1��,{NTv~��w��p�<���j�A~A�)ȑ'��)fb1WO�Z1�����ݟ�=a�������CC:��0��@�;�]M�9��ǰ":5褹��*�7മg����q�/�?~ފ}+�:n�z6�q�;!�SOFb�%��He�gU���M�������*嶌�4�P             ��ٙ����U��G�z{����Bw p�),,Tvv�����& �p8�y�xAA����[�nB�    ��}K��-ȭ�u��J˺-+�b�(5'U�b�	Z�=o��s���ۧ��
t����	e=�FuŔ����`����J�����n�~�`�.��H��g֕�]�<g��:i��_�Q������2�q'�2��8�;�Άg*���͟<_aan-o"0�>�'����v�z{�I�A��u���%���&8�H��Σm謼�aѲ^K��d�e              ��6^��H7|x��)]urc����7�m� ��e"/&����f�9^<�i��읢�вeKEGGU�P    �
�*u.�0�R�uK�[�ǡ�����`-ۻL�ebω�j@���z��@�M������苇���fyBYϱ���N��D���/s��@���ˌ#*=/���˴��`�`5�h��T��)u�|�}�Ƿ�y���z�	s�.�p�FtQ�:��6�oТ�N����ɬ�g�]T;��7��fߤŷ/>����D]��eJ�I)�r��ɚ�i�j+�8^����<����������a��P��]X�o�P             ��жC�����q���j�W��9�XGӮ�fwg����  ��N��������p� �9n�3Ü&���l�?|�p���   �j�udk;΄�A/.Q��R�hU$xTg&�Rٙ�Sp_�3Oc����A��?��_��o�۾��V˼o/o}x���5���$�9����%O�@�;Lf����vd����������^���{u�2Q$��(���}L��"1             p���h-��P/�|Y��vgv�лYo;a��v �ʔ��ic/iiiv��ŧ�a^^��$�����&M�U�P    ��)�QDPD�s>©s9���G����=z;rr˜7{H�I�'��9o^�@yv'�.s>�/X�'L��W��p_rv����xϏ�
�ҡ�Cڑ���]��Zu�*��jW�u��5o�{K�q�)��6�?��[˚�͕�]i#1��{��=o��4k�~��Q���/}Z]v)u�H���             p2���{/�W�w�u\g�ǫ�u?w�s���  �f�����8)����N'��eiݺ��.T-B1    <*�YzD��xJ�&n��w��\��R�sl�P������9O(�X�e���k�O��_�Z�/�bL����ҷ����g?ߑ�Ш�G�XLi�bC�ѭ}oմU�*�~�Gi����qk���ަ��p���sl(�ϋ�l���L������̊}+             (۠փ�����i�M�rۗg|}f'qfg{#;�  U���P�����̴�)))6 �p8�qs�Y���ر�ƌ#ooo�j�   �Q)9)ju�$�!т�

��������CS6��s\����Z�����`��ɺC�ԽI�2�{|��6tr ��P1&2��qZ���(ώ�v�&_L�B�^e�h�D�p�BL;X�u?2�ui�ŭe_��͈�q�y��̹Eo�y[�8�yu̫�>�Dx             �=&���͟��/��R~a�Y��6�����qxc P���󕖖f�/���)>4������6����СCu�y����K�z�b    xԡ�C�ѤG�s�V��ĭѴU��^~\�q��Pu���.G�C�oV���t�'��]eϫn��c�\W�V�k��� {e�+z{\�!�ЀP�0�]3���>��Y��/ھH�Z�/�q�˼��S�2�]��n��C�ztأn-�:n����O'�_�*"sn�w�z6�Y�2�)�o�/             �{�{��^�i�GfNPlJl�]��A�c=��\�{�,��\ �[999ǣ/��3�����UݺuU�^��͛7W��x�    u �@�s-교����r}e��i���zP��b^Z�^\�b�˥d�(57�F���Yi]��<�}t�2�˻@1�p��s��F�ic�F���e�_4��@����2�����=~��en]�#�����˥��?��'�7�n(P���$9��             ��>�>��qY_��ע��=�N7ts�찫qxc}p��fH��nJؤ�3� p�1����;233���q����Pn.!1�L

���q<c�����    ��I�K��V�z��'y�j;�ٛ�W����R�3�~ѿ$�v��unعԹ��G��v(�����u���Z�|P�А�4q�D��H��^�MnRh@h�˚�����o�m�׆e�q��{�߱_�\�zMR��F�.׵qWM�3Eo�~S             �_�Z7K����y�L5kP�ru���ӛ>մU���pf��S1��0���a�]����뎹w(� [ ����!3RSSmƌ��$�����gb0��Ѫ_����GaL&00P�y�    ��\�|�&�ϊPLmVPX��G���$&��i���.un}�z�:�ѹn/?��x�yџ�'Tj��W��+���\��}l ��=��kԿ�*`��K�\;S�\�^�zp��n/�̈g4g���	             ��ow}�^S{��>��V�\��~��W�^���2w
�[f�{��/zl�cvۯ�d�e����ۈ �f*,,Tzz�233�aq��p��iii***�3���Waaa��/����8��G��3
   ���Z/��U�������
5ۺC�J�ti�E���ɑ�'��j���K���`�1#��h�����ӄ��ܒ����uM�k4��2��ۥӂ-���0��?�&Jb�h��gbb�ۻ�|th�&����V�$             ��L;����c=Vn̥G�����ݎ�4�h�Y7�*w�=��h�� @�s:���Ȱ�1s��<s���T������3L�Da�����\��b    x��r����gӞ%�_|��B��ݮ�ts��K�3d�q�f��)O����eΛ���w��jY�e�/wE�+ŜE�"�n����k���S�r�v��#��/K�h�Cn���o��@G��yt�/3��8B1             P�¢B=���~�����(�Q�ˆ����?�;]3;S�.�.q9�-�;�߱;�,ϴU�t��{��� ��rrr���i�/�!�1�8�����(<<܆_L ��_��0QQQ���P�P    �3_�/-�.���[{p�Ps}��k���҂㺎�X(�J�������(O�&�N�r�Z�S��:�q�Rn�����7VlJ��v�7���o��w����(1ӭq7m;���l;�M��|E��B���3�*�Bf���ޤ�����             (ْ�K��n�q�]r�%e.;��D�=����k�������s�?�{�c��*�ٹ�ߪ�7|, @�0!���Kq��trr���vU���Waaa�_�����m�DaL�N�:����B1    <�-���Ꮧ:?��dB15\rv�V�[��m�8o�4�<���R��vum�U�[�/u~��E� n	�,w��1������h5kh��q8��TV(���@)9)����6���Ou0��V�}���w��AuK]�¶�(����'�o2������~�
��1�z^�g�v'�����̣vc�^������D���ƞ7*4 ����D$             �a����=<�a=3�Rwitj�Ik�[����gw�ֲ^K;a��6�[�z�ĭф��ϱO ��QXX�����/���r8����4���@�

������@e    ��L�|A�|Q�$��L�S����@���O������}�Ӄ�?X���Ae� �Y� w�8Ky�{��_<|�oKzn�f���F�l��U�V�p݇��i�2�2u6I�Jҿ��[O]�T���s�=�2g����C���Ly��Y��w|�����ˠփl��D��������J_OV~���>��Gu��ο���9r             ����K���q����؝ߕ��Xl�5�4��(i3��`�,E�"=��9��7g�S  �9������L������L���H ��������m��`L�8%g�    ��~��^�z�s�~��������N���n���WLUDPD��w�K/�xI�)�Ur{�kt���q}��q�q�f�7ܱ|��r�11��~xM��U�t�'w�C�zv�z��W���Om��N�w�/-�F�J{�1��z�����v�V�>�8���u6i�Z�{O�Ğ����G>�[T�m0��?.�G�ˬطB              ���
��������xg�5�C�b@Bpw���-P �-Z(�B��o[�@q� ���S,��	�A������/���$�����z�Րyff�;�3�y淜��yj�m+�}E����h��-6��""���A0�"!0���ɿ���D�����C��#�0Q?K�D	�A1DDDDDd��ÐC4S軖銀#8zd�$�a���*�GG;G�o4��42�k�Ib��M&���V���;~ǻ��@d�������c(���fY��-@�ɕ�g���Σ���(��F��]w����`���j��2��ɫ'*�jh���m�W߂��2_��]�v��W�Hv\�k'��zy��p��5q���<L%D/�������m���
Q�<x� ug�E��=1��(����j>:�ja+�zzDD��˗/U��������S�"��d<%��0OOO5D��H ���#���b������,��|�������Su��`����Q|\qu�,��=cѳBO�pJ�s|��ѹTg�84ä���*ߣB�
����a֡Y �		Z�z��6��:����G|�wm�M,����0��X����cꁩ������2 I�j�i[��
�)��
�+�<G�k��5-:�����3���!��`ܞq���H��� |W�;�m�=���i""""""""""""""""""����Wuy �zv;kʬO+4�����6��5Q�s��%�;waaa*�����>����I���?������D��A1DDDDDd6$��K�.(�����Sd��kQkF-U�N�G>��c���6O��Uo� A���Eo�>���ͻ7 ���V �z�g,��]���q��m���Na�ٵ�\�3~���K�WÑGT`L�@�x��DƖ�\�VE[i����<�=������?�������$I�UsTE�2]Up�����[L�7	öKР���*���5�3d�D��Şt>Wir%��w
n�nѶ���|���n%&
�j�*�����⟳��'0��8"kŠ"""""2R��6�-Bz� �]R�mJg.��]����&{�<�NC�"-Uѿ.�ٯj�
f7��+{����yj#�?�6ک�+O�TQLI�햴S�0G;G�m���B8F��� ��)��`�����O�^�;�e(��f`t�ј~p���擛��L�#�����0���<4Ӫz;���M�6�[�/r{����������8}�4R�\5���J8�;�m���*,8� DDDDDDDDDDDDDDDDDD7yR����K
�)�R��w�v��5Q�q�����ꤓȜ��������0���eppp QbĠ"""""2+R��wM_Lj2I����{߬�K�/1��Ib�B�����_�	l�ý���Sg�����f����e&I�Da�m0V��*�C]WtQl��sF����Go;Y'���һ�W���
	��@$�i\�q�������W�^z!�X ���S�O����_@.�\�m�)�
�+�w>��sx�A�d�Эl7�(���S��凗�om?������cf���rQ�s�6�[Q�H�c��LFr��O#�E�,�岔C���94""k���c�����\\\T�K�ԩ����!���666 �O1(�����������U!��h������UQ���~Ŗ[T�x\I��_?�2 �Se�Fhx(�/h�-]���F�����#f}5�7T�\�ղ�G�?���yj�m�2�%�i����(.Jf*ip[�)�5eV�-����ϑP��=��>���>�4��9�`뀶�ۢM�6���&��5;.�%����|�9�h�����ȍ#���:,Y�T�T�Q��?��/�����=c���k$$yh�?ah���gCڗ�X7��Ŝ���7�Υ:�z�C�>G�����bY#�]Y�|9Cb�$�zG�H LTLԿ���@D1à"""""2K߭������]�
Y+`S�M�p�V�Z��g���ͣ*��Pn�n���*�篏�y�"�sj�����������l� �"������}y7޼{�w�pQ9{et,�M��h��D�@�y�j�!���.(��l���p��_oG��5���S$��g�b�?�UP׏�T�a�RV�Ad�s��\�����Ҭ9�FoP�A�8��J�T�U�_o�O��r�j����an?���&�ܴ��b��A�\5U�L������Act�9m	��"���b��軦/^�}""kr��qܸqD�?vvv�_�`>���'"��EDDDDDf���w踴#�x��ڣ��3U���w�8w�B�C����<{�L����'C�T��͌��\|]w�S��m1W��h���G��-����s;��s������=s�t��H�ܠ��f�a��� ��9�:S%3���f����Hh�4j�(	���E��`��F�+����y;��p��6��.����R=�������3��X{f-,�����~>w0� z���`��>�ĪG��������������������(f�o�)�S����Hǌ�@�@�k1����۾[�n����4��;�ADd��ƽ{��(1rrr�$�����C ���Z
"���ْ/���돣7�b��T�.o	�T{�I������髧 㐛E����2�qIm{�Ψ����J���m�c7���� �/6���z�(����`�+�`ߵ}�Q����;������fbjө��S%�+�e W��[�cىe#�Q������%���퓰E�Q1���G�0p�@��i6�\��B�4�h爰�a��������?��H'�ӚNC�"-�m{��5�X�B=�%�̪���{bT�Q��m-���!�W0z���f����]�z�=�5�����>��DQ�vtt���ٓ ��0����['A^Æs0h� �
�$_����d��h��a�,S֫��z��� 2������}A��WFޑy���+X��P|\q����|�}�cH^��X�?T�öC�� ����Gcs��q���N�a5��q��:��G໵����{0G�N�R��Ib��=_�z��mK�?""""""""""""""""""�^��E�3YQ����J���㗏?�N��w<�T�fI�Esz'{'Lo6�U@������sY���D����...`���?�xzz���Dd�CDDDDD���+�;�.|r�`��p��T��ˌ|��'�c��q�֭���hN#l�k�_U �)H�������F[��p��{����l#7C�S�?軦/,��G��e'��Юz��}2^�IV�]�c7���?a�ٵ0WGo���Gn�9���O5~B�B�T���.ܿ�n+�aǥ�Q!1�
4�W����vߵ} """"""""""""""""""��o���SU��>�!�<s+�0Z�3��K`n���������.�%3�D��8q���,Qhh(�̝��Ӈ�$FBa�~��y'Y��E���f5��\��tC�����)���/���׃x,K�/��gw@�+�tV�Y�&�MЭl7T�^Yg�AL�{��/m��}�����9�ʂ��[�����]�7�\كU�W��\{t�gׇoA_�o8���2�H�"X�a�
�賺_?ss���XO+A+����#j�@�`kc����o_�������-��X3���m^�y��SA ��!�W>���.Z&��DDZ�!��u��m����:y�b��:�-=�4Na��H���O:�=x� �w�Y.WGWLo:�7���?��18�E�#ȳ�=����z#�`��6�gn�y0� ""s���%4[[[���}���@D֍A1DDDDDd��T���=*e���D$a�D�pwr7x>�_>���'�M	m�}e7�?�o��<+xv]ޥsܑG`n~����!�˩ۧL��������Ր�5h��v�g-�E0��On`�3]}z5C(�L=0�+�G�d)5�Hqj� jN���W��Ҭ8���oCЯR�/�I�e)�C=�m����7����/&ȴ� ���e�c��p�9��l#Ƕ�+����s�D�ΞX�q=<�{�m7y�d<{�D�8��ȉU�����Q���!w�ݵ��G;G� ÓWOT��O��UЯr?����=��b��%��GJx*�b����+��K�x��)������������X��#{��Ѷ8��+���6%�8J��t4��	��ʦ�V�c�k8N=�ii'���%x��޾}��`gg�!0���j�KH��M�:d&"�Ơ"""""�h��"���65DI��RdB&�Lp�w�KR������wx��)"�D���Oo���{��Z�_ܮK���b��[Oo�  ����M���7*A
�^E�R��^f` %	��}��W}�F���QaR��s�F
L�G	���|.����x	�iV���}�Α��L
Mڣ�Gꆴ���Lk.�l�ֱ�)��/�a�5}0/d��{-��7uބ\����{���8'u���}��!amrL%""2TTI\��G�C3r^+Z�2�wZou~(C����%��߾��%���c���`�!߱X:	�Hf�̠�����^�'s}D�L�Ó ���Z�@����Z���X�O��E3E�tEP$}�N�[^�9]��"߃�v =�9��K;���~�y�DDDDDDDDDdy�o�em����Ao;y��ە�b��9�^V��W���B����m����B�-�tDD����� 2y�G�`$F�_�a������%3�"J�CDDDDDVG^��ĭ �#��ʃ�2���{�·�/Je*����l�5�װȰ!7g��+��>�ѯR?���~2>�Cr5�S�N�q0]���%R�����O�_%�8	M
��6�
Y+h��t~:/�B�,�����E����7+�Qa1�B��Ս2/)J��=9��ܽs8|�0v_ލ;��(J���0����K�;#ǡ�On�ԝS�������?ypS�3�嬆J�+��%	T5��z$�P��=��W��b�e'�a⾉8}�4,�Q��j�Am�$�o�p��5ė?���e��V>�TCS��sy�evaLr\��9.��}B}y��Q��T)�y�x�D����J"U2�}���T�Z�H����
$�Y�n��F���t�T����WCkU��KT����'ADDDDDDDDD��@�ц��3�_|��w��yy�w��M�m�o1��hա��<r߷�����1~�xY[[[���~
�����b���������L�H��#�W��ފEZ״��mjͨ�#7���~��DЩ �m1yR���MF��h�n�v[�-���b#�w�"��#�D��ma��Fg)`�n�w�<+A�x�J���]63��\U�D�'�{�:/�H1��u�P�!,:�H�����u""�x"��;z��F�<������^��������ͻ7H��|��wcU�ml��u��ѥt�B�u�q��X3镩U�V�uۯ�<y�y�� "�u\J�^�k��S����ٌ��b˅-}n\���`ݨ@2�gBb&A/5s�D��T/���.�s�=��������GWADDDDDDDDD�/�H�z��؝�IG���Ò�K��#�f;���k�_CDD����C��#�0Q?�3*DD�Ơ""""""""���Z���NTq�>����vԝYW��TQtlQ��5}*��hR*S)�3v�X�<�������c?m\��ǟ��T�8k�~q;:.���PX�t������/ڶ����	��fU�̥�0�g8���ڞk�>�9������\sȦ!�A��V�_.k9���|L��M���v��賦��k�_�?ނb�=����	�mT��$W��hF�C��Zn�!F��Bu	rPe Zk��L%�|AB��[�
M""""""""""�$��=W���C3M��.���b��;Eu�@DDd�>�I�:5<<<T ���q:n "�	����*�(�ހ�(n�n��y�Ϯ�]�w�Rɍc�M8�T洘��;;����޾躢+�^�o����+�ӦvN���5eVus�'��f����u�cʁ)_(��=�
L��s��V�^�Wo_�N
������+ꇦ��⃋ ""2�L�0��<�,�����0�!��$a��TNW�}�w���I���~��˒�}"�>E��ή;1n�8u}���[�iJW��L})�gn�:0ޖ��>���h��*��Z������������ٻg�<�9N�9m�e={�L�ߕg*'7�l�2���b���...*F�_���?��xzz���DD�A1DDDDDDDD&"���9�3�wZ���b��m�d���C�1�1��t-�Ug�l��aK�-8��k����&]e2�I�icB�tzU��>���?v~�p��X��)2cG�j�0T�T�A�`ڂ8��|���K�5�����:�T�V�]����;�:�ӲNL�ſ����a$`�^�z "�$I����<s�M��RbӹTg��yX�����g��.Ȉx]��������%�N�""������!�E	��P�����/��`P����E��p�9��&������G����_�n�rYz�~q;f4���sti]�5j穭�b��)U�^9N�� S~.���W�2�l#��k~��#"�E�T�Qo޽��wҋ�lCQ���ث�y����]6������������I�\�	ep��]T8���T��\k�9��ȗ*��%�Һ��wodI���yv(�A�"8v�XX��[�5�����&[F�B͐�.)�Ⱥ��[�Z�C�-���/޼���'�yý���w3r�J�,�
�-��$�m�ѯ�.?���������������̗�?�z��<�`����s(�W)�^�w�,�DDD�bkkWWW�"0�
�*U*$M�g7��z0(���������D^EF߃��6��v]�����VYH���r���b��(����6�=0��|4/��v4I���V�^)���k,����:c��6��P�6H��E�v��Q�5�{x�$F���P�s�Θ�h��4�=fd��iH��>��R �GN��\�\��	�Y�z�
�1e�5Y������Ѷ��O��T�K����%�A�Ϛ2+�Z��j�����揝������aI޽��M�^݋�W����c5�}�s[߂�h_���9���S�?Xwv.>�k��95|r�`���&[��cQ�	���f����I��ʾ2�W>JW����W��R���N���k���vb��]j�^{���v ���|o������[��տADDDDDDDDD�G�'6hn�����^�z���'7��� ""2���\\\>	�I�:5<==���%�!"""""""2��U8�j���߼}��K�Ú{�����O,����!5��0
]���SߝRa1kϮ5�khX��*�v%ڡ���0�,)� �e�*��G
y$T���[�VR��2Jv�_��B�$I4۞�sd�'��ĺP�`ڂ�Q��*p����)����펿��DDDb�х���f��+���U�f����Vo۪9��cɎ� �9���a�$tGMV�^���ǿ�x������&�p�\�4�;�9��Z?�傖�To޽Q�%�<s}1ο��ɂb��ʆrY��w��iHS DdZ�^�sp��h�+�Ku��*~���_���(�=�����QF���/�+�`V�,���$�w婕j���f���U��|�7�w

�)dp���6f��~��$�H �Â�����ȁ�&[x6��H��H�DD����I�D#�0Q?�{���(�`P��09�{K��#�� �g���hV���6m��Q���uV=�Z+�ۆm��a1��<� OgO�n���O���W��ĕ��W�_��ӾD{���UXkm��ń����E�M������E�M�R�1��T�0�(���ŏ��O��Ӥ}����b��̭����1��4�{����,ˑGT(Ʉ,���R�wK����Z#�C��޾���[�ޗ�w�F����q � vtݡBM�4-�}]����۰T�.��>?����������}��E�u>����s�à"�p0������V���W�m�d)ѹtg��5?�?���`d������O�X�9�	�m�o�~q{��SZzb��mx{����Q��ךx7���ADDDDDDDDD��ĭ0W�����*�_j�����<_x�hW[WY:[[[�����	���P888����cPUR��������k����ňv%ک����Uo��l��M(�g�h�B�ȭ�R~[�[T�^E�JPE\H��Zˊ	)���O��#N�I�B�����G
���o�=W� 1Zc(��m���ۧr=���:����@���K�]Z״h\��*:'""���������8�� 2�Ȭ����-��Ĝ�s`�$��TB�CQ}Zu��wJ� �bgc_o_L�7�j��^s��N�N�o3���_�_��W�Z��7 "�"�W�Z{�ك�95�IH�bL�U�+캼�C0��]����������6���⃋�3����o�9�i��T��b���������(F$��ڸwGDdjvv,�7���Ӈ ��`�g�h�&""�xD""""""""2!	E����+G۶n޺��u�Ϯ�{�����zz��Tƴ��жx[�v���ǡ^�0h� ��{<����/+�sjLh4�ҽlwU����XM_){%�o9��3�m'�g�4TE��N��'5��.���~������(��G���
��؛A1DDd<w��A㹍���~8�9j��+�g�A1�v��U��:���]�M՜U-:(F��}���|��_��@c�?V�$p$ %2� Y9.uY�;���lS0mAbv��]�q=�*S������uδ���X}�f��wN��u߫���T�Y�N�x��1����������������#lll���{���`�wwwxyy���C�#""�aP��uZ�	�{F
�Ѷ-��$Bz�������_k���k�[�'o��Ⱥ#akc����m85rՀ�"��7x�X�f<�=���a����Q�R������I���C1��Ϳ5���{���X;	�Y�UrV�5;x66�� J8�_���Y*4IK�UADDdL�n���ѳ|O�6��U���+��z
����f�ڿ� ?]
�) K'-��b$�3�[�xr�h�j]�����|r;/�dP��P���vj^��w �2��+ū�/����;��z#�W^���{/9֮;�DDDDDDDDDDDD�D���������ogg��)S~�����-�0��� "����""""""""����bmǵHf�,���3bO�=賦��k���?q��i,n�Xo�N��u�+X��,�G���~���"�-�kZl�էU7�wp)Xh���m'�=�2#��0Y���l��X�z)һ�7���K;���o@	oҾIz�b<�{ K�,�������e��Q���b"��3W�;#b�����ЙSd��[vb�j���%����W�#w�4�r$��y��:�-:��޿Y��g��=͖2����]�_k��٦P�B�!"""""""""""��%K?~�����CLT ��a0�CDD�A1DDDDDDDD�@�U�̬�mW U�TѶ����M&�M	�x��l˅-(5��tX�<��h���z@�%���r�v.I]���"��W�R M��ug�ŕ�W4����.H��%��~�6�mt:�Nz��_�?~��Ytb͙5h��^�}Jxg���Uh���9M#7�X=�W>dI�E2�;��5�+""#�.w��������p����	M^��7E����\]�kvst��W��������w-��������9>L[P�3���N�Nx��9n>��sw��`�A�7�+9FNW���G:�tpN��K/޼@hx(��9�������0'�Z��z#{��*`K�o���e�Ku,���?8v�Z�̙l�r���ΞH�o߽Ž��p��URq���/W���B�4���%-�9$S���վ�ԝS�/Y/��8���Jj�)��0�b�H�.��bd�#�s�G�D��pU��[���q���6ZPL�<�5��Y s��3�:�ʚ*+R;�V��$����S=x�@c��;���ΛM�eT0�O$�P�%���r"��ze���X��U�Aʬ�;j[{����|��K���<��i�B����"Y
Y������aPY�ܹs[TP���-���>�HLT� ""�à"""""""�x���nW�zR�w�hQ�*e����:�kv��E��X�;�G�L�4�IA���K���?��U/��BA��+��_�
	����mUO�k��Z��t}$B��Cq���m1e2�1x����ۊn,�43�!븖n��<)X.��,�樊��+���J�l�]܆U�Waىe*X#������E�����-�}��޾��N�������ͱ�H�~���'A/���s\����u�Q+O-N����켴�LÚ�k��O'�$6hV��o�*9���k}��|�����:~'	�}��7>�}T@�!��ץ]Xxt!V�Za�0	=�_���qR�?~�x�㤈�[�nhT��:�3x�`���/~߽lwdJ�I�4c����gw����;�o��
}�
Y+�(;}�4�G{������`��:۝�u��-��eK�]Jw�?b�p��쾲[oPL&�L�G������s�l��l����m)�����~=�]�3(F�%$L����?�%�3��1���HHr\���:����f���r�2h����c�ŭ*�F�>b]�s��{�PP	��GΡv]ޅ�!�x,P��\��H�{��~��6�K���s���7�ux�?[x���$�N{ÂQ�\ȵ�.r}!��&�4�9N��~ݦ:B�G�X�� W""""""""""""k�'O�sagg�O�`��ԩS#U�T���Y�ţk�����қ����Pv}l:�	�LS�O��mW��9-R�;��@U����/��h�U`p��������)�tX��#跶�*��7��P�T�'��>�_����{�N�C�~�7F뿐B]@���/���0]��'S���P#W�h�=��p���al���w���B5L%�Cr��Vbj�9;;�PLR-A,R<;x6�N�h^)��Ā*t�;z��A1�i�1�w�
�1��%�D)���{��AB�B��M&"�gn����K�Ed�~q;z�ꉳw�">�qC��~��#
�+��e�����F>�W��j�b~)��Z�d�yP���'F���d]6�փ	�P:si���8�q��� t+�M�=��4���S�WL��9	����w:�IhTb��^�;ސ���V�!��7`I�\˘S�Flm8�Am�~�9�_�5(F�$�D	�H(r��c���y����O��2$ `Ķ*�L�LM��6����<�w�<@9'뵪�΀��$糝Ku��U�GF��1�^��$DN�S�Oa��*��������S�	R�k	]$�)>�bU���=<dY$|�髧����=�5�{�>>>X�xq�.���I��D#�0Q?G��2Y�Q�5��v��� 2Dhx(�>]Q��Ɍ�5
�޾R=*K���nSE������QV}��"F}j婅ýc����]�w�
�E��h�1�Ǡh��h��A�Ӝ�w>�}�8���'7���,(�� 2��פ�p�wT��rVӜ.��G���Wdn)��[�o�V�H���>?�cɎh���]�g�eH���fӑ9Ef��[�X��\�y1��	)$]t�·d{��m'���?�e���J!�c�A���t\�OG���+�Ŭ�Y0�\��0��tT�^�(�K�OD�bm�:��*�O���������#F�%A�Z�r�²6�P!k�X/w����p��_|N�%䘿�������:��"AQ�������.�	��"!��@��_��>ײHKX? NǬf�����y.:�	A�If4�����A�Y-СDt\�W]���(�B�WI�_leM�U|ʱ�ۊn�|��V1[E�w�$�N	�j���V���ў���Ix�>�_>����*��Y7%HƔ�M��`�ܵ4�'d�Ş�P_	�!"""""""""""�Vy��A���b�y�������C���sԿe<Q�����(ƶ]�""��ӷO�p�㳤̂�i�GP��L
7[.h�
ݺ�骷��,?���)\Vs�AmC���ά:*(1�B�Ca�� Zm����9u���$�O�w|ě�8Ϳ|��&	���L����v¼�yF���Oh4�6��T#j����4ʼ$�E�%�����0�����y��F����#f~5S����8���$T`N�9&	�(��$�<��ͱ��ćv%ک@�,b*.�>r^���dK�-N˕���#�U��ζJv0iPL�����9��q�g�e���H�Ǘجs�?���RNs��k�a-d���5�����V�ӎK;p��-�7	�Z�ne���Q%G��A��M���N�Ͽ�����F��L�ӻ�G㹍վ>>�kTu�:���"ck����B�Y�T)ş�r��!}����#�䟓�ү�~��ɖ/A�����'7M�� Ӓk$WGW��#��Y��u���������������C L�������]]]�vo������$"""""""�g�o�1�m���,)������H�$$Gzz������= ��>x��+	�^s8W�����q��q�������ǰ(0��l^��آ8�Ϸ�/&6�h�"��"]�
����ʾ�o���7�ckL�1F����Paf?o�٨����wUo�Io��;�cM�5h0����b�歋��f�:,)	b�>�L�;o�UH��|��qh�fPL��Ց�=���$�F��K�9D
�z��W���*��һ��oM����҃K���eЃ\��v_)� ��	��o��Z�q��%5�2d����&�����ͷw��Yo$��V�Z���բV059�Ȳ�ok��HP��n;Qir%�
'�v>�}4��yﱛ�`N]��}t��J��)�bd�Z�:,�%[2��z�{/?�""""""""""]�\������߿���ŉȢȳ^�k�F�p��!���!22�`>���"""c`PQ<�p~��z7G7���䭃#}�����~q;�~���9�3���k �'uf�I��R<;��T�Q5ڶ��M(A��;un���>�k���zq����s�_>V�4�����]��PT�FG��f~5�S1gZ״j�6$$�ڣk8q��<���+	y�����5�+<�=�7u^U|��!9�K���W��4ǟ�sZ�G�_�����"Y
�Q M�P,ڠ��[�����e8LE�ѳ|O�� 58,X}��7�G���$�D�ȓ:O��Vs��$��䵎�?ڠ���=���P<�x�g��� �Je*��)2�^BV�[������0���F����{~O}&��q0Els�Z��9�����P�ܣ�Gj��3���A�re����~��R����vޮD;���t��T���Y����ET��ϱ�J��?���9���[X}f5���KHh���?׸@cu�}��E���_�_�~L�t:�I�ͫگ2($F�1��V�(�(�wM��)3�dƒ��C����,G���T0f\�����ǋ.����'7�k�c����^:Si�Ǥ�EZ�P�!���r�ihH���#��%45U�T�)�C���Ҹ���ΛQ|\q5=����7�n�9^�s;&-8�@���G��|�t�M�*�dD�%!B�(�j䪡w��GADDDDDDDDD	C�.��<�窮��d�Ȯ�3�}n�G��\xp�Ba�ŭ����b��X���g.�~��`gY��3����(>1(��������(�I��;����'ڶYSfŶ��aىe農�*�Nl���ۊn*,Ư�,�0֞Q[������)�~����<�#��o;~����R�`ڂzۘ��PBJd���^Ut&�[ё��f��u/�W>�vN�N������x��]�^��~P�Z�Pt⾉�{x..ܿ`�<�!�9����
4R�ȶd
2_	������~x�хj{<{����r����w�Z��ސ�!Շ`ۅm�wm�M���7����}��1v�X�xrCsz)����hZ��fy�jz��*�%�qX�^���m8Voy�%dN֝=����-��B�2�ЩT'��@�$,�ȟELR�<��d�$u���R����b�=�_���"?/�N��U�~l�)�Fm'���H���m��p^��"鋨�Z�j_L?���A1�}���e�/�A:c�@�����s*D 1��}$�b�?�|���G��Ŷk���&��	r��ػ�
U�)�b�:t*�_?G|���em�E8'�*r��������l#���12�[�y����6K�1&.׮��Scn�ц��9�#�����yH([�h��ɸ_k����7�TT����6%ｄ�I؍�"�E��e1�� ��[Ws~YRf���3�7MH�6�S�u��󛛫���sp�}}���Lr'��
<q�N�>�<_�Js�뷯�FDDDDDDDDD1#���[��}�3Z��|^��h��!���Ig9�L¬C����+��cPQ�w�*��N�mP�f���p�����bFc$�;�{�-ngg4�� �(4<զVÝgw���\O����c�H��H����W�h� ����eY�0y�dT	1u��}L�?SLQ&��F2�d:�M_����UQ��J��������ƪ;&d�'�22L�{�
��^z�ؼ�xQ��(���a�?���^
O��V;/o�\��\
�紘��
� c����å��;�'o��vz)�m6��x7��su�7G7Lk:�g֎�k��g��B�ےζ_��n3h�Ҿ늮j���Gʞ*;~��z�2�z��+�
���|����S����_�#�t�lb�ly��s;/�D�U=p����@_
�eеܥǗb\�q�3���W�Q�.n����۾�v��	$v��W�;���+���p��F��/-�����_�6r��Bv]�P�Ӡ9���S�Gc:b��`1?d>�	�&� ?��T�7Lj<	m���l+�79�o��bkB�	*�O��&�qiG,9�$�yIP٠�0/dV�]�z�"!:r^k
����L}֝]�Ν�Z1:d(a�{g�U�h#=�R+O-u^j�A%�@�ee�jQX{���]s$۱VP�|O5p��Xgj��}��,���$�R��pɾ�����������ܧ��bry��yR�Q�wU��O�N`HODDDDd�CDDDDDDD� ^F�T��{V=t����[�W��7Ɔs��H!w��0�2�g��i8�!�?���F
1��+�o�ك�.R?��t�����Ǡj���Yyje��s��=4e�<{�,��Xd^{����n;5kV�
�c��K��5TX�.���L�QAq%�-#w�T���W�1}��Ja���\��|�B�)U���~��Y��-�-���'���AB�*O��Y�����y�fh�a˰���X��IM&���]s��c��yigDDF�x��SqRE���2���曲ߨ���0i����d�;�.v_����&@��e˺��Z��C�+ￄ�u/�]�4Jv0jP�j�L�� ��L�y2�g��&�F��Y�� 5-���F�T�4��>��F0R�+(�z��H�V�J�t�ys_y�]�vz�H��=�z�h��vq[�zzK�3ii^��:��qib�L�2hV���x�.�k���h��f�)�p���%&�(�r�s����U��.r�9|�p��:"V!��WqrEl�Y�����`ىej0"YW�d��Q�G��I-��JP]l��⃄��o8^�*���n���h��U�L%5��b��:�_tAXs���o=�w���cJ�'^�j���%��ɳ;DDDDDd�CDDDDDDD�@.?���j`s��H�,���I���;�W=�\?{��Ab���t��`�rx���['�Xdpˀ!5���lb�5��K�mE7�y]4��̪�͂#q��o��Iz':}�4jϬ�=�������=s�\�r����1��@j�e�QBb>&�[.l��H�f�-c�⃋�-��z�*��Ez���	O3������̺1�����Nt^�Y����g��c���7�t:���U�x��Qgf����'N��������s�MH�1��;>�!1�H؁VPLc��H�,�
q2�%:h�[{fm����?�/����i
�,�N����a�y�C����Nױ�cv&�,W^���Єq�}&���[`잱�G���]��k�ΰ�����q���ޱ����T@I���4��\�g��a>�_�\'�4$&����ձQ��brS=+���[�����a\HЛg�{�<�J�]�tŘ�c@��}�9�+�9$�KRu��}�|S?_}dN�9�i�_�=֝]s%�%�ϭG�&:��vm̠}�		���)�,-��D���5���ɜ�"""""""""kӶx[�l6Ө�����Ʃ~�T��<������L�A1DDDDDDDD	�ȍ#�:�*�tXcP��Ǥ����wc����a�8s��]��4{e7w�޾Xqr��\�6ߔ�F3B����۠o㵐�#��6=����n�?�q���8/�!1Q$�D�����E��c��5��8)ƶ4��ga�ٵq�����w��v�H�����qhLa��8y�d��1?d>�k ߂�:Ǘ�XB-컶/F����O���5�5$&���H̎�;`����_�
}��5I�Ȉ�#$$����跶�Q�)Ao�a�:��X�W��M��r$ģi����e�L�zW�*9��m#Eɉ�bu��Ȗ*�����J�e� $s%C�mP������f��G� �NWX�i����2��J�]Q5GU�s 9>���?M~��YCs��3k�/�p������g���:��������?eY�n�����_���9^�����Iϫ-E���`J��jځi0w�#�ﾲ�Q�%4V�4_�Ѹ�R������m���r-CDDDDDDDDDѫ��f}5˨!1Q��@����aؖax��-������|0(��������(�IAx�qű�o�ނ>-�7D����cUL�?�L�V,Uݼu��.)^�}kU*S)l�	�N�1�V��z�L�E���;�7F��>J
鿮?,�;�P�7R����9��x~^�^:���3�+������`�>w,�Q���C�&	����ю��@�|��>\���:ƨ^��d��kU/�x��"a-*��8���^����;�t��i��=�MB�,�b��d=�#d=6FPL�"-��>��q7����[�XI�ר���m7��LP���6ÎK;�XH�����"鋨�CB9%TF�'J�U|iW����6��WO㼜篟c�����|�f�?��پD{��#�E�c�1����{����d=�0<]�5Ϫ�Fn��2zU�쩲1.kʬ���v]�2�7��`���m�
"��oP�()���b��5�� K�/��rj殩
	t��]	$#�!���Z̃���f9w��JDDDDDDDD?��ׅ~M��|/�C�P m4hn�ϽY���/�����V��*��*R����^E������7��A�f9=r�J�*�TRl%E��C��Z
;�>��ܷ���ܜ���e}�
X���M`�)��v�v�*�G��ҙK�N�:����A��Y��n��%��m��,
ϓ:�z����{�/y��:�����&후;��e^RD����1���^�%`*s���1��:B��凗1;x6���s��C]�w5xy�K������&)��k�ΠQ?}��H@���7	R9|��I���b���O�$u�b�M_Go��2:��9n���0����p��*�+:F��տA�#�פ��0��T��{���s��2)�R|1ο��
W�G��P1]�Z-��úr͡E�ӌy="��[��
�ŷ�/���n�C�Ӵ`S���.��{�a��}����bm��0�v��i�����zz˨˓mw잱��Xw`Y�|�c"�%er�v��]X�&��X��e��/�=cŴ*�Js�ʵY9'�����x�����������(~�Q�����{,�1��g�U�����e(�3�^��N�4��ب�Q�1(���������L�MX�����X�j�f;)���
~��޾��bH�!���쯳�T�EGY���6am>�[
U�7��s��M��X�i]N�`ǣ��m�d車bbc��1��o",����uňi
�������I���/a#�bѱEF��l�i0F�>\�iF$�5cy����iR��#� e����˻��������9^�LA4�>���)�~1�\�rjۗ���@t�ɕH�B�l�R�x,]Jw�9�C�8�����TR�8	4����"�C���婃N�:�����{$ae{����7*�hىe�<+Q=�)�	�w���%����?��LK�B�t���4r�/��F�4�����;bJ�%����G���膲Y�b祝��+�W>����'�!���=�6O9�j���zߘ�;�k̿����>W=Wu�iH8�G2�M�W��]|�DB���b|r�������z�r$�ZdD��A����z��X�C]s����ʋ6���m#�bM;0���f�]ґR���u���}}j䪁-]����F"""""JX�]YCDDDDDDDd�v_٭�Ȥx^)�\m������1
2�T�=sï�,]�h]�5��k'���0L칲�!1�@�fa
��"�wM_����9塚��_��.��Y�'z��Kp��9��}ʨ����*���t����Q�7�۠B=�i�~��dtϨs���Ŕ�X)���9N^��[a*��t�H�A�t�p0��Q����*DDF ������j�.cơ�A1~E��om?�z�*V�-��Xr�m��
���6�-R%O��/g/����h#�����Aq#a1峖W��4��5Z�%�s5	-е�˾�R�Jz�N�_�]�w�Ɠ�/UsV�'�.�fl2ϑ�F�)Q�)GU��b*e��9N�*�GL�9��S+5��!�Z��<���P�B��pu�&�����ʏd���؜�5�}+�U�IC6��gwa	�����+Ȗ*���8�U��0iߤXϿ��c�.������������5� �5@ ��`c!Bd!hwwwwwww��=w�����������٧��p������nu�����L��#�\����
�C�9et�і�S�ɻ&�譣      @����G��ͨ�7OKPH�쾰��r^>(���L~^����g~�r�]����2�=�v���   DA1      >�ܭs���V)�����
�)`~x]r����w��gF�,���5pDW���j}e
o=�%QQ���䃊Hろ%F���~�@��E���?0�"��Y�Kڄi�Z֦S���o;l�V��l;��/
�����Z��q��u�M�4�FG�r���P%{˶�G������S��оD{�m��-(f�i{�㮝�w�;��U[�l��vH�tE^i�0�FɄ�^n��X�!*ds���
Y*xt��vN�o�|#�W��ɥoݾ�0Ci5��_��j��u��	m���*���e.�M�g"��kH�8�/�~�tz���T��m�;g�R�sz�Zw�����h(��9��'�y�QP�^G�w��s�\\*X��/�&��Ň�������L0�#z܋HPL�bm,�4`��3c�A��e���$�疮S�
      ��7f\iZ��e�ѫG�ʠ*nfp��Uyk�[淭�M�¬MWTV��Jj�a~'   ��      � -v��NG��IG'�~�)P�QA��w˾+u�ԕ�"c�2�� SpU$��@�o`�+�QGtqOL�~Ϟ?�!��ЍCM0��iQf�TyMA{���$0V��4Ò.Q:�6-�sǊc+,۴@wT�Q�X��%������
k4���u~�e[�$�%~��r��][���p��9�K�ϥeN[ز��������"���xCd�W�}zwDâ�S?_}ss����&���2B�L�b�MN�7�:# �$��X��Of�E%3�4Ǯ��Kg*-���$�U����KT�,4AC����0�K���x��=��{�D&g�#O'���ny�?u~����9+�蟄�����}�݃b^�# Z�$��P��K&�S�b鋙�Ύ��������~�6v�Xˠoʞ<�)(pW��i�Z�j���6V��4qQ�Ef?�r���R��      9j�i��v�ᓇ�ttS�Bb�N�)�k�j���J�TydM�5Rmp��b�	   �     ��Fn)�V�ԭ��LI2Iߺ}�:?ȆS��SwO��/��ґ�	�E���EZʂ��(,�J��5��E�R'Oˢdg�_���b[���Ѣ��|퉵^	�ɐ8��2YZ��+E.����h،;��Ro������<�
53��v����B�>������r��>g����?}�T�]�'�����s�s��:��y���+�œ�ܽbٖ6aZ[֡!�^'O������M�DÍ^V%{ɒ4��7�u,�ѲMC+<y �_7�ߔO�~"m�K�֝\����֩T'�\����@�����R)�gy9~�DeV�	��$27�N�9镶6��8\֬�����;Y�|�#E�v�CQ\]��gگ
}�t�R�l��1^V�x�8n�/+^�xN�]>$�t9��e�]�yv����kJ���>Qzs�~��;���z�4�����-��$�j���¼L�)�������r�{�@�vv���i_w��s�`�����O���eυ=       �T�i}_�w˾��<��V����Z�H�j��������VK�AU���#    r     ��tt�6�ۘScDw�+�qVt����f��{gȌ=3�j���a�ĉG���M˩�d����/��R�a�o$�s�vX$�*��sݟ����Z����jJ�`y����ש�0�Wx_�f�jy���~���o�Z�jan_�,���c��ܭs���BYvd�	��"Voy����|�#˾~�	.K�0��v-`�#(������w�:�F�s-�<��+"����hȁ���۲�{�����^��p��m�(�E�ۗh/_.����i����f%ds�����5l�0黼�\�sQ1z� �_W�*?����X����=���8��	努��&�)�敠�ҙJK���Y4t&2�<V@,�vO���|�i��#�o� ��X�k������\�r^�^��y��Ǖ?6����,d6Y�d{���,�F� �(�7w8����l1R���.Ǯ_6v�X��<ޠ� ��o�sɴ�����<y�D��in�a      D��K;�������umY��?�ga�ua��h>��1��{M�5R}Hu�{q�    �<�      ���6H��-d|��N���B������'s?�_V�"�NQ�u]fF��t�y����Z��u�T0�Ì�^ֺ�����D��o�ЍCÜOtS�O!���lɲ9-vUoK��M"�G56�b��'U�t�-����}}͉5ft�>�����t����%�6�Ҡ�Yvt����*�Eo�d���X�hȊ]��[n�p-�u$�����: ����xKx���o��0��=l�0�A1J�b����s��o�Om=�Uv��%�;=6�9�F��.SvO���o
쥣v��՜�F�e�Oj��{�ߓ�V�&Q�UhB�\�$E`��	�j[���e\�sIZ,�)�s��{W=��ºtۜ�$�*0���{��nײ�O����Ů�<���7�}��5d�����jC������WM�5I~����k}���h�J�ߊ�+�M�G㶏�.��m5֜������s��       �K}ț:��6�=�ڽk��oʮ)r��y��i���4����]�   D2�b      |ش�ӤFh32���]1��<�sݟ��4�bN�9� )��P���ሆ���J�eZ8�ӊ��W�^榃��b"+�h�G�����ݫ�s^O�����H�U�H��On9_�|���7��.S���t{-�����/}i�v��	��!q��~f֟Z/#��47�h!�'iP�'9���<�����'���a{X�!Y�d�bǈm�r"3��uGbH��Seυ=R M�W�2&�(5r֐E���=�v(���=ds�Dڇ+�JC�4 �Lnʍ{7�쭳���>�wi�<~�X�yZ���\=�Z�Y��\?У�b�6q�D��	���5�����0�慛[.�S!zVc:m���s�Ȱ�����o��s��=�'�b��#Y|>��s�ǫޝ���O��i9R%{y#�2��|�U����B	��]�	�	�iS��e����yZ���o:��`iZ����>����F      �4�E��Yqt�G֩�UTUu^dy���Ŭ�Zj�iD   �y�      ����WK�~��*�J�r�%i��.?VG	Yvd���6����;�N�:f��$q���B�_�e�)��uկ���,�#3�͔�R�R3gMɜ4�ˏ�"q���M	����]�W�l"C�qZ,ֹtgYr���:ʶ��~��o0���q�봮���v���O�#*�B�{�����G�?d���������	�qR�'f[�a7VA1a=���'D{>g��oy��A��oئa���v�ֱdG��b�d�b��vL����ؖr��9��k�_� _��������)�E����}��Y�&�-���A1�`6f��la�~y2�+���81���m{�P��)vń�������D��z/�-+ޱ���V��O�(���*(F�>���K�m���*�ʲ��F��Ǻ?J�R����oU?�y��      �;��WP[�z.�E>��,�DR�p8���(x�	��vv�    �,�b      ���GwMȆc����P)k%	���q:r��;e��=>7f\���&'z���=���'�3��3{ȥ;��W�r�L�s�s�ˡ�eƞ2r�H�xj��?ݸCZ�ma�I���b9߀Fd��Ur�����R�J2��@��Z5dér��A9}㴜�y�l�7=}d�+�$��'�;�O�q���;��44�jD'W�����<��H�o.v{��x����q�������za�ÿhA��j�e������L�=Mn=�%�7h �8Z���Z$*�(3p�P2cIə"��kh�#�/���ͯa��<y��>�^oZ�31�o��m�����=��<��Zyl�쾰[
�)�]���$L#n__5g���pr�7�kP����|�򖁲zM6u�T�o�Y��|R����2R>��|       ��l�+�W<��]�wIŁei���.Q:��� x˺.���js�   �a�      ��Ї�2x�`3%��܌Z�?u~��c�{�ߓ������eѡE���9p逜�yZ|A�<u����%iy�i�m��5̈���B���`�7U^)�����UK*d��(�e���̌4�#�����}Fwɞ<�T�Q��<z��x���#"�Ĉ#ÛwZ0�E�Z�=l�0�qn�<y�$\�J'�x�ބ�cF�nQ���.�Z�f.�P*�Y���TZޝ�n���#��œ�N`�fW��������<�ｂ�i�֔]S�]�v��iX@�bm�5X>^?�oxӲ=ds� �r���rf���X�a���4�QFԜ}s����Ge����V�&���s�X���Cz�T�J�X�~��^ga-���$g�w��'��Y~t�eP�~6�e.��!)����vɷ�k�ƕ��ϊW	��M���;�GC;M�$ϟ?       ��(�����Vq�2��	�ɐ8��yt/�:Ցu'�	    � (     �O]�{�(;�yA��g(n�4tF�btTk��޻j�y��e9{�칰����J�*I�j�����?Z���J�ҝ��eߛb-O�jQd���LH���20��R�OaF~�I��]Z$�)���(F��c[ȾO�Y�&T'O�`~��\:X�&�jٮ#5�D��:'� �=��a����8�L������	ܩ���)(���2�Kˣ'�L��]�*���5����C�8	-��zZ��L�&1���6s�:���4(�e����kұ��j�i����A1$�#y9t�DUzL�~x�R�^i��s�ϙP��i�}��q���V��îݻ�u'���i����ϑ΂d�ƈk�J��������<��)��]fAԵ���G�X���TƧ�b��\Y���W�|V�<�c�x=&j����{'D�i���7J�h�,����V�Z�      �=}d٦��u_�����ʛ�p��]jq��Rx}Yvd�    �A1      ~l���ҧz�������yS�5�����К��h�PP� �G���aM\&��d
p]��L�9�֑_����	�	Ͼ�9��x�ޥaR��XF�m9��D����p7�-��e��k����N��ݡ��M�+�3��ґ�*d� ��V2Z��3�^��V��l8����tO�8Y�vמc�'���ǋϲ=���1<s�̲��N���cҁK$O�<��i��m=���c�
���������x��+����N�:J�(5p��v_����c4�I�8�����N۝��#*Q�DNۯ�w�m�Ρ^�76{*L-��W9;�k g��1L�"��ˡ���[�(�K^�2&��J����,��:���urױ�����|K�<u͵���O��9�M��'       "ύ�7,�t�������~�\��
���Rɗ:��y����gK�e��%   �^�      ���W������
�{d�@ѐ-��ѳu��EZJ�xI�˕"�i2D~o�L�3�B�8�B<y��n;��+������s^OAԥE�p��&�hȑ~��^��
�S�vئ�|�Im�Q��y���?�L*M�4� _i[����\6��S���k���ET�q$y�䦐�nZ|�6aZ���w.ڲ��ҋ�貵X�JX�Ao���WC�ɜ4��<OP���i��Z�W�mz�t��I�rDC�a��R�%��I�F�>��&��qJ2%��J[��>f춱�-n_pڞ!q�u~�G���5����Mϑz�iV�A+�
�I�؞�Ù�g,���K�s��IA�VP�?|������KϪ����k㴏��V4�֎�اr��2�������m�z!����{      �7ܸg�20������,z�D��UeI�%�~G4,fN�9�lL3��o�    �A1      ~���^R*c))������"_.����iq_�Ty����Y�L�����ƌ+���6��hX�e������n�G�����?�}S�nW`�����i���+�Q��Ͻ��u��YΣ�%SvMq{�q��5o�<9r���)K�,�k��z���f� 	��V�Z�r��ɲJ����m�i
������hٮ��v���x�ҝKb7}m��|?̑���V�ȳ'��=g���3z�h����44�������:��h����� D����j�4��>�����˥���>u�T񖻏���{�-)4��E0�ݬn�U�뼬�2z��@���h���z��`N;h_F��P���s�Y���/߉��6�2(�J�*&������󫛧��r5l�C�C�Q|���\: ���6��       |���o/�b��V��'�}�W�ŝK�tEΣ��Ln;Y��nj�W   `�b      ������+�L��9kFxyZ����Oe��N��?2%�$��7���'el�0NB���k�EX/
�t�vv�)�<x��)�9s댜�q��Z鿶�l9�E�7�/�3��6=x�@ޛ�	BԧEfP'O��^ҡd�a�[�u�1s�L���[v��u�A�����{�߳�O�l�I홠g�ZX��	�֥��A1Ξ�{5&,;����������'����nBa^�(N"i\�������z���Y�<
_��[΄>
�ׁ�&��7�z��~ߥ}R!K�m��c�!4V]>�R���K�-�b��/��;en�Ӗe�>�c׎Y��sV�Ň��d�9mw����s���v)���+m�L�ߪ~��5)��ah�Ұύ�6
|���w�/	b'��G��j�!WB�       ����cs_���f�g)/#����m�z��	�Y�PJf,�p�y�[S�Ř2c�   q�      D:r��ސ.e�H��}�(��u���Q���6�����($��M ��8���ΊJ�48FB���y��5Ġ�27��4�_�$��3����oƈ����'=�����
^_-��2(F}V�3�y��I�U��d�l;r��)z��7��=0�)���	�r�b֊���D��	�^k=v�Y<��a鑥b7g�aυ=.-c뙭��֑
Y+����_�m�0(F�]���	�i���e1���L��$L��ƽ�:� 0=v����2ަ�#���RKI�h�L��N��2��X�ﾰۥ��k��#�곕�`�r���jS;WmȊ�)m"����S���[�(�s�,��� x��<먾I�%������RcH9w�       �M:@�UP��ܸCj�)�X�n��Ni7E�Oj/�<    CP     @�E�����GH���]�vR%{�Q��xj�vo����l;�M���.�n�2Ӆ;���[�����Η0��p2&�(��d�lɲ��}]�m>2i��'B}��<#��L���!.$ j�rf�,>�Xj��=K�,�`Нъ4��ʥ�Kb'W��+�������j1�a{D��^V/o=sް���p���Z[�ո`c�a��.S���rղlw�98��#�Y�g����V��+�M���*e�d�Ǯ3�ݱdG���:����*l��׏��B`�
��zEZ$ަ�w˾�M�mJg,-Nm�u��L��9�&W�|V��a�K5d�ڽkb�&�����^*-
�pئדY�e���^����DC���g1a����O�d��+"�R�}�����آ���h0ո��ާ���.K%U�T���1V9^�[      ��]�w9����s�� /ݱ��W�y��֒���[��D���Gr_   `�b      ��O����Ǌ/�rT��%�K����u���#Y}|���?O^$/4EJ�z��R�50�v��f*���D�M^':�K��}e������~���A1�󪟛��Ϟ�+��1D;YQ�*gE�bbW�K⸉�{:g��K���${����;����a����
q��s��쭳�>Qz��V������/����)�~��:�� }�1��sT�\�����z>����e��	��>/���;'J����&�}��O���8��O��SZia{PL�����/?�ܥ�9������>�a�z��K��R5{U���sM�_�h�_i����ʟJ�i]Q���V��4P�_\�sф����)�F>�����U�V�y��BG�/u�Բ��ɐ8��<�ܖ��j�O       ߴ��:����W��S׫�;�yxG�����q�T�V��<�[����    ���     �(���{f�u��u�E��O��Q[F��]��H%v� -^ԩ��ޒ1qFi]���tD��A��I�J�*��|h���H@9S䔦���iW\�wݲ-e`Jۊ5��a���O�޽�]���Q�Ju�5(�s�Ζmz���Ë�n����缞�-��s��#W���=O��>N>����ҙJ��O�&�Q[Gɷo|+�b���V�����_��>�Bj�_����! �ﳢ�~w�����&��\�r���6Z|�<h0C��e��˗�����oڲ>���eZ�{q�����ca�l���
���!��{Ktt�:B��K�V�Z��<���oMh���y�;ET�O�2v�Xˠ���D4I9;�r�]z�^�y��H��r����K��e뙭      ���wy����G�2�-����>�:Ց�fJ��5   �g     EiȐ&C�J�*�i8� �[�O\:)�<}����3i����7���]l�k�Xl��{�E_�k���Ϟ
^o�-�NtZ`�ޫZ/��k�KE���P�e)g
��0��&Xş$��ܲ���Gr��]��U?_}�����>�:��ʛ*�t,�Ѳ}��Y�0�n�O�\����y&��j���T�R��]��1d����'��!?�,��Xe[�"�ވ��s�BM_i�p�7r�!틷�|�� �@b����t�y���݄v�/4��*(F�Y���ќ�lY�W��r*4v�{!�vN��)���	 �#�R�U=��(�w�����#����O��i.��ƌ+���/��h?ݎ~ud��w���?0v�+m�[!kZ$]��\�F��4�'a��� x�HS�r}���nb�O       �A���Y*���z�M�mȝ2��|P�I�$S�M�zy�	    �E�     �א�hz��}L�RT�-Zp�wy_9��׶c��ufʔ$�	��P��߅P�#~���/���� xJ��8�C��Zxp�l;�M��/�]��4hC��r��i˶&��/+����V���X|�cW����_�~����ʓgO½�hѢ�c�� �?��)����� mƷ��r�Ĉ#?��Ѳ���n|��~B�o/m�9޶�i
J�F�����2l�0�A1����9if�m�ܒ���
`%i��r��u��G����Mv8��b5e���� ���|/��$r�޽|ws������e�Z���÷�7b���hP�ն��N�C澩��$��X<A�o����|�H�B�L ����MC�F��4�C�u�����A�w���Ү�㐬�E[��X�Z�`~����U�R��C��w�Ή�^���gw�-%2���G�ێok�+       �eѡE�bT�bm�����m��b�Q�eJ�)f�"    �"(      
ɟ:��k=β(-*����.Ǯ_q��)�2�����'3�x��-LPBT�� ���,?.�Q�Z�U�%�߾_��L{k�e{�j�]
�Yyl�|Z�S�m�2�2/���
�vV�ZQ�4"vK?����wZ���^ۗ=@���nپ��z�ש���ӺJx}]�k����e�lm<�Q<EW���"��#\����Q-GI��,��m�\�������ҤPD�Hp�`�y��|6�3�C�^Ȗ,�|V�3S�z��aA�-;�L�_;.Y�e}��*$FM�1�* V�Y㟦���/e�I���*Y�d2��$������4���v��m�~�����a{��X��Vn@9s�	��3Ȝ��8��"WB����;� P������z�ɨ&f����X���p��������N,��w�K�P�u�ǶC��W�X��n*��~B��H��5�Χ���W�,�HC���b�l*���iY�����Zڄi-�VU��½���J�*YΣ��~5y�d      ���gX��_�vɷ廥���oк���4��m'   ،�     �(@�H�-����e�yD�H��o���o�����U��I���H���$s�̒&a۷C�Xޙ��,8�@|��״�J�nj���'Q�������������!0�/헼��:l/�������0?�������E�4���+Ԣz��2��L�+��ME4�DGk�������tz�-����u~0žVf�!�ХLs��f�7�z�X���O�~*��k�_�❋2i�$���{����Y�f���}tW�Z�U�������gAs޶�I�O${��<9X�ݻ&v)���)�o^��	!
o�^�� ���߹�8}=����b�y��=0WB�Fx�z{��[�S��L�3@��p�}?�����L�]�l�;/�z!��<�p���%}�����⿖�K�C�=�t��/_�(#�ߨ��������A2��`��y.<�P�n+m��qخ�ߑ�G��W�SGԴ�>��٫��U?7�gگ���=��S����GXFn)������rs-����%������)=��?W�����Zz��̇�?�
      �1��`����0�W�4�����H�U���� MF7��m&ʛ���cI��لg�zL�x)����   ^o�      ���qʨ���^�ߗu'�Ɏs;d��}����������5Y�e1�1E�1�ڻRLe�M��?��(62�<�R��VD���y�Z�^O�=�37Ϙp��w���+��O��'�'Q�D��2i��毎r�Q��Q:Si���i?������
�.-���񱭬G��@���b4xc��i�#�'��L�t[#oM|��B?���^:��l���Ϊ�1��8�A�f�c�ĝe	r���p-O��YZ���C��r����7�9���׵���)s�{3�3Ǟ��1^�m����t���������n`�����Lh=����^��9��ECδ�<�Ѭ�]��ه��տI�ܵM��-�����X7����8�#yi^�����/�[F�ύ��B�Ƿ��*��j�i&=��͟P���v9x���/�B��d��Qm�����3���O�}*�n��>=�<�c�r��<%2���l7!�s��qi�z^�x��N���|=���+�W$<�\�aj����<��ט]�v���¾q6v��&<�O�>�\���w�K��=�l沒5YV���o���GҴPS�y��&���~�#%3�4�v:�5 ^�-Y6s=��o�o���T,}1��%G��������P`����ԑ�e�Z>vʮ)� Y����J��=nXɖ<����׭����p��=�W�^Ҥ`��yZR'L����z0      �^c����_P�S�q���c���ci6��	ҷ
�]��
5�;bō%    A1      ~,g��2��Lɓ*O���A�0��|YulU����N�e\:`&]��w/�����zp�N�9I�����ga�!��dr�qϟ?��+���C��䍓r��Y���.y��f�s-.���T�V�x��M{k�|��;�rї&<��|j8�a:R.s9�����8���r���_���*XItZ ˎ,37����r����GC�*f�hF"jR��	�y����c�?dr���	ZL�M�o̴��N�xj�	��zv�9&>z���h��#�p[o��������Uxw��q�pr�+!/�S'O֥�[�}�5C�oろ�K�.aTiA��xsM��U��o��~V�3iS���0Hf�!�����M���+j�k���5�pj�����m�#��n*뺯3����q���*~ K�,5��5�ט� =?���/I�%1�C-f�I�'�A�p��	\�0Wh0 qc�5�]����5����&$D��W��I 	c'��)$O�<�O?V|��7j�(�a�����5r֐���ZΓ.Q:��q�l>��]�9F^\j����r:��(�3s�SwO���Fh��|ݨ@#�aj�79��A�u�	��|f��S��u�.G-]�i�F�=߯��M?uC�� j�ߨ�|Q�Yth�ٞ�'�ʹ��^�y[?��,��8ϗ�Tʄ�9�w]��������+=�X�83v�X�4��C��v�Ϣ����sA1i�	s��<���b��T�      <a���r��5����w��y'��5�I��h?���W�]�v    b�     �SZ�7��I'Q��q��=ST7h� �vv�x�����OH��z���~�gZ�W�&H�|��aο��n�5�W�׫EKˏ.7�ٓg�7r�!urב��+�D�d�@�BiI˱-M^d���ehS�����z��!*HҥL��U�Q�L�❋r��u��#�;�	��t�w��+Ǯ��P8ma3I���7-���Q�n-d��_8��W��4s�L[��ׂ^���Ad��-�I_�K���ҝK&t U`*�`��i�y�Q�M�'�O	�-�oy�([�῭���t���cd�����;i6��-=�:�ZKw^f��#�50��<�ݽfn�Ҁ;���a����㶏����`(��6k�,�<����t����h`�3%3�4�zS����ԝs˖3[�㤎Qz>o=��l|o�dI��r>=7�S�3)�~�n���5�Ί^���^Zm-�r��Ay�7d~��a�O�O�#h�}M}������1b
|��1k�-{/��aJB�c�:y���=�V        ����oxV���(�F��8���>
�RK��n��v   �날      ?��lÛ�X�����׎K���e�֑+�Y��	̨���BC�т��@�G���$�Y�� :�����v;z��y�u҂��%�K�2]_	�����A���2������Q[G�5����;l�`�2��ȆS�.��Y�ҙJ��^-��U�,�FFo-E�o	�h��3����a7v����^�f'����<��k�?}l��7��,����c�˂�������;4�'hx���uV�˪8��Lo?]*d���c�y�r�ȱ��b9}�dL���|3���ɛ��a�����S��hJݿ�����.��TX�&�l=�Մc�yxG��Nz-���r��u)S�),D�ab�y~�G�b��{*�YQ�t�cB{�;FlI�0��,=�T�Mhg������ʏuty~���       ���.�F�b�M�&    "��      ?�A��_P?S��.���%����ͨ"���
�PWm:�Ij�%�ܒ�D_��&�e�v,��r>`�P�%��xt{4��տ��k~�j٫I��=�~���,[G~Y�}��R��#���������~���O�>R7����<|�P�j,�;/�|��ٶ}Z��������:�}��g豢�CWI�!�e~��.[���rlK���D-�m2��Ll;Q�Ĉc�2��W���v��4P�꠪�Uͯ䳪�Y��M��4����B6��׵�v:_��|ե;����2e����*��HH�iU��G֡�I���M0���_�/�U6A7��d�e�z��4��L�5Y"�>�"����K�"-#m�ڧF�8v��Y�G&��BR�o/?���ٺB�e            �Y�      ������n?N�4X໥ߙ`�Ȗ9if����.Ͽ��n�9���~p[�"-��,�bI�bm,����&� 2
�t�.��e.'���3A/�+E.Y��r�4����uN��8LzU�e0�F�7�h�����v��9����_ZB��H�B�"�]��u��E��'v}*wN�Z�j����W���ޗ���m;�M�('c[���`�Ž�|LsS$�f�e�Wƴ#ْe�в���v|[�x�x���Y�G&� ���Mj��u�v\Fn)���"��C�o._��B�8l?q���8�B WL�5U�&L+urב�؁]���Z?H~X�C�틿�<y �ǵ�Y{g��0��v�zE>�����>N<���R���2���Z��yF:L� ˎ,�Ȧ��V�Z��^�HS�c��~܈-#L�<G�gYpp���:��;�:?*:{��h�mX���b>�            �,�b      �Ļeߕ~A��~���҄�x�HkQ_���\�_���B��|a���H�Y�e1�,�迿U�-�ed�nۺ��L�2&��o��&�'"4�ay��RyPe�p�� j�������73�#ѢE���{K�Q��\����B&� ��������=Z�<x�`鷪�)~�}�z��=�T�ZA��+U�W��i
����Ϟ���Q[G���S����Y�^=*����e��'U>���3��x�����'�s��������)�ka���ҭ\7I/�[�?t�|��+Y�]�g�Ҋ�/&�Wx_�o(	b'��25lׅ]���b���ĚH	!{�iQ��k�$g��۵�?���~�7�)N�8&D*(_�T�RAr��m��u_\r�9ߎ�6F�<�#��&�l��}G����~��\?Є�j�Ӯ߻.F40A1���/��r�^[jP�n޿)ޤ��B��ڹjK�rݥz��&@4"�����Fs���o�׮��*���F��z̄ jS��wݕ����c]
��m�            ���     �M5����w�0Č�~��}�j~%��Uvi^-R�Q�O�<-��\�2�|�GR�p8��6���*9q�D�n�L�9���o�_ڗh��i���N����#���u�hd#�=�ö�#�e�/��c幸P���̽3ͤǒڹkK�lUL��Q�LC[]>$Om�Ȓ�K������I��88��3��M�<{"+��0��+���PB�d*c���s�#EI/��2t[w��-��m��g������ܭs�-���|��!&��~��R.K9ɕ"�����M߫�7N���M���s<��������W�M�9_,�B~Z��	�	�$�2��,I�����=r�,?�\f�a�z+Pe��m�nB;�#�T�^Մ��X��K�����k�!?w��A�sq��<�R.ݹd�v��������x��X�/�~�[s���� ����$=����O�vO�t��~���a_��s�[uR��`��鋛���y�Y@�#��>���Å=&�`퉵r9��Df0}�t���&���_r�[��VC�t�����T�ZQ��+��'w�j9p���.Y|x��9��+��_���f�7Mp��>�n���'e�٭����cy,�>��˾w��=i?U�Dq��m��eM�DC6��������iߥ}�ߨ�y���u��y>����M��{ߙ8�����üEC�f��|�4���V�jd����������l�����x���{Ao����           @�     ��Jf,)�Z�r+$F�ޚ��L�=M��fΚҫZ/���c��Xx]h��{3ߓ	m&8lO7�Ln;��h�LdӀ��:ȢC�dp����1�
�-$�[�7�&Z${�R ��mܸ���j�N/$����&�����ޣ{r)�����zb;_�c��۬4@&0v��
��q��NC.nݿ�@O�`���IiA����k'F���9�y����m	�����`�t�S'Lm�����	��bF=��(&A�c�$L#�b�}��>�Ź�>hѴ'?7�Df�qDu(���MC��<#Q���Xr�*o��v�z�aj�0NBsl�c�#�8����c�2}���3��7??�_Ґ �^о~���̾��znѐ���o�/�P:���I�'Jo�Y�u�<x��E��Ru>o�j����'J����2}��1�y����aOo���z����4*��uSx��6��S�=���5%           �A1      >L�f��i��\��|uC���Sśt�Ǵ#ѣEwi~��-���;'J�R��Z�jۋg(.��"=f�o�m�tz�Lo?]
�-������hF�"J�:�S�������Ұ���̓�O�?����A��XҦh����!x�J��KIt�'�'9q��D%�O<~�             �#�      ����2��XI�0�ˏ9w��VK�]�'ޤ#���4_R�t�1�^�o�+J�ӷK���Q��u�u'֙�o��*���쎳�B�
�^·?�U�Vɜ�s ���y��"0�ö�w����s               �b      |TϪ=�R�J.���I�2����M�bɴ��I�4�z��mc�u���J�}a�LS�r�-F��[ge퉵�-7�ߔZCkɔvS�n���ZF�h�dx��R�_!9��  ��(�òmĖ���C               �      T<Cq���W.���-�7���Cb4 �fI���z܅��صc򺛳o�Ӡ�81���3�\�rr��!����K���d|��Ҥ`�p-#y��2��(�9��<�\  �
�d*#%2�pئ�a�	               ^�      ����2��`�ݵ�n�<{"��4�}���}[�[i[��ۏ�x�@d�������ϙd���N�L�2r9��x�㧏�����.Q:S�sT�VEZɸ�� ���G��m�-�#W�               ^�      ���e�J���\���Y��co���gҫZ�p=6a�����κ4_�dYeN�9RmH5	}*����i8��lzo�dN�9\��%�����zpK  �gE��f��Y�\?P               �� (     ���L!������'�$�o�Q�����7܏O�(�Ď[>y(�3w�RJf,i�b��UW�=�'�r9���u�ׅ+�'u���u�����!  ��x1��_������w_�-s�                "�     �!W�X�M�ҼW�^��f�'�֡D����ZF�q�t�Ҳ��*y��L�����U�YgIPH�<x�@�e�Ž�cf�bT��N�w�տɩ�  ��w�[��"�X��͒o����               DA1      >"E`
y��.ϯ!1�C/�7�)�F�j��D�=��jU��k�+E.�S=Gu��n�4�X?},�2z�hiQ������+ �|Z�S�6��  ��l�?���1bK��TR&S�����o+;���{�               Q�      ���+},��]�w���2a��&��|�-!1/��{Ao�z������������K˱-�ɳ'�-]�v�=q��طK�-?,�A��:+  �=�j����>{*��v��ϟ               Q�      ��x1�I�2]\�W�?��xSp�`�d�m!1J_��� �S��u�!AM6��l"�[?���[�㧏�N�<-=����ot���cĖn����?  ��~����3[               �A1      >�y��(N"�杰c��zD��G��G�?$Z�h�/�cɎ2q�DYvd��n:��,��&��2�j*qbƑ�����'��n*�Wx_r����c;�� _.�R=}$  ��9��H��               �A1      >�k��.����S�n�w�-�T�D~���ǖ=Zt��v������v\^i��/j|a˲������4<HB�Jd�}��e�˨��~l���~��2u�T ����2B�M�&O�=               �.�      xY�4�dƒ.�;e�9x��x�W5��/k~���$��T�w�/UU��/HT+ �Lh=A�Id�2+g�,s;Εz��y%,f��qҧzɑ<�ۏ.LP �/=�\�].?��YZ$               ���     ���<ﯫ~��=Zt�w�K�r�"m��R�﬐ZCkɩ�$���vhӡR)[%ۗ��\�y�����ܸC"��gO��e�ˈ�#�~l��UMX��{����<�#SvMq�v��	�ش��$F�WV��յ{�dυ=���Z9{�                �BP     ��5�����]9$[�l��;Fl�r�4-�T"���l~�4�D֜X#QM̀�2��HiU����Q&SY�m��1�H/\�}��T�'I�­�i~���d����~n_�fc�	 ����5               �*�b      �(S�LR8ma�����Ȕ0NB��~�T�^U�%e`JY�u�|��[�~������
�%J'�[���Y+z|]�S�u=�I�a����Y?},�wM�n庹���                 ��b      ��^�z.����s�}�D�T	RɂN�H�"�m1b�׵�����K��e㩍��Zn!�����G�:3&�(k���z!�"���c|��bj�%�bɣ��                  �AP     �U�R���6��$Ǯ�Ȑ;en���<ɚ,���b�����eҮI�υ���W��?)�����T�Q�+�O/�,�L��n*�̏�un8�A�_;���?V|)���߇                 ؉�      /*���K�-9�D"���Li7E��M"�(Z�hҢpiZ��L�3M~^��l=�U|Y��e�g՞R/O=���/f<��a��;�]�i������s��s������ǖ�\��                 ��!(     �K2&�(��wi�u'׉�u*�I�9Pb�_=@�jf��v��-#e���r��U���2�\*X
�) �$F�2��Pə"�|6�3y���G׷�Ȳp�h�N�U�                  �AP     ��h�+�>{*Om��vD�]���+�T�D�Q�tE��k�_M����se������~y��y�l���6T�VE�o e2�1��/���ǒ=yvi3���}t�c��tz�<y��Ը���                 �날      /)���K��Wn=��m�(cZ������Ӱ��Y+��z?ɍ�7d���&dg��}�u<~��	މ����K�d�$��R0mA)���	�I'��}�W��J��/�o���:4�f繝R<Cq��:AjI�B��^            ���w�Q\o��oHB������]�\K�ҖiK�O�8(��N^�	\B<�{��
dg}�@��\!{Μ�����<��b��������M�t���`���N����R�'"OgO4*�HM�D�D�v�m�"?�x�ШP�F�":6��������ƑI�K�{fW�%�RYJ�Ч���f8v��M��/h��A1B�#�!"""""""""""""""""""""""��b��������I~��F����՗ݰ@C��0_�$'������USR���K<	����O�m�j�ӥN�~�B�,��z/���̷���`P�A&�'�}���������������������������CDDDDDDD�(�R�!w��F����Ֆ�"E
�5?��)S�%	����?�~y;N�9���N���K�����_��l�ِ'm�)���UՔ�5�U�������C�,�1x�`����Z�~�#_�| """""""""""""""""""""""�1(��������(d��
G{G��Z+(���s��A��-�¢�p5�*��?AdL$��=���<�=Ք�-#�\��;|�0f������γ;F��2A��Դ��6L�7A��P-��D��7]^����*��x��h3��>�5��66L������������������������(9`PQ"H�����)��4�-F.�\H
�?h?v_ٍAp��%�
�ep���U�I�,�а@C��Vv)�𾋍�ŲS�0�<^?h�q_�|��wO�釭?��O�>�T���AD�T�UGE��[�`KI8г�g*�����>!"""�j2
_T�Bg[��}0��ti���?ޭ�m�ɥh;�-�������������������6CDDDDDDD�|\}��'��a�)R೪�adÑHe�
�$���j,:�;/�DTl��c����-��;����ӢI�&����(���G������q��q�/��ͣj�eV�~����JV������7ǘ�cT(�%$�H�"&�c���������$�4�wn�T�d���'<�=�d�>���4�)�>��s�����k�{��J�&P(}!�P�}��5�������q'䎺�y58,DDDDDDDDDDDD���\���쥾�x������b�����������^<2{�\�aN�9hX�!l�䝓�gV�Z���p��-����j���>��9>*�*vK�xPb��oqȊ��hq��a�w,~��z��
M%�B���B�<��eq<}h�:1(�(�8�9 �guR���R�H��KR�,!_AO�&�����}u���I��S��G�����E�oDD����ʧ(������~&$<!�Nb"! �لtsvpFUߪ������)�Y\\��_�Uv�R��2��z���t���[�/h�o����ᛇ���R�u�/u��T��k�,�P:Ki�z�j���?v��`�U%g���CB���<HKDDDDDDDDDD�����;y5�j����
�Whd(��9��w`��E���������:CDDDDDDD�����3�p�A���f&2�e��칲���?l��-A�P\?���F��0��xU(�T�ym�Q����A��Y���OƟ-�D圕�G^O'??	��~��Ӭ1̹:}�4�H3,:Dd<)4����*z.��rx��~"�&A��p��q칺G����?��g��*$�V.>���W��B�헶#*6
DDD�Y7o]����Y�ܡ�=%`"�e�3��e�bmЬP3T�UM�Ř������R���M=0���N�+d�Tc��E�\�M�O�E%(G������o;CDL���;Jf)�:F~���eTX���2(�@��]�7����A1DDDDDDDDDD�X�zd�/~A��m�_��誂�e�����x~#���5N�9"""""��b���������wjo��Eǚ#oc��E�ҝa+r��/����C@P ʎ/���>��h8�;!)�qh��ȘH$'�D�)��e�/�C��
A����lèݣ����n�����_��tX�b���h��]�W��22i^	�ɝ6��Zk�n;s���3s��Ž��@֑/]>5�*�K=��&a��xUXNDDd+rl ���q%��
����_f����3���g�������ː�K��%�!#6��Ā�	�*R�H�����5���K������R�Zmu��,GBKg-�:&O�<F����l�ФP�7]^|/�%�źB"B�E��<�����γ;F�+���$����	�����?�m?%��Y�A1DDDDDDDD��ؠ�����lY�%&���i2��J��o�c��ETl�|I<y�d���R��vR0f�^?8��M�_w����bA�����1䄁�j|�f����Ҟ&]���"T'��D����ʩޗ��t�j�s���k�_�}��U!��=Y�����U쇁�b��� ""��\޹0���*4F��\?��`V�Y�+� ˒���$�z���o���?���\\���R4*�Ȫ�J�`�� �-�ê3��:v�l��~���������������X�b�<��@���%@�g������7`��a8��ޱe�ojc�:�Ō$���O�=�)�G�CDDDDDDD���1&\CBR���E���SwO�ゎ8s����wN����X�X]q$1I�|i���}�'�ǒNKT�9�ˇ=��`R�$u�_D�08Ot�yA1ƾW��'{'�5\��
����..?������i�Sf�"E
x8y���GgvϬ�	2�^�;~��;F�����z2�eĲ��0�>_�y�#"�O���1��5�T��.�]�/S>���u��U�a� ǁ���Bݼum2����gǖs[���Z���Cb������������D���uF� cI�f���~���0���.?��_���Զx[�E�����H��<΃���M��3�'�����CDDDDDDD�R�~��&����n��=T������EpdL$�����bN,�[��EZ&�:�92��y%$"�f5�c0��@�Ɛ����I�&�i8�X�7����#]`%Ge��łT��.�����S˱���_�GpX��1=�=Q9ge��S����#�1���P����ӡ�@�5�� 8�;� ""J�9rR�IputU�pߣ��$�nNn*d�������f,��=7�ꤪFl�jZ�iF���}�~y�
~���2�gB���Q)G%��-�:Y�i)*L���Z�����������(鐿����/t)���1��,9�,�c���Ƿ��Bdr!#[�V�^?���#�r�r�g�i�/n��@DDDDĠ"""""""�D��θ���>������H0@�
}Ք:Uj[��
�齼7�>�7����(����;�WWIH�e��X�/!D���������/
��;.���1t�Pl��Mg���qf�Ϡ����$�I޳��#3z�hl��UoИ.O`ݹuj�b����&>���o������~�C���}��D}h�=���7��WN��p�@��UQ���T�SwOa��� ""����ta�Q}�󡧋'
�P�!c���W\�����<�9�����6�}u���_��ޫ{p- 7��DL\L�~�޾��[�KwF�\��[2sILn9]���.r·���o��R��KN,�������=����qvpƒNKPz\i��$��?��{[x��!�����������^���/�ļ���߫s��!�>�n;���F�Mj6�߀�!�ADDDDD�cPQ"�+�C�����c����t�D圕Q*K)�W�����bN�ڏ���I�]V�����b�,�a�C���R�꼯����
q�d�E�H����[�3p'&�O����_U��U�Ro�TƽW�>tv)�0��4�(�#^���3h� �q�*˒m�����T<Sq�m6��"h	��ۊf*���z�,������Ҟ&�#�?	}kY�%z���Q�H��s�q�����6�ژ4��
g(���~��+|�t������{g���}�����{�?v��
���vΑ9j�P8cH�L���F�l�0���XD�<*���b�C�q���f��������o��a����@�>��`ՙUX�D3�._�|����#!]	����d��%�/�[pl�X������������l�v��Rc��Ɠ���<��Q�r���n��#�>
TA�O��"�\����k�9�r!����K{�������Ǡ"""""""�&Wo�����%�C��"W�1�.?�����Hp��O#�G6�/ﳵ��xߍ�3/����&�-�f�j
Ʈ�]��$�F�����_�U%gN�NX�-
�x��Q/T����Չ7�p��	ԜZKv���U��+��t���7��o���pP|򼜻NM������_���)������F�ar(�+��9u���d�#W�Te�ޫ=�;���?'���˗/���jL�?;.��8J��ʎ/�)MA�2]����a���j����ѯo��K�Wӿ��j���f4����nWǟ��<�K�؂�
�9z�(��:�'�O^���Rއ�"""""""""""[���l����̑�3�:?E.l�Y��4�`��q�;�B��TྜoҽlwuQ"-~�����o>��������
�b���������Ȇ#�~��J�5��|/Cb^���>Z�����]J;�-G�/W	�P��3�d��տ��xѪh+��iV���V�ޫ{A�ɉ=�;-V(��`  ��IDAT�7Iq�l�lU��&)f���|\��NKP&k��mM5��NK�bN��ŀ�������U�󪮫�������C���#YB��>_�9��<���#e���};���|��?DrL����?>y��ƍ��PW�tvpF��m5���\�rT¾k�,Z^.�\�\��f�<��7)$�9����_`R�I:��n	�밠,u��5�y�u0�Lo���6�N"_�|��E�����9u�F��iU(��h�R����}&�L:�뺸+��\�w�ѱ��;�����u^�y�<9��k��s$������8�!"""""""J@r���E[#)�b�Sj �Q �w�o�8�q���6_��?>4J�'m4/�I���@���Ua'Qr"W}��zz���]���|Ns<�x���#żU'U�B����Q�4.�3��D�%��>5��s�U����4�8�;�m��C3ADDd��/R'�Jp�9	W��������'9	����6?�e�,��YK� -�K��8(F>��E�n0�>4{�)��Р����loS�������f/C����������������#a.��9��7Ǻ��T@̻�d,�a5��]�v���7U�YW��ěGƩ7����u�w
�'W�ƞ�غ�.֚A1DDDDD&`PQ�B�QMF��b5)x�M�j�A�ļ2b�Ud��H�\s�α�(.���F��~���_]�>�(��,:����(9\m0�����mkϮE�ymi�X)S�����]���ԩR#:.����Q�Bn5������֘�z�[�&' �����d����ѯb?��ɯ٧n޺�!""�� ��~(���f��!��84��ː�!�`y��}j�e�2��s�Κ�������!�C7��w�l��m�*��6%���Q3wM���7���V:b^9}�4:,��C��a�S�Wf����|�ݖ����\��vz�i�qL��x���q���� """""�CDDDDDDD� rz�T_�V�Q	I���t\��fWVO,a�a�rݗX�u�UǍ����v�*	j;�-�}v���H*f���^9���_�]��K�_޺mg�N�Cb$�Z�jhR���SьE�h��_c.=���k��������:��{�ײ^pwrG�"-_��s���?h?�������p¾	��r�f�r�ˁ��Ț�����"�E�}Je)'{'�'���gV�a�C�sM��=oڼ*�E>w�C�|d~-c��QA/��se��<��YK�l�P�����zMQ�$�]�wNࣹ}��'��5&4�����7&U�g4,q��u��=
?��!^�\|Oέ\uf������0��X�R��g�?Օ6����b��5��>�Z}�-W��%'� �q>d�]Ơ5�0��L$v���Ϩ��.:-�Oo��C%ſ;.T��W�JN�g77x"�v����+�W!eƒ|Jf.��������쟂헷��/A'2���n���o��\]jA�(�GA<C�m��Mo{V��6/�wvpF~��j��I]�K&y=H�ZXT�?������R'~%..(��(
�P'��9�!�S�xI�QL\�E<SW��d�o<���ޒ�
��L_�2�5տ'���d}��?��7'鐆l�P<sq�x�x��(y|�G<ǵ�������cI*�MN�,��0�˫��^.^걗m��n������gq��$�`:��J X>�|ȝ6��ox:{�� �٫��b��������{fG��E�'m�O�^-[B)�=FГ �~\ %]�ϯGtl�[�oJe�
�3V!!d:�v�1T�2]u��Iι�s��9�o��&ۀ�V�Z���#��
�+  ( DDDDDDDDDDD����]�{�~+������ѽlw�������u���Qg�Π�b��1(������H�!"""""""��2sr���]�7��M6aԞQ�Pɗ��o�����ژs��Ar0��,4*�-
�@RRշ*N|qBf콺D�o�|�
�_�Е6�ڨ�_}$HiF��p�R���hY�%<�=t�	�h;�-�~\��Y�	=_��
�_�@� a�H!y�,����z��z���[�sVF�H�"����c�ŭXyz%֞]���+���S�{-��P�׺:�Y�㷏� ��A��1��!��ɺ�"�e'�Ż]�4z��%;�L�2w	��rq��&9�Il�ӯb?�.��22��I��>�Z�T�X��(�2m��A�**�4$���㋰��:>dMsTD��]t��ܩ�	�%ۄz��{����>�S����$`fR�I:���z���~��MB->��1�j�b������������7���+�
�[kR�	l���v�m���G$7r\q���:Ԓ�3����.}Q��m����NGrv��E��޿Z$ܧF����oDxt8�e����|����"�$�%<���.�Ё�LO`&L���������p��M�q�rT��&�!"""""�0(�������������o�j���A�t_�=I���skq%��*p���'ױ��n$}��U���2ڊRl�tTaD)����ۅ����\МG�w��3���Y�k+�]�x��X���m��¬C�I���C͠���f�2�d,�v�۩���is[4���7ڗh��{����]��PS�Ff��K`\�q*(���R�\�rjPy�Z�m��a��1&�U��iZA���fP��'�V苟���?c�8����$�f��*|!1Hp�7��Q�r�k,�_w+�MM���n0�=���������O�>*,�T2O�b��t5��
�����v�,aGZ�!	�z7(�f��|<
g(l�2t�$�Hk��nPLF���d�چ*�f?y�h-Og"(����.?l�ɕ����dH�A�����zn��\��b�?���]��(��<\]5����Ú�~�1h��t�KhՈ-#@DDDDDDDDDDD	G����}a���\�ά��VSu~/("���z��uLgP�|�KDDDDD�aP��IQ��t~����\�Sy褠wΑ9�@�R��/B��8$&$�c��ER�d�������z`*�>CkU'�����>�>2[���j3K1�#�-�/m�ᛇ���#5	w'wU^(C!�!��ԩR���hг\O��S[�.�?��0t]��ߓ�'z۝�,����&K�B^7c��QAt���ǭ:�����7���v)�`m2~ろUp���*$hmy�娕��E�H�Á����1jϨ���뺯S�K�,�R=���z+H��d�(�ɑG�crk���ŜvsнlwtZ�	7��@B������}25,,�����f����˕c����\�깪�p�K/�V*d��#WE�ux��Ga�����r����5,*̬q+���7��k���� ͠�RYJ��epEDDDDDDDDDDD	#m괚��o6{\9�D.�&|x��{��z���;'u���l�w�DDDDD��b���������(�cl�ML%eRԿ��:$�?��A�OL���V$7��OB��P0}A��'E�rR�����#�EωL�h�c��� z��{�cɎ��0�����0}!1�.l��[�7�d gg�Юx;�.���u�fN}q��{�C��n�w���:H��������-?�O~ؚ,c���h?�=V�Ym�1]]���FT�Y�+���ξ;-XyEC~o�;r�͍~+�����IȐ�J(�5H���%j[7f�X���f���Bil��oUt-�T!^�������V�N�:f͟2���X�4��x����\����.��]3^?	��U��\�%lEv�l��7��Dr���.�����������Z2sIͶg��I��&A1���$����# """"""""""��!�'j������������>��~���L��QrƠ""""""""+Ie�
+���($&�qn?�_/_dt�[���u����xz����r��f���Hn����cs���5��l�8��������VSQ=Wu�Ɲ�|�>��S�A�>�^��ڗ����z��sB���U��t�E�D����Xt|�I����֫I��%�r�К�kТp���(�#�� iK�:�����O�>p�w²���lv3l<�Ѣ�$<B�D��	\Z�m��Bb�$�#a1�$ǡzn�ZH�+���n2Z_L�7�j��U��َb����ҹ�S�Dg6�ޫ{m�	h��q��!1"���3G��mձ�<W�X��Suň.������ 2&����6��h�O;0ə����v��C�+���f�����+���f۱��l"v��!��N�!""""""""""J8Z���=,=��:o��zk���Q��v������?�!"""""""�)��~.j�m��R(6`� �;�N�.��-��ĴV�����V�-$7�.m�((&�Z�M�X�[.n���Q>{y���?�����.>���Sk�[�n�t���إ�������#쾲D�%:�������+A�ZL�Y�/�ݵ��Ɓ�,Z9hɉ%F��{��ѡd|��;�|�_V��*tB��s�}U�7=�|��wN�0�k��!$<!!��1WGWu�.		)���e/�,�Y�g���:.B��%p5�����q��U�!��î�]����>����^D�P�9y���S���P�3FьE��c�����g��{
�oP�-�1y��q��Y=��
5������?��1.=����� �ٯf���M��A�� �In>����(,#�i9�jT���F�#���G��ta���+� ;��D��E��������>�{~�/��ދ�<Hx�L��?u��*�܄r�y��a����=}��Ї8{���F�������z��z��>���T�}�cN�9�!1�X�}\-�዇j;%W,,�S E3Uag�.w���굮+Sw���O,����􃋃��6	��|�������'�O@��G�<�4�%T%&.��q%�/�WN�vٗ�����ն_k��7]^�69.)���
2��O���5"�#ن�zzKm�N�=�;������������~N9�RZc�F����J��{DDDDD�b���������`dÑhW����I��Ā��q�*n~���V�ʣ+���*H�	��w,��헷�z?�=��&g#w�TE�搢�����M^��{���"�E�H����X�m5�O(����7%2�x��V����߻|o��ʡ��ߊ~�ĘC�y%�
ry�R���RYJ��ͣ��j殩�]���`-�����?Xyz%֜]����#��5r�@���T��V��~Mo5����'�����N�}���<�O2u[/���WD�BMмps�I��P%g��ױ�����/��M��lѷb_|W�;�j�5�{����I�2�Q6[�x�K������;�9�x��*�pH�!Te�
6�E�	$):��E�H�����!1�oƯ;��sk����]�����Vs�
��En_�e%J�+e� ����O�>�n������S���Ru�^��_����j�ɚ�2��,8�;�k�zi+�����j��)'�6)�$^ Ltl4f��o�|�s>ٟ�"(F��"��u��_�������<m�����]L�!a\��i��s&�%aT���I�*嬄u�ס�o���$TK��$@x���V=$"""""""""��\�A�7�=4��Z�M����%G�!"""""""�P���e�/M��a�Ct[��o��s��	��2����5���7���/��V��67tG
�3)V��C�غ|��U$���KT��&6��>��R�'����I�\���}���!�ѿR�m�Ϭ�ܣs�d}��X�ᵆ��M��bt��}���	u�v`��SƙC�۝�;�� �h=��3��[+O-��_�/l6y9-
��,D��H��U��9$������l�:y�`P�Ax	��r�U:k�x�M
����~fp_(� ̞1X{v�*0��_g?9�OB=J�+m�������_�_B`��e֜Y�B�ҦN���<�㚍C����^W����[W�]��>^�
2�<3��l�W!��@�B
���ߪ�k��'~В\=�_38���n�w0���'*���m7��@����q�!��Yx|�ζ�f`X�a*��]�����K/�Z�9�:f���Q!�ə3��Ϲ��@�� ���k���T�}bH�z�o>�	[����VparW.[9�瑠-	���A��5z�h<
"""""""""""C��P��1���9��b��������,��=涟���M�ϭ�lv3��m������j�Uѐ%��Գ�Fr%E�R�(���H�Œr2���l3Ӥ��XY���!�}W�U����cT����f,����,7/l�(�T�����[/m��[:Ki�N�[g��%��w�#�k��Q��}T��xa�l����y���'�O`-�.lR�^{?ًl�t�Zc�YA14�l��sCb�%�4y�����[�@���|R^�@ԛ^����)�����Y�g������!1o���ƳcG��A}m��UǺ�#�P_��Z�]B�Ϩo�1��:֚Z+��PI�|Q���r�2��Lu\��Wջ�貺����1�x�y�����sT�r=U����*�K�M�Ø�`�/�}���j�URA��Q���6i�}�l�͑>Mz���d+2�� 4�!M��I0�7��Q���6S�[�8������������������>�!"""""""2�}J{,�[oo��[~j9�,ꂰ�0��G�Fa��i������\�:"&�ٙ{g������n�ɥ�|�f��.R�oja�}p��],� v��&z��;����/Jf)���/�^���#�}��4$�����HL�|�o��K�~/��$�mh�W��������ͣ/k�Α���O��������c�v	���Ua��*���ğ��=3�'I�����R��pfC����t��`�9G� 6.�0e���8��:bu��:�%$D
���Ģ�o�~{��y׳�g*��Ҡ���p����>;�^����_a�ꁰ������	 ��&WS?�Eutň����Mߨ���ܝ�Ѷx[����#9���"Zi����A���	#j�w�}��������Ko��[ي���YF�i���Y�f踰#��?�b���������$E�UrV1i�
t��}MΐpK�b��u��YH���;k�|�|={���y�s�ҹtg��Y~�Y�Zvr"�#���r�"p}�����?�<���N���gy��l��c�5���VN��w!�I�F�@L_P�.E�..6�x�|T�#�}rsr���u_ �������ÐC�I�G��-TH�)2�ɠ��c���}��D/��쇘���9u�F���k��]�K�x|�镰�{��a�ơ�����~Z����S�SB]*d���%z.�;k�Q�����W��w�q��C�������$xH�迪�UCbĶK�p%�
ry�ז�5Zia��?�R~j��K�� l���UV��X�eR�H���M'��6��H�%�~�Yl
��&Ǳ$*�nd;�ϓ�P��p��MQ�Ơ""""""""3��ʉojc�<�����U�)�Rؘ�+̱��*^y���
�e�|R ��ktP���q��e�;��u���������F���A�������k���z��)��v�k�H
���P	�8s��+;4���T�u��1�桙�se����×տԹ�����IA12F��iu�=z��	�p��%��5r�Ht)��@�7�~�A1�7ǳ�gVk����]�%ۉN�:a��aF��qŏ5��]ۧ�I��^ڪBm�%�M5�����L	�z�	m��6y=I���S�G�?t��.��*%2����g��������-��z���#�=D���ޏ����f��Ǿ��E�H�Fo���ڊ��e���|&�}��=�Y�38�9��OO�Q�/�}w�ꤪ*̍�����������������/��ab��pvp6�����ʁ����}x6~l�|�������^U����a����f��`����O0y�v��a֡Y�~y;��2o�~���f_��v��;,���kH
���
�x��XCj1�OOܝ�������K���e����d�'x_H���
��V.^[�leMK���Z^�����D��x��VO�����t���>ܜܬ�"$�`���VO�O�N�B����kctP���VE[i��ٴ0GcI𑮠� ��<}�姖#1L
�d���3�O�ҹM�����c0,M���˫m�.ѱ����_Hnd?�y��ѥtا4|j����s�6�~�5\�]��uqW�}vע�H�>1�CA1��|�$q�ŭ������8�<�b�t��m^�Q-W5�.����Ǘy�wY�Sj��%O�!"""""""2Q��-Ш@#��o��=���($F�qX��V)�����C��"~	^�W��J�@�,s⾉(��z��a����FCdL$���ԩR��{hd�޾Z��I%���������d-�&[Yqj�,�YL�T�}\gP���2�g���F�%��Ln���.���w���������$K-<�?��)R����h�*9�`��V[޲�ˬ^����B�cY_o_5]�jp	k�
l����
���=W�� <�xm5rװ�$d21 �u���V��/��'��s�����ݫ|/|��+���]��fۺs�,�H,�z�����~NN�t�T��B
�r����_�vC�Y�gaW�.��$nv��z�q�㬲}6�b(���b�wP̩��0���9�F퇌%�X2�=:�������6��WC+娄��|g�`4""""""""""""""""J�CDDDDDDDd)��l����_A���R�)c�c����{B"B̚���ۓ�M6cJ��!�W�G�L�Q*K)��˗.V�?v�����Ё��0;N�N�m�n�M�����M~~��&L�8T.1<}�����kRP̥��t�H8ҴV��bNX��-9���c�q���GP6[Y���rU�jP�ғKam��$��
�Х�oU��b�o�ٶ��J���$�)�Z ���-�GVU����#�,k���H�/lFl\�M�1��T�A1�k��f�7ff�;��m���L��J����l��2^?����x�_�m���W����nj��i�c��9CcZ��ћGQ~By�q�ⱞ�?U�Y[�y�f�z�Y�K�����؉�������������������y�������ٍ���sZ��Xk�rˬ�$ԃ��2EJ��sHɠ�7�è~������B?����M����_b���x�DIQdl�[���O��W_�*�F�"�I�ڛlY��>���������&Z�X��$t���fdL�f[F��&-sg�NT�U]g[ろ����[�^DRv �mƽ~@3(F�ԬE�B�8k����
Z�އr��i�����?����2+{,^���}�AB-lM^�'���|�sM�EZ`�	�Ö�J�ivH ����A��ڏ�3��m2���v�ݡ�b��}vm�1+�HCAir�h��P߱�xB�l���cV�γ;�3�����^�zi�Ke�
#�P������������������(�aP���0���W�q8N�=e��#EiƆz$�^�<u�Ԡ�\r�^<B��i���fP�������5�4c�|RtܷB_��3DIѻ!F��\����)R�k�r��Hl�hT��$5!!�w��n�rS�z��d�(��
g(����p��9�Ye�4Ų���}��5jj殉�_�U!xs��U�8I-dG�P$L�$\C�<��r��e�E���>h�s$$_�|���-���fq�b�e�mDbH��1e�Lk5Mg[���
���0��Ľ��M�'&ퟄ�������g��}�#O�<�}�ÂQgzRd-��$L�Y�3؂��N�Z�l�$/C�hR��f����b��aV��MDDDDDDDDDDDDDDDDI�b���������ԩT'���aT�=W�`��x�._�9�
�N�NF�#Ş�#���enP�̻:�"4�a��}\���s��o���b���4���1y�d�G��(�		; �[;R$,A�Ӥ�ז�-�
TJl>�>o��X�I��Ll1}*�A���p���Yn6�l�Q��*,��a-�
��%�ߥ'��]�v�}�Rڡq��j����ᛇ���Vl��GnQA-�����6�9y�f��;�;Z%�A�rl9vv��痀#y�Ck��T�����}��r�!�H`BXx|!~o�����F�*�C��U.[9�cCy?�>2��}��aȆ!��d<	@��{�
W�"a-�gԷ�����͔���`PL,�b�-&.~�py��x�֯��7�k�@T""""""""""R<�=0���ƨ�����Ke)e��o��[������2�!"""""""2���9̨�R��ɪO�~�z���������y��:���bTcevˌ�/��eLP�-B�$������o/R�Ha�|R�ݫ\/4C��\{|���ͫ�`p�Π����cW�.$��is������H`��	�pstC&�LFl�P������{u/lEN����O*h���4s�S��ٚ���gYܳ�+�w����]��T���`�����Q/���ܱ��r�E�����F�ǝg�s�90�������X$P�$d"�$Բ%|q�?�пR�xm�Z�Y��
11V��5�֜Y�����ݏ�8�s�����A��ϒ�{m�X�Ƴ��ͣV_���V������؉���������g�?5�4/ܜA1DDDDDDDDDD�H����~��د��'""""���A1DDDDDDDDFh��A��w-��O����_��JSH�4�'�{f��eP�.=�d���&�¾k����4.�ؤ��WU�QR�����5���`���P^�z��T�Q)��U}�b�ΑHLܑ7�A7����C����\�Ө�ƒ�'�嫇Υ:�-*���u�סƔ8v��o-
���63�Ia	͔@�W�=��泛ccύ�q�1i^)d����jfѱ�8t���\��'�A��ڳH��*��t��JP�-���-A+��������#a8I��Bd���q���H��M=0UgP��Z�+���-�b��#�ж��j�O?8�;	 5�u!a"Oß���S�����p������zn@��e4���圖��o�u0t<eN8����o�ݐ��ن�P�x�x�l/����}'}xCDDDDDDDd�ne��O�\~�����C
�Mq��q�2�e2{��`g�Nпn?�m����WS|��;4*�Ȥ�<i�p	�!JjN�;���k��K`L~��8��ξ;.���*���^3OMju;����V�g*�4�i^�~��i$G�%��2��;틷��5�Zܜܰ��R�[Ҫ!+��fc�2EJ�O$���RX�i	*�h�8v��cF7���7��4	[�	i�)Ɨ �Tv�t�[+�Ė��P���+v��}�k��^D�@bH����q�ս*��]ռps,=���8KvT!C�>
Ď�x�I�K�ƅ����vgm��:C�^��~����������S��L�*�P��� ۑ��[/nE��u��~�P�B6	$"""""""""""""""���A1DDDDDDDDH�U����;1`"�>�ٺDǙ�q%�
�?Y=��=o��%@�1&�A1R���v��[Ǥ����ΠJ��X�UP���k�l��!!pwr�v	����g�n0K��5��]�Wr���K,<�Pm�6�ڌ��u����[N��B?�,�m��l�Q�Z���]GWTح��T`MXtb�b��{4��]�t���
��ʓ*�M�6���O*���)�ѴPS4)��έC�U�q��MX[XTlI�O�;(&����M^F�����}��������\�;e��A1�w��F�H?-3�P�7"s9�;be���o��2ݗt���+m�.����۞�3�͖�u�"��ٖi�_o_�%��O��ʕ+���������	�۳������{""""""""�J�����`�ȘH��o�u1%xC
��G>��p��f�[2sI��>�k��-�bĄ}L�i]�5����P%%���+��&��+��Y�f��j��k��������8u�C������A1�����l����Mg��%;�b�y�̳hY�6��4�!1Q�QXrb�
b��������n�a+� ���2T�U]JwA����$�B	����":-��6Ú\R����/��,��v������]��!����G�4��I`Z�(Ps�r�ʡX�b:�d7���K������__����,�c�~�A����[�jH6��k��@�e( 8�{Q�x���lق�g��l�s�ҤI�:8F�W������ ""2�b���������Z��Q���Z
mɔ���!�Ao+������P������!�e�M�a������2�e2zWGWd��aJj����A������+�_o_\������cЧB�N����%�ay��(3�B"B�����lֲ�ƞ�{@�9w��,�U]Wi��l,֟[�'�O�^��~��"��Z���߃�R;���I8����j�Oi�RYJ��j�����4�iL3m�X�m-�j�m��Ym]��`+N�NHe�J�=":�*��
2���C���%�I����4�)�4�2��,�5<^��(ի\/�0Ds���{k��:�J�W��a���;�G�B�4�HH�'�>��C3d�n��BL\���/��rl)�L-�3(��m��3.%���`̝;W��h�]����x����*4���G����x$#��w�0""J�CDDDDDDD�G�(���Q}�:�lM
��u?Զ�5���_0�C
��窎M6���y7����� E��T�Ĥ��l Jr�=%�c�+�W����W��W���_��~��������̓��h>�9Z�^��4��~`�o}1���2�Β��gVc��hW���voo����/�_�3��~��R��gy��)��t�DB��ʡ��4r�HU�_4cQT�YU|����Ӥ7j,;,��F��'׭�~�����]o���VY�-���P��� �i2h�kQ�5��t�1D���յLW|��[��y-�-�Vs�i���)S��춳ѦX����)�� ��1����q�.9�r�d��7}'^|xd[���$H��������������VTT�͛�7$�111x���egg��b$4F�c^ȼ�)!3DD�|q/@DDDDDDD�Gݼu��'E����ak�oD�D��S.[9�Ǩ��>�b�?c�b\S����+N�09(�V�Z�Oio�} JH8�*(F�(����w������ݿ�n��*��]�2��O㇭?`���3z=�@Z�'T#A���68������{H�OW�������Cg{���1i�$=2y�VE[��M�ˏ.�e[+$Fx�x!1�������j��o�z���ZM5E�R���#���ݝ��}���mI7�����Jf7���C��߳�r��g��d�����0��ӛ�m�~��'�O@�	i�xa�
�{��[�n����ձdG��F�^��+�Ad*ه�l3S�?��07��$�c��iŔ�RR.�~њ}���/ٖ���+1 """""""""��c��-H18��(qm߾O�>�-���"88XM��I��uh̛22�Nm�=Q�cP��Ŭ9���Y��:�!W����W��1�o�O��v)��I������^<}�t�錞GB��1 ( DI���	=��WN�N���o輨�����i5��~����.�	㚍��Zñ��B켼S���=~�_�)��+'�e,��yj�"!�[Fն3p�Q��c�������m�����# �$`�]�adÑ:�����/踠��c��]C���}�d_/_$%�s��!5��2�7W�\޹4�@��7}�;��X���>��h�h���b��i�I�JTl�U�S4SQ؊lg�H`�!�_�۞�'^?z�L=0UgP��]��Π�]���Ux�)�xhj���VFp��/F��� Ǌm����&���f,j���J9+i�����;�-	��'42DDDDDDDDDDDDD�p^�x�cǎ%�j����j�~=�97���*H�U�������������2eJ���A1DDDDDDDD�j�R0o��V !��Ǡ�7��_��1���3f1���t�4�'���b$(c��Q��I���W�A1�$��������J�a�����Kg��`ԜZ뺯C��et����AU�IH�����$<I�-�%��U��[����g�~�'`@���Ig{����Ǯ?p��	�ƕ"q-+O��59�9�L�2H�d!�h��o���kQ+O-��䘯N�:�{t��˔Ǥ�O��7c���ػ����?2!H @(A� �	((ME�HQDDEŵ��E]�u˪k��� XTT�4�]�PB-��>����>a�̄��0I���dfν�N�{�^r���vn����4���?y:T��+�&?�W�ےf�W�󓠘����� Z�WW5��=�>���k�ԻD�"\��ce�	�?d����<�{a�zy��:_�����\�����b�\�`4��q��y�L8(          �g�����ʒ/3�/..Ζ������*W�l�cr�d�|  ��#(     �3�=,��a�i�Z�k��CA�b��>G�Z-U�J=��u{���ďO���Z��9�)��Z+��(xP�E�5v�X�f鞥��q�nlw�}n.9�K��O{���Ѥ���~�>�u���v���Pw�$e�f&��,�r��adƦZ�Dț	�0�@��������!_)P��6p�zZV����(����z������սQw��K\��2��t���m�'�g�s.��ۀ��2צ�vt[��P����VkP�A.��7�o�P�d����+?�+�_�Ug>M�S��:��ݝ�v��w[�S�������5T^L@�?��S�Ӫ��������Y�u����=��Z!��4������s�;3D��         ����S���9�N�����Jpp���S�T�r:L�<>W�D @� (     ��f�Lg��CA�7��QVk;�cm�r�-v�jV�o��m�*T;�2�����ӾN{������#|�c?<�~��)4(�>�[��c�v�rf;]���������n��W�yU�v+���M�=� ���~t� b3xټ��g�?�SW>eǮ�0�y��І|���6(�
y�mnPIa�#�Z��Fw�vhm�m�=��������ym�x�b�n�ƶ7z<(�o��y�0.�������_�Ř ��U2h���z�����6��n�x����ye83�qx��n�1�3@A�y�z��Cy.��oo���C�����l�r��z�e�L@�'m34�~s"��U�Qކ������?��!          ��СC*�RSSm����UW�|ysfx�)9�9 �A1      n���2_˭?�^���t5pҝ�y�f`��#=�^͐��߼�~���ʲ&՛�sO���֣[���f��KV�P��#����h�����2b���Lp̄!t�w����{W�	�mX�X?�� ����m�߯;h�����ϟ��Sw^���F�q�k&��PB��I�����W5�	.��9ll����|��W��m]A�!��D�ۥSI���j�u��=�������<��_��3�s�=��IC��虣=�xS�����٥��{��ά���1�j7�=��Y�9�N�d9�|L�n�V7_|s�:s�=�� }��[_1���6�ۮ%QK�	�{�G�w�.{WO���|���vS)���os�&���m���v�u���i����w����<C�Mhj^��          <�ԩSJI���%Qff��=j�+�����cL�Q���W�n�d����� pn�      �Ѫv�|-g����nT�X]�z^�S�6�h���x��Ŵ����\P�3�}��-�T�S��kY�%A1�Y_��J�v�=]�9��y���~���=���R�J=u����,�S��BC�2��I�H�����q|�`o�b��n��0�3}��SMZ;I(��V���z��g��uq����й��R2Sl1!.e�LX������.���Ԅbَ	+y���z��'<Ҟ	Ÿ���n�g�9[I�I�$8xk�[5q�D��רZ#i5�m�	>ȯÉ���m�+#;��+_��3(Y>\�ˠ�&(&�c���Y@~���1W��s�~�@��zD�d�����lCa\y�����~J�����׏�kU�7�TY�_�|�˘�4          �'==�{�yHMM�%:::W�	�1�19!2�q��;�  ��     p�e͖�Z���b��)��f�vx�pO>��lT�Qo�{���ڰ���Y��ʄ��Kq�[�l-TP��[�����f5�ف�9���)��j�G+�Tv��1�/��ɏ���k���=K�{B����W���Cƻ�77����A��W{�_?�~�������kގy**��R��T�DT�p[w��g��Fw��V|��1;����W>mC�ܙ��;M�������y}��6���yfʺ)j��1���S����J�JJsmm��Z�n����W��7�]D;�����k��������2An�����g�̾�����o_�����i�z���k^s[����OV}"x�9�M�yj���l�fl�!          ��!1�fd:d�_9������R���@��ի+  @ ��     ��	��\��e:3���.��<t�y��e:(����ݍ^i����Q�O��,2�]>G^��=�h�����0(�|1��M8�o��v����/�ߞ�n��6ŧ����PQ\��n�p�Y��A�'$��>]��r�um�k��n~��"�G��1���"Ŕw��ÿPH`�<�B�
v�7]���uێn���p�{�`�V�Z��x���֛ ����I�P+��^��r�C���{]������6��1�|-ܵPW6��e���.�GC?����V�nY����W����S|��[Ŧ�
8�����g��LZ;Iws��v�{s񛺷˽r�9\�_���\�c��
����?h?Gݙ�q����UYuI�K����|�6����sX��y���-ߕ��        �Ad�H��@�ԬPS��� �&N�Sqqq�DEE�>c�	�1�29��,"(     ���U�k��'���n���BK����z��v@�7�m�W��w��}+Uִ��Z5*�8�r���0� Tm ��%�%��'}5��jS���������׈�F��Pۈ��z�T{^9�G�P�O�k`Mi������������$�A��N���m͍����vY7��P]��*;x�0��뛑ߨ[�n�43������ͦo���J�F�տ���v�g���/�Z�Pw}sW���U��_��EA�An�7���&,�B7��a���2�m����4��B���G��56�Ǖ�G���{��G����ڡ��p���q���ƂgL^7Y�^��0*X��G+?p.�������s�i�iԌQ^�l-�=�{���/t�%w��7�O3n��~��Sjfj���yaO�>�u��ΌBn�&����\���,s�)���SFLQ�{乜	-~qދ        %[��̿��X�� ��IMM�%:::W����BBBT�F����"c��w P     �BX����v��¨[�n��1�s?\�ʢ�!55�Q^k��8�p�uz��O"�3�=?�W�n��e�fva�X�\E@Ip4�z��C?��ᬀj�����x��z��g���m��ڀ��]G����[
��.׵�]��E���TO]���`�k�_��u;j큵y��k�z��7\֙s�w�}�����������חÿ<���h_��$z���zo�{��q�%*r�&���w�9\�N<�y;��� ���=2�;�>���7լQ��][s`���m&0����{k�[
�1�W���}��S�OѪ��
��6ެ�}ކ��3����h�;g��P-�]��rBs�ŷ(�?P1'c�IJOҔuSt�e��{��G�jٞe��h�G����s�o7���Fʙ픯3�~׷����i������'ߘ��+j9Ȇ���6w�]���ۮ��������ž/�����W�w/.t�]�
�tO�{�x��U�B�s.o��&�          ʺ��,����yV���Phh��1�1&8�<6�z��
 �T�      �P9�r��;�|\�%"4�������ʪg{=����^���u.�a4fpYҧi�|-g	Vk�mG��ێ%"(&�������qPuG�;N��W�O�v�׆!�_>^o/}�#禰�0�p��]V�b��������*x�	�zu�zo�{.��g�	��ـ<�1�	?o�Y���wYo�q�>�T//xY�,}��[y1��/Pc��
�+�UgBC�D�Q�f}�I�6Л׾iJL �7����m�u"�@�ԫRO��x�#yz���+ә)O0�'��v��fxqY����OOj���y���������1�+�]��/&��au+��P��]N?7���}�k�O����phC�뛰>zd���L���<��cEz�����.�����v�5[h��v ���ߴ���|v���K�]�������e�.cӀ��s��;s�G��������s���bBȾ���ez^�S�ߤ澠Ik')%3��r&�ĜwL V^3�E���^������{h�����.b�v?��@�����v��Ra�
��.��)'�p�Bm��h�̶ޢ}q�\�g~��j4��c�u��m��u��	>{���       ��0�Pk��Vx���!�f���q��}��d  W�N������}ς��Oǘb�dL�L�����FP     ��f����'�/(�q��^���ixS;��,i]��^��gg�K�SYP�r]���|/ogGPLfv����8|�	65}��D-��!�U1���РP=s�3z��6�c���Z�s��$�w�5*����Ѝ�nT�f�]k��8������|.x�	3�֕k�_c��޿:�v��a���Fu�#���<��	���g-߳\{b�(6%ֆ���m�!���juk��m�Ǆ�'hw�n���0a+�v������s����z;��<7��|5ǃ`]�J];�ڼ����y���,���)�����6!Kgj�Vs�k��f�9�~�N��A=��]'��<1Ǟ9�����н�A%�%�
��դ��?�^k�Ѽ���z�=�d��^X=�ߚ�U尿�>����,���m�9S��j�rFL�_���"�ǅ=l�pf�߻	�1a5f2�|�kSL8L���>d�P�L��	�2
�b΍��M��r�_>:o����P�bu�����/��ڙ!�e�L>���{��m`�G�����=כ�
�z.�X6i��ӓ�)��ʫQ�Fk/�?����|U�*T�mo��L朚��`�9ט���UաМ{���:{.       �|1��M?���&W�Pzw̽as�����`{w!�  �����DGG����WHH��1�1&8&'P�F�� �'>�      \�T9_�9��*���\״�F���VP�ۃ�v;���L���׿���ܤ�����������k4Wq(� ?3H�"�A�@IbB�Zd�3�xV�9�mq�-Ǝ�;���'v+:!Z)�)6TÄ �P�Z��ԸZc�dB�2k�,=<�a:�x��E�E��߭;c��k>�&�v�Z�翨�~>��*VҰ��l)��;������ݯ�b�[Vb�'�߯&ݠLg����2f�u����6욫��5�ѴH��mMX�pWFN���Tês�u��ɖ�x��l،'�����5���j�9�7���w��������+(fƦe&�p��o�a0& ./!�!�b�-eBI���zℂ3p����E���?���>6�       ���ܓ}����9���ץ~[̄6_��J���_ �/���R\\�-QQQ��M�Lxxx��<((H �m�      �`��GyGy�U���1��H�g�TV���W6��X�9��p��6[S�MQif���>Q
;�9�	�AId�Z}>�
~���l�WLǜ�v�qg���zqދ�9G�OV~���|J�.��7�K�]�U�W���?��ӆ�&�\~���0n��Tf����x��YzV��|1D�]�6��x��w����~xL�v,��$��|��bad��������+?�'�s��IC���Okl����v�zk�[
���r�ޗ��&'�%�aY����_���|����q����.%�'	        #�?�N���S�i��^ŀ���OtS��O�f���I�����@��k (ݒ��lq"|:8�$cdr�+WN PT��     p�ԩS�Z��_��%l�mD[��h���Uڙ���_��y���!�l�2�ݫ���6�8p�y��*���qf;�dfЮ)& ���wk`ˁn;DJf�f�1K��H�w/�OZV�^]������eLF�O��َ���e�-:�pH�t{�#7�M���P�zX��Ly�)��ګ����|�������1'c�}Bw�9C�/�]���~��O��^\�ݦ�޻L?��Q�k�.r{'RN莯�Џ�(o0���濤_#�;���e.��E���g�?<�.M\3Qc��v�-������(�LX�u_^�g{=��z=�@[�6l�0m=�U8?L8�#���?f
       �3}p�����.��}�����c�
ӯw��K�]����^�o��a�=^  J���T[���s�9�����c�cre���U�|�M P�     �B~?{j ֹ%(Ƹ��]z��T����\�*T;/ۯTYߎ�V=�'Uژ]̠Âj�T?��Y
����|Y�k�-�3̀�ԳqOuo����y<RK��hѮE��ϟ����}��=u�S6 ͕~���s��Z�oe��ϸ�~x̆��q�j\�q�ߓ$��̇�~��o�^���^�����_��]���S��b���z�gl JqHHKP�O��.��~/��s��`�;H��#�������~^��x��JWP&`h��i��O��E޶��Zu����B�p����m�H�v3y�d-ۻ,��(8�Y�WP��+?���|�8�E}��;�g�ԧi�B���/�����?�pfg{��'l8�	��������=má6n����       ���۴��g�޲�<�-�'k��f{,$�L/�}Q���:a
 �	� ���t*..Ζ�����L_�ʕ+��1A2g>
*x�- �A1      .�e��k�
T��h^��G]2J��Stb�J���>dj�O.��#&k�C�}*[���6Cպv��g:\X�B�8�C�T�r�B����*�4ILK��Sm1*T�� ��6Rx�p�<�`��P���ǵ'v�v��,�!W��_�!G9�7�7�\l��\���6R/��v����|�7k�,���']��z�������IG5w�\}��K�*�e<5�)����2mo��h��^V��*6��z��b~f.Բ��zB3}�t��7�}������n�n�x������:�3�t�3�6��HK�,����y��n���:�yzV�=6�Y����~�6��9�aUL`�����Cn��}�3miV����k�_c��
.g�����&��O|/k�u{ܬ;�N��<�t�]_�&jX��ۺ���PZ|��3-��:�+>-^�&�D��}i����5Y�Yn���`B@��ϣڐ�V�Z���w�ϾF��s=smh���l�FS�M�ǘ�Ŝ�9ￗc��
��9O�b΍�+VW׆]���\����^1�u��k�y�\�m9�E        �ӱnG���n���~���5�-���[����z��r �Wذ�x��o˞={r���1�J�*��d�c4�� (     ��)'�\�*�T�D�)��A�As�=<�a�FW4�B�x]�`H�!z���򥁈EU9�������@o���_�u�ғ�H�43�N7Eo����oo�W�Rx�3۩�f�b�l_�_d8�bfK�HQ\j� 0�w��ps�����i&(���ڒÜ�L�)5+մ�G��++�?оw�d޿	�1�&�W$�'�Y�L	S�:�l�I�J5b�1��q����Vpc�����Rf0���^�%"4�ș�Z�j�XI��L�=�>�[[�lՖ#[ι��/���U[���բf�`��{���1��2!5A������)�x�"�Ez%,� �� �9�ڢ�TR��ҿ����q��*-�gsIr �@�ڗ��iIz��`B����-&t�e����_5����6�t��dB�r>����d��%��b�nr��r���a�y�^X=U(_A�A���2�S^N`������o�S�ګ���       ��Ż���w=���\f������������6��3 �+VTbb��▚�jKtt�c����
�1��Ǧ@��Q     ���fЏ���A�fPQ�Z��܎�i�֒��7v�J�&՛�ۑߪ���|Ř+����z�7��)�׮yMu*�)����u֤���M�6(�:�w e���l�2[J
���:[J230~ѮE��TщѶ̉���ĄE�!S��L���V�����C���K�i��	�ۘ�Q�7
        o�դ���M@��m�=��'�k߰_�Ä؛>fb���t��i��{]���̋���L"��� J�ڵk�������[\	>cʙ�2�q~�� |A1      .D'D+?̌еBjٙ���cݎ	A1����>P�O���ӏw�������{���גӧi�"�ӹ~gy������ w   ��{�ܣ@�@�u&�g���         �ӏ��.vY7�Y�>���\��:u����}��;=7�9m;��e}ŀ����-z��+���;fb��W~,g�S ���ׯ���H%Ijj�-�ѹ�N��1��Ǖ+W&D�Q�      �����|/� ��W�b<�ѷY_�|���j�W*�̍�w�U���U&,���Ы_UIԤzM�eZ���ߺvk{��d�Iy�i�q��^� �9   �G�#@�_v��zf        @Yզv;a�+�m��c���~�ai��1����<�3��>Z�~���~��:\���rf���M�j��� _תU+͛7O�N�P����ȑ#�����Phh����N�ȘǦT�VM���'��}�      �p4���ӓU)��9�m_��V�[���ɠ���h�����W%UNHLǺ���l(&Lh����tf��
լ;f�9�K~����S�N�m�o�K�]b�QP�   ���퇫N�:.��S�5y�d         eѥ�.u�z\j���f�Ж���s����9Cb�d&���i?-p���̕am��D0�]t�"##�vN�Sqqq�DEE媯T����$��Ք�+
��     ��Iy�zt���g�R�����}�����<S�B5ͼ}�.������Q��f�9�D��丧�=j�D7L�A�)��u&$�����5�{���^��\^����*   ��G�=�n��%��0         �'�I�\Y��c����8R~���֯ڿJ/����O>�ۦ�f�bʕ+��~@�r�9��v
 |]�^��k�.��e��ɶ8p W����BBBN��T�R�t�L�5l=���     pc����
����e^{��5R���o�mD[}1��8�Fe��VIѪV+�8�G5��@%͕��Ԛ����i������W��i��sԩn'��۷i_��?N�P�cp��u  ���f��έ��-��         |��O���k=�����Y�ܯ�:�ež�z�׺��M��V��5[h��- _��]�j����ZVV����l���:����O���6@&'H&�)����7�b      ��o����Z+���$��{�׬���x�D�9��1��Y|}��

UIe��%�/ѫ_��^��,.�Ҹzc}��j]�����\����K��h�A�A����^/6%V{��
   ��d�3����6L���         �U�6t��ڃ�	�1}���n�~á��c^��1~�x�A1F�z�	�Pb���S111ںu� Lvv����mq�bŊ�Ccr�dr�� �      ��$jI���uQ/MY7�����A1�moS�#@#��TVv�|�y/�}QO�|B~��T�9��G�����h?�!����៫rPe������M{k���m�O�>�
2?�S�N	   �_��m(dDh��z���          ��*�(��U꺬[p�G�a&�2��ܙ�aj���b�
�ۧ�a�sյ��B PR�+WNC���˖- �9y�-�U�p8lXLN�L�*UN��T�^]��b      ���S����^�z�\vX�a�	.�+_!o3�sT�XM7u�bN�ȗ���RSFLQ��vi/1-��jb~��ߩ��x�zRz��jMBCl�Z��Wo��K���pA�B���b����/֌M3����no~��{�o���|��i�M����xP̰v�
�ނ�  ��a�;��t����S��z�ި��N̫������;         PVլT��m��Lg���<�m�{wy��qF��a&���c����\uM�7 �$��C�^�t�j�6ԂI�r:�����%**�:sL��� �5'D�<PZ     ���;�k�%�ι\�z�Jpŧ�{l�=/�
�+�8����6i����|�XI�\�������N�3���%QK�1z����B�g�������uQ/]}��
p-u܄j9H��M֛����c�U��b�a���_�V�Z�l�o���+��S�iτ)]���B�;o�<  �x4��\��)��Wtb�����         �����s%.5�c�]�wq[�+f��x�6Gov��	����aÆ���;�������� ���[rgdd�w�k��c�sfp̙�2&`�ۓ��DP     @f�13_A1&�Ą}|��K�m�_�~*NT�@��_��{]//xY'3N����[:ܢW����ЈB�a���8j������|�ؔX��?2���z[�^���V��!��h��#tŅW���f��ۥ��ڏ��OW}�9�s�l/��;:ݡ�]G��j�8ըTC�u��݋=Ҟ�ه�x�?�����  �o3���7۹         (�*Tt����{��w[�t�Ry�G�p���� %YHH�Z�l�.++�ɘ����X������5S�sOp-55Ֆ���\u�Æ��Ș ��P��ի+ �h���FP     @�Ĵ�|݀4��
�q�9t]��T��;�뙫��moӘ�c4u��b�����GꉞO�I�&�j#Ù�i����oj��-*&��՟�Һvk=��Q�h?�����n�L9�rB36ΰaE��./RpOp�`]��
���v�����;���Ʒ��   |����?�_��"         ��s�������h�g�����.O9�|���� (����O�N4j�(W��A2���JLL��1&TƼ������l���i�5S���r��>�M1A2&P&�qa'�
��     �<�g�۠br.=.�Nu;í5E���]�:���|1۞2b������[��&�����d�o�E����5�Q�R�Pmd������Ϲ�ԡ�C:_L8ͨ���/��>/����V�
�t�e�ْ��e�+s�}�����S;��A5iYi��1A?a�a�Q��Z�j��m�.���7+�� _0��P��9����9F��&/36�   |������6�         ���E�X�#�w��c��m�����\!(@Yvf��+&�"%%�t��)&H�<7%&&F�����DGG�3�oHH�=~Mx�	��Q�����U�re��~L�A1      ���O�c<��I�<��ۼ����j4ӄ�&h\�q�n�w���l��1W'3N�=?u����h|���V蠏K�,�#3��C��+��u�7wi��	zk�[�ya�"�i~n]�w��s����p;k�/1nhs�>_�y����/�z+����#[   �s0�>[�����}K>&          �_|j���CC<Ҿ�$ϝg��8�<%)=���f24�W�L� 8���A�DDD�\ƄX� ���d%&&� ��PSL= ����:}�EEE�Ug����гBdrB��U����@�AP     �9�0�mG��y���\���שQ�F�:�ªZ���(_R%����N[ҳҵ��jm9�E�o�?���8{#:9=�._9�����T;��.
�HM�7Q�ڭuY��<2�Ijf����	}���:uJ�hc�F]�ᕺ�˽z��7�Mlo)i3��q�E
����U�դW���x�� �(V�_��f?�ń5�����n����D
���z��#          �%�%�|��7,�(�Lgf���\���:31��7�)�r��;��r�r
 P8�����c�,���l�Ell��1�s^3�}�_6PR9�N�!2�9fs�cL1A2&P&�q�r��BP     @>�����9�s�9�J�Wt�������dCV|U���5�f������<�fP���͒~�@�v-ҔS���ԵAW�����.*���C�j�Ǔ�k��� �(LP�) �/:1Z�-zM          
�L���OլF3;�[a���m#ں�_h�<�B��Iגғ(  /���?FѨQ�\�&�"11�Z$''��&<Ƅʘ����- ����jKttt�:s̆���cքǘ���c8<<\�˗�.�b      �a��z���T�R�s.;��0}��s����oǯ����~���6�[�ݪ��T�$ۏm���/ק7|�[:ܢ��$���b��O^�u�����P�.{���;             ����Lg��;r6!/E	��\���qgٞe����._7�# ��q8�C(�1�&4&��@���$�8&&F�YYY������\����gǘ�*��3�     ȇ�������7._˿5�--ܹP΂����6׫E�Bn�.|U���L��1$=+]#��=�{�l�gmXJY6��P�AaS��|�Ӹzc��+3�̄�             %�3۩�w�e����4�)���-�Y�x�byR�*u]���FP �:LaJDD����  ��������A&P� �a�7S���s՝"cJ�*Ul�L��>��4 (      ��/�G�=��J��\�Y�f6���9��}?���!�Gg=������΄ܘ}�X�1�;��2�V��C��]��U�Z�b@E}���X�P�3AOq�q            ��h��ͮ�bZP���xe��l9�m���vr4Oj�������	 P��ɸ���e�bLpLll��1�<6��`��:�(�K�
�q8
��1&<����T�^]��#(      ��l/��|��?z�C+�����~����]v���l.��韟.!1g2�C���z��7T�]��J��d�&��x�e?����ݺP�9�tT�^�o            @I�8j�njS���$\w{X�,|��m�>\M�7q[�p�ByZ���._�<) @����:��Q�F��N�mx���c�dL��y���) �g�3sl���ބ=���� (�����     ��pŇ�ut�7Fs���ӔS��펊:���6�K}_�6n�8���U�Fo.~S!�!�{�J��o��}?����V�[�mG��]Ƅ.����_c�URz�             ���9���*W�\����zZ��Mҡ�Cj��W�=���f��:������Ƕ P�9�<�(�y��$$$ؐ�Մǘ�9�	��&55Ֆ���\uAAAjР��7o�6mڸ�.E� (     � 2��������_�|Xp�f�>SW}t��'w�L�����+��
�3k�,=7�9�f/�{A�j���m�WI�}*[��,ӂ��t�R�8�CG��*+;��PӠjum�U�[V��}��؄�̹k����]{c���g�)Lǵ5�tէ            ��lO��>�Z�ֻ4W��5�����~%�%䫽�/�Y�/���X�1N�Iu*�Q��.�"�G
 ����ȡ���ԭ[��2'O�t ���` (���4m߾ݖ�˗k�������A1      4'r�����[:ܒ��[�n����M�>�É�Ϫ3!1_������"��	�m�m6��43����P��բf�&f���v����w��Ɍ��zd�-�����m�k�r����V�����Ճ�?�o6#g�S?����1W�)�{5�5ws�m             J�W|�2(�h�V��_�۾�M��7��Έ�#�ٰ��\f����'�I�\1�m>�Y  UŊmq^����+<�̯��ɥ�;�	ǎ����C��iӦB�"(     ���1{�2�Rx��7! �����kîzw�j_���?��0�|�jR�%�'��w����(_u$�^^�>]��R3��ofz��`;��\����V����2Mo'�mhWo���"��7����             ����S��>���s�b�b�<�F�o�^36Ͱ�����W�O�Ck�~�wt�C=.��v2��zg�;���+&$&>5^  x[@@����mq��t*%%EIII�����������L��	��׌����ot�m��nݺB�!(     ��'ם3�Ԭ;f�\�r�Z�I�&��}q�lPF��ZBn�.|������?5n�8{�ט�s����/)1-�Hm}��+���5M͐����C�5v�X            @ia�s��=FSo��v���ݍ�������nyR��uԣ�뀚Ż  _�p8bKDDD��S�N)99نǘИ����P�dP�deeٰ�|�1�x     PH?������}=p�Z�~X}��mG���/�,29C�U��m�+�\���F� O1�4�am��[Nf�Ԉ)#���.             (M��������-z����$;������V9�.�D-  %��d6'H�nݺ.�IMM=+<Ƅ�$&&��9y����ߋ/��W_-�b      ��ɟ���/W��vŲ=�2o�<ܱ��eeg)%3E5+�T�*uբfui�E�j���_����#�)����L=:�Q-�w��~+rf;��q����i����7�J���|��"�G
             J�S�Ni��QZ��
5���������:�pУm�A�#;�tY�}*�� @�lK�Z�\�gee)))Ɇ�$''��������0���l%ɪU�ԵkW����J�h!      ��������W�F�^ن	��r�����؀�����\��z�k֯D��,߻\sw�UY�p�B-ڵHW4�⼽��IG5���x��D��ʏ�x��=����޵�             �V'RN���}��E�V�c��W_o�Z�vM�kԼfs�u��`�� PV���+,,�W�N��1�1&@&���9ń� ���[�l�%�\"x��     �q���i�C���*�(�Ѷ��n�h"�Gh���8�a��/�=]��=��Qx�p���s�
�s�>�e.;/�^�o�ݗ�����w�����>��cf��z�χ�             ����G]���n�N]�w)R[�N�ҿ��K/�{A����ϻ��vӷ  ��p8T�J[��w������8%''+11�ɘ�9���m׮]��b      <`鞥��n�F]2�cm�٩��w����Ej�`�A>�ڢ�4���z���Z��|��C�m����(&���7���s��w(-+�X�w ��~��G]��:�����(+�t|             e�����>��������U	�R�6v���?>�Y[g��7�Nu;��35�o�^  �`���mq'--͆�$$$��z��I�v��{}W�\9���     �������t�4��!1gJNO�+_�+>п��K�_v�~���V}&�ϧ�>-֠�q���9��?����屠���1��C             P��ɵ^��u����N����]D;���s���h�<NY?E��N��]�_��ۺ��W���  �g�V�Z���t:������8%''��&@&66־fe���Djj�RRRT�bE��1���b      <džk��e�jc�FyC|j����&�����~�K�]��)53US7L�gƦz{��
	��vL0̘�cl'��a���JLKThPh��Z�oe��             ���K��[K޲�Z�jj_��Wo��A�U1��bSb���h��*%3���)�?P������  ����PXX�-���SL�LRR�}���UZ�b���	�     (��nCX�W)R;&8��/��L���/�SW>eg�(�(��������'9=Y?l�A7_|�׶aBUF��	�'�|1��,ڽH�Z*r[ff             �t"���o��d�����   
'88ؖ����'O�T||�r}5�͠�)EB~�a�      xH��l�ڿJ}��)R;S7L-�����,�4�%���͸u�Uk��67r����s���v��o����u���1�#A1+��                ��*V�hK�:u\�gee)))Iqqq���Urr�-�ÿ́ʘ�OA1      �bߊ"�|���uש��5�I�b@�n��B\3:���ʕ�h�&h䴑��a�|��]��܆	�Ys`�                 矿�����li�(���N�S���6<�|�	�1A2&`�<������     ����^���%;o�q�q��@���=��Y���u"J{b��I:��G��U�Vk����j����|��cە���J��
���Û���$                ��s8��d�IMM�29ńʘ��ĉJOOP     �AK��)�b����>����ԩSz~���}b�>��c8���-G���q���<��}*$�0�����ְ[���y��                �����DDD��7A29�1�������!2�)�#�6�      xPzV��휧!��j�u��|��K�?��w�TH`�׶���6��?��鱶���W|(_�9zs��bfo�-                @ّ$�F����ʲ�1&<�ɘPS�c�A2(��     ���.tP̦�M�w-��]�_��Ea�a^���c��<3a��k޿�v��]�u�'ת��                @�����*Hf���v�����'O�`$c�&$$(##C��!(     ��fo���S��+�W�u�NDɗ� �+>�B��J�o�P�!��É���ƌM3��̇�ˊ�����g{�                �_���P�V-5l�P*TP����W��i�dLxLLL����l�LZZ���FP     ��I:�uשS�NZϤPG'F��l�ޤ�����*,8̣m'g$�%�%i����֩��|�ʾ�}�^�3                �	��������7Vpp�U�jU5j�H��???egg�����d�Ή'l�LRR�}nƊ �DP     ���cf��b����._�1z��~�W�РP�����$���Z����t����̐�;�r�P�e�iN�                PL�KVV�-9ʕ+���[�֭k�� ��	�9r�v�ޭ��%$$��>P�      x����K}_��˯��4����Wk����]�*���6S2R�R2��1�C7L�A1'cTĦ�j���VbZ�              (I���T�Y�@�TtT  (�&�ؒ#55ՆƘ�h�"egg��b      � �D�VX�K�]��uҝ��u�v-Ҩ�4���
�q�b 7-�R)�R��{j�SZ��J��'���(p �	d            ���[�n�b�����tf�h�QM>j�Mn9�Em����Bޚ�4U��zZ'44T  ����Z�j�����      /�z��
��+秒��_�~X}��7��m�q�2/���,ݳT�.{W%��0P�����$��6[         ���;����?���� E�}�ZQQ����.W��^�.�k���^[�����jk{���*j�D�wqd	$�$�,��NO������L��p���w��y�O{f&�  �3��%6�id����c�?���a&]�  2�P   �Z2z���;WFvVv��w�����~�n�k��᫵OQ~Q��J
JZ5�zYu�:��hlj�L���Ԫ��M�/j��         �����1���o�o�~+~��c��1���  �eB1    k������G�ƾ�m���y]#S$o֞zש�Sߝ�_i�UާoI���-m����'.M_�%�6n���         h߶�`����w�+����>%����   V�P   �Z4�͑-����GIAIT�VD&(�.���~<}�ӑJ�Vi����*�j[�޲�s�@���}d���K-�^ONy2         ����=�8��8c�q�k7  �j�b    ֢{޺'�t�"/;�E������9��I<��3q��7��=����-�ky�3jMH���uu��
s[��g�=��aY         �9
r
�cnJV��O�:  ���   X��,�'>x"��շ[4�oI�xg�;�I.x����oÒ[�v�>�_��ߟq�����=�����U�GM         d�K�]5q���  �:B1    k��7G�8�E�-���LRQ[>ra�v�m�^ۧ�Ol��V������_i��kP�����_F&�ѥG��Ϊ��~�l         t&sω�'��A��.�%�K�?��q��#+�ժ=�>��x�7��� @gWPPK�,	h	�   ���w��e��7EWf����Lt�;�?����ӆ;�z큃�Y�7?�E��N�O>2�&=6i�ܻ&��M�        ЙL�5)�w���=J>��z[ƶl: ������k�dge����[��*�K �άw��1}���   X˪�V���&�^��ҹ۬�Md�$�q����S�?���6x���:h�Z4��'.�L׿G��}a�        @���^������[ґ�C�>4~���b����uw�8�������� @g֥��/L̈́b    ��;��ӢP̎��9���~id�q���sӟ����ݪuC���֏9���Խ�{��!+��������L�i�M[<w���        @���nI�|sd��8:���q��.����=��q�sפ/� �Y��P   @xg�;-�W�S;��9^��bd��>��������d��I��W<}E�O'�|B����\����l�g�ͫYV�L         ڿƦƸꙫ⽹��}'߷�XLIAI��N�׿t}  tVYYY-%   �&Ϟ��{��;cC1���hL�lB��N�Zw��ƈ�#���)����n��tά�Yq�[�D�K�R�Sߖ�{y��w���!         ����H�s�9�����O���  h!�   �6����xW<}Ed��^�.�����j����q�GƘ��Dgw���}�_�[^�%�5,�L���vo�ܷ�         d��_�>��������c{n�g���3T/  ��	�    ���3�g�&=6Y�ܽ��%%QQ[�hԛ���\����ZwɁ��}��Ʀ��R�T\:��ͽ��ۢ#H��o�W>y%         �<MMMq铗���c��XvVv: s���  ���b    ��S����8m��r�s�-��GG&�^V��q{����[�n����cw86���ߣ�:l��b׍v]鼗>~)>��At�lyH��>9��          3��6.fUΊ>�}���N}w� ��   h#I�%���w��nƆbwL��ա�Ĉo����{8*j+����5���U-�;��Q��e�Ű͇�h����1m��          3555�����;��Ƕ�`�   VN(   ��$W�hhl������Vߎ��ca���D��|-��ߣ��mX�a���ŏ��(:�K�]���t��7�������l�(.(n��$�        @f{z��+�lT�Q   +'   �Fʫ��O߈���ҹ9��׿t}d�$frפ��}/h���{��G���Y��q���h��&�'�>����]On��'�<         d�)��xr�9  `�b    �И�cZ�I���)�I<��C��I�R1򄑱��w�Y�����խW�>qtdge�h���>A�.=�m�j�ܪ�U���         �mA��/.(  `�b    �Н����EQ�$(���{����(y��QRP������tO��k���*'+'F�0:���k񚧧=�I���9�-����X         �m���b��#+��M�  |5�   �6�Y�g1v������?g�s26S�X㦍�#�9b����q��7�F� �����I�Rq���ƾ�m�e5��'�D�+�)�s�yn������        @櫭�]���3u�E��b  ���    ���^��š���=*����O}�蹏�[�PL�]N���8�3;\,f�!#�G{��Uk�h�����钿wߒ�-�;�|F<��3        @��ѥ�
�746Ĳ�e  |=�   �6v���Gyu�W���E�ٹ�����9=2ѫ����{$Q��
"�=x^���\:���ɐ��z�k3_�LW�_�wa�����-���
1         �W}v�zYu   +'   �ƒ73����.n��Sv;%F�-�(2͛��������z/C���s�oI�8i�IQ��&2U�}��a�3��J��g������^�z�h%���         t���^��Us  X9�   �u��箍���-��J��f��EC/�SF��&��|���ؼ�櫽���oG�rD�_2?2Miai����c�������Y#���>�������Ƽ�y        @ǰ��{�����>  `�b    ց��������9�E�O��=qt<���i>��fB1�o��FL8wB�4�xz�ӑ)��d����;�����GCcCL�?-2U׼�q��n��TV���5��U�
         :�!�Y���t  ��	�    �#W?su���Q�[�ҹI\��co���!�,��dM�y�Q�F1v�ظꙫ�G/JEګ��ܸ������.�����kV嬨o��L��G�wl�s�Ͽ��[��
W�        �(�v����������   VN(   `I�W��2���j����֋�'������Ɔ���sMK�9�9?������?��'���ЁC��C��m7�v����#S�h��	;������.�_>��         ��8}��#/;o���:��   VN(   `�ݸ��ɻ��nԢ�C6?�����'����b��=�l@�u�]���Oƅ�\o|�F�k�m�]��[��om��5��ܪ���v�h�����o՚��^�+g         ��E���]����U͋�g�  ��	�    �C�˪��4F�0��k.9�2oJ��8:2���Ek�: =�MW��2��hjj��4t���ɐ�ā��T*���_R�$2M�.=�!������:j���?         Cnvn�s�%%+|��w�Ʀ�   VN(   `=it���i��}[4?���r�-��O�/D{זo��7`��HB:#��&���羿��7�l`��1q܎��V�mkSu]ud����x������Z���G�5�         ��[~�����=�l6�+����  ��P   �:�����uJL��(.(nњ�������^�+�Ο�Y^v^��sP�A����fM���>�|�L<?��(�._�}���|��7⛛~3�;m�S��L�ZJvVv��/�7ܪuɛ����X         ���⠸��k�e�*/}�R���+  ��P   @;0�|F��s��cnn񚲮e1�G�b���׮c1���������>=~�Ϗӱ�|S�M�)��G>��UuUQ��*��-��y]�K^�(�/�^]{�f=7�e�����$��.$�'S\w�uq�և�jM�s9���        ��շ�o��1q�NǷ�bl?{�g  ��P   @;q�k��w��N��-^���:����X��>��hÒ���Je�c/������$���ޥR����1|��Z������t�        �/��΍ny����H_<.� [򙶒����j��b�������:�Zo��g�Z��o�g?z6  ���   hG������l��ܬ�k��I�b�^?4ޙ�N�7�t�$X}�)��"�Y���#���qZ�����_ċ3^         Vl���c��Xt��O���?;  �hhhh)�   �v���<���x���(�����/Z?^<��8�������d��	Vߖ�m���JcSc�7ɕjn;�8v�c[�v��Q1b��         �s��d~�C���2  ����	h)�   �v��9o�I#O�1'��T*��u������>�Ӹ����=�ѥG��g�`�u�����,�Ο�I�.=cԉ�b����^��goƩ�O����         ��^>=�s�wbʼ) �?UWW��P   @;t���Ņ�\�;�w�Z���W}�إ�.qƽgĢ�E�.0��Jek��[S�o?��7�1�=��ؤ�&�^;s��8��âz��        :���}(N��Ԙ[57  �_s���G��P   @;u��WD�.��}/h���v<.�'�:9���t�+���9�osx\�������I������^;�j^p��X         ����qѣ����{  �euuu-%   Ў]�ȅQZP��l}p�_i�;|l��ſ�ŏ_���іv�p��ِ`��g�}b�����缽ΞC��>�@̡[�J�+k+����}         t\/�x!n|�Ƹs��aY   �O(   �kjj�3�=#R�T���i�^��ʊ3���xl\���q���GCcC�m9Y9�ף��~ެ9���a��Q����N~���zJ\��+���t��XX�0��x��7        ��#���G��?�����)O�G>
  `��   h����1�Geme�d�OVi��]z�uG^��}N�xzD����Q�PkKٹ����w�6Gı;�&�j�s0���!���6�i���|��1��bҬI        @�3�~��h/���U.�����]9;>Y�IT-�
Zfi�Ҩ�k��+'ׯ     ��+m������fa\v�e�J�Vi�A�ō߻1.vI\��u�`̧���癗���Ĝ�����#���t�M1s��xa�k�\C6���:p�j�3�|z�aXL�?5         h��~7�|C�1�����h�
7�S��  ��P   @����c��iq�7G��.��φ%��ߺ<.;��7m\��8:���d|���Uگ{a�8n�����46�q�w�˪c^ռ�Mj��Dm}���_%%��ʊ��z�G~N~�k���1���q��+�7O�f�^��[~�8~����gŶl���=7��8�֣��o            V�P   @��k�]�Q�Gq�����/�#	�84=S�M��?�gO��f����Y<'��-Y�&	��-��{��7�=��x�����"��Es��ƄO'��>H�=��'�>Y�hI�.=b����c���6�o�m�]z���+�JNVN�l����=�ǟ_�s���m�ߪ�٥g|k�oő��6�Ѭ	{�oqƘ3���.            X=B1    ����ǎ��1n=��8x���ؾ�zJ���fYM,kX���-�Y��|5�����&Ifm(�.O�w?�K�%�m7�6o28����m��";+;֦���C��s�������x{��1oɼt'��%!�$ԧ�Ol�}�ش禱�;���v��{m�Tj�=�$,t�}g�-��           �?566Fuuu��Ԥ�&#9-%   ��� �!;$��缸���!���0�0=ړ$���{���>/~�b446��s�I�'�<�z�WQZX��/t@:�q������Zo��X�&͚��ql�?��           �� �xkVVV�k}}}��եc0�/�y���g�}�<������b    2X����㯌G�4�������v�����1�8>Ƽ5&y���Q>#ڻE5������G�b��M�	;���t|�EGR�P�?uyz,kX           ������I�$�D`�.]����dɒX�pa̟??�Ν����6	�    t ��y'�ip�5���Ձ������(>��,nx�����[��G�J�>�O>=~��O��]N���J�E�{��g���ώɳ'           d�����ڵk��0I�%	�TWW�{��/Na-Z��� X��b    :��Ɔ��k��	wƥ�.������΍L����c��#b���Q�PIeme\���q�����=��/�e���#2ʹ����G.�{޺'           �=�������t��{���Leee̞=;},��	�    t0�̏3�=#F��wa����-�[d���f�ŏ_��~[465FG��~i:sפ��/G�%������}?�x����;���>           `]KB0.L�� L���ҥK2�P   @5�|F�gx���y���?���1x���^555�/��?t~,^ڹ*�sω#o=2.zQ\r�%�J���I~&c�wL�#�M��y          @[hhh������,Z�(�����***���.���   �ખV�-�ݒg�uF\u�UQ�S�I�����;�-���謒�ʯ��u����%�.�������1w-�(           `M���_���������!��X�ill��b    :�?���x��c�c@ـh�������~�j�뱿��������^�O%�����>��XZ�4           `U|1��_�Lr��Xr?�;���b    :�	�M����s�x�q��G��'�:I$���G<=b��b�,�SF���}_           �ש��I_������2~I�'�9�>�   �N���2�w���ψ��:�s����x��������j]�s��{Ǳ1�|z           й%DMB/��K�5	�|1S__��'   Љ���?����O����ox����r�s��y��y�������.           �����:�I�/�H0����c��e˖|�.]�DG�J���   ��&|6!v���q�a��ɻ�ܦ�2oJ�e;�١��9�rv����#�=           t�����/����ͣ��"�I.<
����0:��hǄb    ��������?��G\���w��mr�n�݂/;~����|wM�+�sF,�^           d�$��^�Lyyy: ��N�%#�/��TZZ��R��hǄb    X����g������#�9b���[[|+^����,Gowt��+	Ü}��1�͑          @��dɒt�%��������R�~���!   ���[57����8r�#�G�1��Yk����ꙫ���"����ٹk�<wN�3�}�ܘW5/           Xwjjjb��GUUU,^�8}{���QWWОm��VA��   `��|o<5����+�=N�T*���ѻ[��������"N���8|����9f�ψ���x���          �����!***bѢE��H0�ǒ L22UQQQ4(hB1    |��ڊ8}��q���5�_�n��?Ǚ{���x<��Cљm�k���\k��,�����*~7�w��nI           �����ӱ�$�R^^UUU��N�%1������j�}������m�    �R/}�R�q���]��|ylP���;�J�m��{^�g|0��ʺ��C�>%%ke��'��?t~|���           ��jjj���"=��/����ɨ���6�`��y睃�#   @�465�-��c��{A���9�-��ٻ{a�xb�1����ӊO�3)�/�Ny �X�{'���=��x��g          �/KB0I ���jy &�����򨭭��
�裏N_@��#   @�,^�8.z좸��k���3�:#
sW{�~�����O���ib1Ih�>{n���w�g���.���{8           :�����񗊊�����OF}}} �STT�w\���#h[B1    ��yU��'�$�~��p���N�.�]Vk�-zoϝ�\�~h|�����zv������L�51.{Y�;���           Yyi�|1�|;��466��4(���oGqqq���b    X-�*g����=zQ����q���cÒWy�Mzl/�����۾�|�LtD�{�G���ؼ��kd�f�W��"z�!�          �è��KG_.\�<���(LUU��P�Z�a�w�m�Ql��ѷo�`��   `�����k��&���8q���o��n��*�Uֵ,�����1��-���ЁC������խ�j�S��:FO���1y��           �4555����ŋ���<I�0��d$��``����^��ѣG����o'���,����C(   �5���6���_�c�~�ǩ����pl��j��������c�M����;+��-�L�J�����<.9����^�}&|6!������	w��<           �U�I�/�h�4�O�0����}�����/�Hb0I��v�;d�    ֚W>y%=��ǹq��ĕ߹2�vo�'�zr�����ߏ�f�����q�17Ő͆����@\��%�P          @{��L2-Z���$c���QWW@�XQf��֋^�zEAAA�1�    ��-�[7�zS�5��x�'����U��E�t�Kq�s��=�_Q��:2AV*+��9<�8�(�/Z�}F�92Nyb446          @[hhh���ʨ��Jm�����oWTTDccc m#'''�����=z�C0�Q�$���t|B1    ���g��p`<q����dgeǏ��q��q���=o�MMM�^��o����]6�e��5q�H          �������ŋ�ї$��D`���ǒ���3��.��$#��$Q��۩T*�܄b    hS��|-������>������{�N�+^��B�������/E{2�l@\|��q�N'���7�rc�>�t�          ��jjj���*~i�$�d$ǒǄ`�meggGqqq:��`��Ks�gϞ����u�b    hso~�f�}����i���/�b�&��ų_���>�?uy��6.֥�e����<N�����Z��ݮx������          �P�i�4a��'a���� �^NNN-�����+=��%%%������b    X'�Ο��48�?��ح�n�����O��g�7�|C��8*/]m!+��6g>+�����U�X������^�.          �Ω��!����%��hѢ��d̟??���X7
���QZZ���4�N�Rk�P    �����1�/C��cn�cv8f���e�]���C���ߺ;�|_��:6j��Ě��X��F��w��n��ѱq����ދj�1�OLy"          ��+	�TVV�0UUU��I���<}���"X7������8~I0I��9
SVVyyy�P    �Tr9���b�g�7�&r�V�%�n����� =��U��)c�ُ��W?y5�������Je�������{�77�f�;`��[�7ִ�f�G�vtL�7%          ��V__�/NG_��K�I�7K�755��.��$#��$Q���Ʌf���   `�K����xi�K1򄑱aɆkd�.�]�ЭM�D}c}L/��,�$>Y�I̭�u�u��n�?��u�����^�=zu���ŀ��ck�M��g�wV:�          d�����>}z̜93����HG`jkkX���KIII:���/�`�QPP�i�b    h7���\ls�6q�!W�i{������ʉ�eӣ=�W5/~t�b�[c          ���/��ҥKX7���_��In'����쀎D(   �veQ͢~��7m\\s�5�^�z����=q�g�ܪ�          d�����뮻b����}ݺu[a&]�v�L�b    h�FO��x\2�8s�3#;�cT�?\�a�������H           ����!F��q kFvvv/����.��E^^^ �$   @���fQ�s�9q�+7Ư�U���J�"-�^�}�q��Em}m           ���G��UPPP���4`��0�ג����]hkB1    �{�gO��n=*��}:s�ևe̋�kƟ��S\�����          ��f͚o��F +VXX�/!������ �O(   ��1i֤8�#b�w��� �����ɏ�hʼ)q��7��⥋          �lcǎ������*'''|I�/��b&��<�]�+    ��ٛq��FIAI��aq��'����T*�N�WEmE<��q���SӞ�&          t.��ӧtt�����K���1�u��}��b    �XI�%��$c����c�?&����o����k���iŧ1n�x��G�o�#j�k          �X&O��B�tYYYQRR�<�D`�C0�������   �Cx����WO�*=��u�o��F�;`����ؼ��ѫ[��>G]C]|�ࣘ8kb��p|:3u��           :��3gd����(**Z�)--]��ݻw�q 3��   �gIݒx���ӣY���1���X606�i:&���%��u���Xְ,��VŢ�EQ]W��g��9���ySc�����          @�2k֬���!��L��]��1	�    �),�Y�~�jz           �TSSS��������(..^�)--]�)++���� :�               �
uuu�����.��$1�� L�5�ĤR� �"�               �
"1��/�`����իW@k�                �����t�%��$�$��Ib0������                |������d$1�$
�|;�J@[�               :����())I�_� Li��$�

�=�               :����(**�R�w��ѳg�t,���               2^aaa:��<�L�i��J� �	�                �^vvv��/I &��4Ga���"/// :2�               �](,,\IF�I�0ͷS�T tVB1               @���1�޽{GYYY:SPP ��P               |�����urss�ї�Lr���t����� ���b               �+����&��*,,\�IFs��v*�
 �,�               �]�v�����L�8N|�b�9����� �m	�               ���h���wމ�&'''�����޽{GYY��LIIIdee �P               |����gd(&�J-�$��L�����  s�               ���n��b�رQ[[�Mvvv/�����.�����E^^^ �1�               ��Hb+{�G�?~���K�.��/I拷���"�J �P               ���{�|�A̞={�������������FAAA �P               �Dvvv�p�	q��ǜ9sZ�>'''����% ���ݻw�q �:��               Z�k׮q�)��s�=���j,]��_OB0I &	�4�`�o'k`u�               @���������o̙3'#???���� X[�b               ������O�> mE(                ���                h�b                 �9�                �vN(                ���                h�b                 �9�             ����݆Jv���3�qf�I�E��Z��(V�|�����Kɦ.jC[(�鋢/��R�j�m��aq�!�I��c6�4�<h�n��&1���n��y�Ng.�U�Iv����|��̙��������  '                �8�                ��	�                 $N(                 qB1                 ��                H�P                @�b                 '                �8�                ��	�                 $N(                 qB1                 ��                H�P                @�b                 '                �8�                ��<�~����U*��fB1                @)�������3��2�z=��P                P
�f3:�Nt�ݟ\˲,VVVvb1�L(                �6�Y����/V*��ꪫ�ӧO/���׆�)��߿���ػ܄�~3&                L�޻���/��                �M妛n���q��T���j�����{�ޓY���Ї>�dL�                `������O]�����#��N�V�0<��Z�~�^��:�~���~$F(                �9��`4�^��×���q�R�7�x��z��sssy�С�F�b                 ~���g����8���7�x����ڿ����ַnM�{	�                 <��`?��|tcc��o����]s�52�`�P                �elooׇ��'O�<t��я>|���r}�              (�,ˢV�E�� 0M���n��� R��t�/\��w7�t�\}��o>p���^�+              %2
�,..���\  L�Q,fcc#��~�f�Y]]}��;>v���߾�뾵�k
�              @IT*�h4��y  L�Z��f3���v�1)���j�z��;��믿���\K(              J ˲X^^� J��=�ŋ���G�z�^����w=z��>|�n�#              %����J%  �f�YZZډŤ���W�����[^~�����XC(              ��h����\  �U�Z݉����HU��i\�x�߆�oߍ��b              `ʍ6M�b1  eV�ՒŌ�������㯻����B1              0�F� ����<R7bss���o��B1              0劢  Ұ���;��rK�����q�+              S��� @�M�=O��˷���hx���W(              ��h��`0�<� �����O·�=[����Xů�z�������P�������              ~���f,-- @moo��~J��n��K/�9��߿���s�t:������t��_��B1              P����z=j�Z  �I�ߏ�����̑#GF�ύƱc�^1�'��J��K�E�3~�(>�|�G�R�槯]�~�8��9#�{�śo���~���cL�b              �$���byyY, (�Qxeuu�Yc.����lxx��������U�^��N'�<����q�+              %1�@=�H]��c~~>�Uۉ��4
�loo����K��������xx�K��F�`?��?�y              (�N��3�,�J��s ����`0�c��xOL�����O(              ��]���=̖z�~㇣�U��3�.��'.<�����CO= �������Ȋq�{���`0����
�E�+�O(              ��[�[�5�-�v|�?���iT��]�i�����=(�[/���q$���Lj�,���s>�                �����EQ\��/|a��|��8��                J���?\�T&���������8��                J��}���o��3<�Ob��(�b                 �O�e�m��������
׌k"�                ���ĄB1Y��b\s	�                 �Uř,�&��Ҹ��                J+˲��Z;���q�%                ���I-\�Ҹ��                J+˲��(&��P                ��E�>���b                 .g�ɲl"k��                ��<��s0�ᄖ�Ѹ&�                J������S1�b                 '                �8�                ��	�                 $N(                 qB1                 ��                H�P                @�b                 '                �8�                ��	�                 $N(               1�۫����W `D(               1�A7y�xU�U 0"              ���|�3���D  ��               $��7��o�!^}ի @(               A�A/����/}�K�\h 0ۄb               uv�l���;����xY�e �.�              ��=r�����g���x�k�Y� 0{�b               ��ߊC�z(^������q�+����zt����  �O(              `J<p�8�/#˲X�.�Fw��l�ڈ��RL�(t \�              �)Sŋ�Č��Vw 0��b                 '                �8�                ��	�                 $N(   �	sO�E  �H�NU7�         �l�   J��F4��  �\ν�\���          �B1   @��?6��Db            ��&   �V�b5Zw�"�             �jB1   @)�<�w�#�f            0�b   ��)"Z_mEuͣ            ��   J�y_3��            ���   Je��B,�Z            �2�   J�v�+��            @��    ��o���r;�^             e#   L��Ȣ}W;*�             (#�   `���ھ���            @Y	�    Sm��K���b             ��P   0��O֣���             (;�   `*U�+�>юl�            @�	�    S'�g;��|+            �Y    L��{V�v�             �B(   �*�'�c��            0K�b   ��1wf.�6            `��    S��Z��]��"             f�P   ����E��v��<             f�P   ��"���VT��            �]vX   Ik<؈��            �,�   �5��|4N6            `�	�    I�=U��ݭ             @(   HP�ɣug+�^             �    �D�N����            �%v\   I�w���{b.             �B1   @2��K��            ��%   $�v�+��             �$   L\��G��vd�,             x&�   `��"��W�Q٨             �N(   ��}����z             �܄b   ��Y:���Y             ��P   0�s�h��             .O(   �s��J�O�#d            ��	�    {*�g;��|;             ^�   `O�ܽ��             ���   �L�d#Y             ^�   `O̝��ƃ�             ���   v]�b5Zw�"�             �%�   vU�͢}�y7             ^�   `�������G             W�.-   `�4l����            ���   v����|r9             �rB1   ��՞�E��V             0B1   �X��y��lG��            ���   �&+�h�hEe�             ��P   06ͯ7c��\             0^B1   �X,~o1���             ��P   p��?�Ǿ��             ��   ��T�*�:ъl�             �C(   xɲ~�;ZQ٬             �G(   x��}m_���            ��%   �$˧�c�            ���   ^���sѼ�             ��b��Y��۠�fw3  �r��W�����?             �#B1Dc�y��[o�� ���zY��hG���H            ��$   �`+w�D��Z             ���b   ����F,<�             �=�v�������J����;q��  �|���	�             0B1����?o�շ\�3��?��   ʥz�+w�D            ���    �)��Ѿ�y7             &G(   xvED뫭��y|             0ivz   Ϫy3��             &O(   x�������              B1   �Ϩ]��ʽ+            @:�b�sk�b��p��E?ή�  `z�[y��܎��             ��!���0;�O  �Tʊ,�w���Q	             �"   �h�ی��z             ��    �^���,             i�  �W�ͯ7            �t	�   ���W�}��              �%   3*�gѾ��V             �M(   f��=+Q�Q-             H�P   ̠��Y���/             �A(   f��ٹh>�             ��P   ̐�j5Z'ZE             0E�b   `Fd�,�w�#��            �t�  �Ѻ�է=
             �Fv�  �h<؈�G�            ��$   %7
�4j             �K(   J�z��{Z            �t�  ���;y��hG��            ��&   %���KQ]�?            @�-   e5             JB(                 qB1                 ��                H�P                @�b                 '                �8�                ��	�                 $N(                 qB1                 ��          `O->���� ��Yg�w6   ��	�           ���AY/ `����   0-�b                 '                �8�                ��	�                 $N(                 qB1                 ��                H�P                @�b                 '                �8�                ��	�                 $N(                 qB1                 ��                H�P                @�b                 '                �8�                ��	�                 $N(        ��c�nB��������ή%K��H��đ�(k�"BsU�Cq��=de�=$��D/S��Ň
���KC_�\�^JEӀc� e�4���tf��M��2�������`��{����
       HN(                 9�                ��b                 ��                HN(                 9�                ��b                 ��                HN(                 9�                ��b                 ��                HN(                 9�                ��b                 ��                HN(                 9�                ��b                 ��                HN(                 9�                ��b                 ��                HN(                 9�                ��b                 ��                HN(                 9�                ��b                 ��                HN(                 9�                ��b                 ��                HN(                 9�                ��b                 ��                HN(                 9�                ��b                 ��                HN(                 9�                ��b                 ��                HN(                 9�                ��b                 ��                HN(                 9�                ��b                 ��                HN(                 9�                ��b                 ��                HN(                 9�                ��b                 ��                HN(                 9�                ��b                 ��                HN(                 9�                ��b                 ��                HN(                 9�                ��b                 ��                HN(                 9�                ��b                 ��a�������Z���<�������7�                ��P{n߽?i�$�Amw����                `��b                 ��                HN(                 9�                ��b                 ��                HN(                 9�                ��b                 ��                HN(                 9�                ��b                 ��                HN(                 9�                ��b                 ��                HN(                 9�                ��b                 ��                HN(                 9�                ��b                 ��                HN(                 9�                ��b                 ��                HN(                 9�                ��b                 ��                HN(                 9�                ��b                 ��                HN(                 9�                ��b                 ��                HN(                 9�                ��b                 ��                HN(                 9�                ��b                 ��                HN(                 9�                ��b                 ��                HN(                 9�                ��b                 ��                HN(                 9�                ��b�Wt�ƍ��؈y����V�w ��c               0W�b�W��K/�͛7���b�                sG(                 9�                ��b                 ��                HN(                 9�                ��b                 ��                Hn�C1�$��fp�х��=Z{4���1�~��A��               `��:���_�����<����{��sq��.�4�¿|!ֻ�               �_s�                �B1                 �	�                 $7ס�����(6�{vvv�}O76�����                �0�:��v�����z�������?�eY               ��1ס                �i                 ��P              ����X,c����ȮSvb�� ���              �O՟��4?���cii)���c|{����_ ��	�               $�TY�k���#�G"� �!�              ��N�N����(zE  �K(               ����qu�j}� �wB1               	U�j�-�E1� �b               R�P���  #B1               	]�] ���b               �9T��� p�P              @2ã  �	�                 $'                ��P                @rB1                 �	�                 $'                ��P                @rB1                 �	�                 $'                ��P                @rB1                 ��u(������NpO��Ȯ��zn              �}{뭷��T*�LbvY�߻r��gǱ�\�b�׷������S�Nd����nM�s;               �!)��ceY>1���k���                 ��(�VY��=��=���b                ��U�ek���b                 ~��(ZeYNj�P�8|���X�S�˸2< ���7{7c���v                �`0x�(������Zs��տ��~����v���               ��(��㓚]����֚�P                0�>:��EQ��ZB1                �,;1��eY~\k	�                 3�wީw:�G'5�(
�                ��O�����bR�+���k-�                `&�ߜ��λ���q-&                ̪���_ׯ_�k1�              H��c��S/�Տbx�"�Z5v��4�T�S��_ f�����?��w/_�����CeY�����8�             ��j��h�����(�V�E�R�;�B �+�hY�1���G���y���Rr��o�\L(�*E%Z��G�����             ��(����z=  f�(s����v���nܸ�k��bB����q�'�S�P�R})��Vgk��             �t�V�����J%  f��w�v��w���o�}�,˿^6�y/��`��1:G�#�^o�z���?���F����l�              �EQ��  3��l�YF�_�7��d����������G���r?��A�0���0�U�V�'N܈1�             �0�8- ̺����t:?��������W��v���Y__����<l��ѥK�vc��b              `�E�z=  f����v����k����{�0T���a�k
�              ���V�{�� �A�V��w��^o!���믎{M�~�V�              �g� ��J%2k4뫫��4�u�b�s��/�W~�+             ��)�2  �E�w�F��W��P̜���+�^�/�ޗ�ZQ�             �F�~?  �E�w�Z�����O��A�=ס��}�s�x���J��F+����N�����#��ŧ�:��|L����ע�o             ��h��`0��3 0��nd�l6��g�9���P��G����g�����z��`��̙x�'���0MN-��g�>�l��             �ص��h�Z 0�F��N�---}cmm�/j����oeY���N̺�G����J,//              �cww7�V� ����ގ�Z��?^�z��/�������j5�|��8s�LE              ̞����&�` �,)�2677���E&������߭��=w�ڵ�5ס�^��~?fݱc�����/U��S�ܖ�             �h�(3
�4�8th�� 3`��t:�n���u2�k��������e^̱;�w���N̪j�+++q�ܹ��̂�?�w�L�s�Lw�            ��F��G�h�i�R�� �J�H���hii�G�z�����>��s��eǏ��/Ƒ#G             ��T�e���t �qi4�V���7o�|�����b#3c��j���Ĺs�               `��������F�O����$�A(f�?~<.^�G�	                ���j�~���^����^xᯋ�('y?B13�Z����s�Qr����?�3���&�$K���Tp��A*��b�Z�U+R����ފ�zzN�p@���{�-�
�E�mk�c-�F�X�AE
Jи���������|=��Ͳ	I�a^�9�3�������a~	�컻;���b�*                ��K͎���ʾ�ɾ��b��١���]}��Si��o~�bD��害�3zzz���#                ��r������XX?��o
�T���&j��ľ��|>�Ծk�---��v��o\~��b	�Y��}Ѣ��;����"                4�\.7��w���h B1�Pggg���DGGG                 +�P�2��磻�;���R�(                �A����p�\����]�v'&&���:::&�>����z�\.��e�}8�(��e���3zzzb�/                ����r�k�}qjj*�P(Ě5k�k���1<<�֭{����7B1�|>�����Օ�C                �-a���g]����, �\-�O� :;;���':::                �_�\�wM(�C*��GwwwtuuE.�                ��j��Z[�b��c�9&�?�����                �D(f�������]]]���                �N(f	��쌞�����                �g�YD�|>������+r�\                 �E(f�tvvFOOOttt                �|�b��|>�������\.                 ��P����===���                 %s���������r                p �b������鉎��                 8B1�I>��������\.                 K(�0��쌞�����                ��K(�*
�m۶8��3#��                �� s�tvvFOOOttt                ���С����=��y�G�P�W��Uq��gG.����ݻ��}��j               p@:S)Wb�<~Я?������}lܸ1�#�\.����߷K�P               p�:s������/�W�����                 ��P�ڲeK��/�rlܸ1                 ����<5�T�s��m.4��^����DSSS �cd�����U�=                DC�b�y���ΉO^��8�� ׽�{���               �H:�\Z����?�=���o�                �b�ُ�O8;n��8��                 XLB1s��rq��F��                 XlB1s��j�w�i��7�"~�����㘵�                �b�����h���o�u\}����all�                 G�P���ǲ`�����wo��                 8��b�De"               `ll,}�ј���|>�~��X�n]�r� �CM(               htt4n��������Zm�z=s�QGe�4�~���9 �`�               �Ƨ>����j�{���f.�bq& ���Q�t��� �"               ϡ\.?g$f!J�R6}}}��ZZZ���O
ɤ�L>� �P               <��o��yGb�K���ڵ+�g��r�nݺg�c��)���&               ��;v,�g��j188�ͣ�>:k=�b����蘉ɤ��`y�              �y�HL�R���T*e���7k-��g���I�z@�>�����'               �����Z��޽{��K�X|F8&Ee�1�t�����'               ���닕�T*e3�����2���c�������!               �Q�Tbbb"U�\�]�ve3�b���xLggglذ!�ʴ�� ��P               �G#Gb�T*e���7k��Iј4Oʴ��G.� ��C1m��hijY��5�5,�b��-˻885�Z-              X��^���/"���XL=$���1�ٰaC��,� �(:s�����N_��M�6����rE\��Xή��U145              ,}�\.8���jd���;k�X,΄cҤ�L
�ԏ�wQC�b               `>�$��T*e���7k�P(�ڵk�hL�ǤpL=(��ٙ��D�v               ��J������Z/�Y4f�ƍ��#2)*��� ˕P               �b�J�l���f��#2�����2��\. KUC�bF�Gb4?���,����]�}�Uk�              `yYY�����hooϢ1)��1��̆���% SC�b&�)��,�J���M�Z-              ���Z����@6����֋��L8&M
ɤ�L�XT8�:               ����T*e���7k�P(�ڵk�hL�ǤpL=(��ٙ�<_�&               x*�Jd���;k=Ed6n�8+"��[[[`!�b               `?��|��522��\�իW�d�s= ��S`&��@"               ���Ғ�b��j��0>>��Ν;g���^{{�L<&�d�q�6d�O�q�               �<���bxx8�HK�����lz{{�����b�ڵ3��\�ȤI�[`e�              �y{�B1,9�Z-�^��Y(��L���c2��Lggg�,/�Z               ��	'�?�p�rR�Tb`` ����g�555e�4)"S�ԏW�Z��#               �8�3���o�Z��LOOG6ώ�$�bq&���A�t���8�b               `���q�)���?�J�R6}}}��
��L@��y��u��pw              �s�袋�G�j���*�J�޽;����g�c:::f�2�8��pp�b               �9lܸ1�;Ｘ��;ؿR��M__߬����g�c��i֭[MMM�P               ,@OOO�ٳ'~��p�&&&��'������|���cRD��I�����b               `r�\��o�"w�uW �N�Z����l�R,g"2i���q�?a��              �J1��.�(^���׿��x��ǣV�px�J�l���f�
�,��1i��I��&              �:����+����������3344�M�Z �_�R�ݻwg�l)�v��g�d�q��X,,B1               p�����E/zќk)^122������٤�t-Eej�Z �O�ǆ���y���g�
���Lggglذa&&�nݺhjj
X*�b               �0H��H�u��Y��j5�W�xLz��cRH&f����T �O
:�{/Moo�3���|���g�p��ttt���G}t�Z�*�H�              �E�"�����J���E��I�t�w�ޘ����H1��Ed�b�8s�I!����r��CI(               ���H�y��9�SH��������,j��Ӥ�Z�����4}}}��R���=�ƤxL
�ԃ26l�����%               �T=$�q��غu��J��cR<&�dRT&M:Nׄd��V��=����w�z�o��4)$��2�s��P               �P�Ba&<1WH&�,���gb2�xL
ɤkCCCQ.�8�J�R6}}}���}�v������"PO�Ȭ[�.�����$               *��gA�4�7o�sO�Y�#2���ψʤ����D �N�R���~��g��{���=�ƤxL���cPG}t�Z�*X��b               ��*���/$���xL
�f��Z�t^��x����LD���w�z�W��4)$��2��\.,_B1               �A+
3Q��[��ZzHftt4����xL�ʤkCCC1==��W*����뛵��յk�f�j�ǤpL��ݸqc477K[C�bR%ijjj���?>��:��              X\O��%�����LL&M
ɤ�4{��r����{���w�z�X��WӤ�L
��w�rd5t(ft`4��b�R	X\�8W�lY3             ��|>�}�4�7o��^��btt4�]��I�������d �O�T�f���ߴiS�~��q�YgEKKK�8:               ,m�\n&$s�q�͹'�-�
�ԟ���8xO>�d6��ַ�~��/|ap�	�                �Z�X�fӦMs�W*�92������j�ott4>��ĥ�^�����%               �h�B!6lؐ���J�����fϞ=Q.��,���/})֬Y��zjp�4t(��o�ڦ��?T�_�� σ�c���X�&�=              ���X,f�y��9�GGG�x����̤����	�GL�H�����w�������y��hDu���T�����~"��z"               ��5k�ds�q�͹�B1�x�ӟ��)4+I�T��۷ǥ�^�               8Z[[�9�c�\�V�1<<�c����@����ώSPfzz:`9ٱcG\p����~B1                �Y>�����g3�Z��dR0&�c��)&S�J���� �w���8��s��O(               `��r�X�n]6���{J�R��B2)��ӌ��dG�#�<"s��                ,�b1��)��Y<�>CCC3��S`�V�J;w�̾W)v����9��!               ����Dggg6s�V�1<<�c����@������xjj*�@�@���x����
��%L(               ����X�~}6�S*���L}RT&Ed��޽{crr2��VJ(�V�5�&               @�X,f�y��9����bhh(���q�<�fh<�r9V�                �����l���T*122������٤�t-ej�Z N(               �C�P(����ٺu��j����31�z<&�dҵ���(���&               ����c�ڵ�l޼y�=�Ri&"3::���L
�LLL4"�                ��b���|!�z@&�c��L:O��k�Z�J#               ��Q�lܸ1�n�:k�R�d���IA����,��2����PLOO,7B1                ��B!֯_��\���lOSSS�)�JYXfll,���ٳ'��r�R#               @�H!���Y�&6l�g�qF���D{{{�j�,$SȤ�����#M(               ��W�¤I��ڢX,ƪU����#�?����r��磩�)�_.�cll,ɤI�ݻw���`���P                ,@��T*����Y�fM6�7o���B2���D�ٳ'{�,$�"4),355p��b                �I1�j��777Ǳ���ӥ`���x|��_���逅h�P�%�^[�[���Mg���=��x�֗�rv�c����d               И��b6�\.`�:s�Qg���N_��M�7��Ni?%~~���rv�On�               HC�b              �Hj�j���z͚��   �              8BN�{j?|�����=  ��C1ӵ阞�^��Z���J��ܷKQ-�]               ���������_�fM �k||<��~�.E��j                ���                 ,B1                ���b���,�P                ,��7
Ű`B1                �V�^�PB1                ���b�B	�                �"��r%                ��	�                 ,qB1                 K�P -ߔ��� N<��lֵ���ͫc�Q���?1��RLLM���P���c��c���S�O               �0B1 ,H[K[��/��oyy6��u�IG����z���x詇������|;{~���2]	               ���b د�Go��N�(.{�e���B��[�{�n^/{�˲y���Ȯ�x̿��_�~1��_��C;               ��YN�<-��į��W�P̑��1����lj�Zܷ�����-�y2               �Q	� Ŏ,����+�E,�\.�mٖ͇/�p������������(W�               �D(���t�I��s��<��Y,f�*4�/zm6�Fv�_��W��>{��               4���m˶���k�ug�.�M�XN�Y{L|�>��yo|��?7~��x���               ��L(�������揳@L.�;��"  ��IDATd����S��ȓ129��R���c�2���Y�&���Ѿ�=֮Z[:�dמ������s+�>�������ߟe�               V"��p�Q'���旽9�M��z�������ߏ��}/���w��]�����ӡ��De�ޫ��=�[w\����8��3�%Ǿ$��:Oˢ2�%��s���U��*�򮿌����               ��D(`+6����k_}m�Z�c屸����w�����1]�>$�kxb8�x0��|����\/4�ksW\t�Eq�)�y'�����������g�3>t����w}��}^               XlB1 +��_��cq�Q'.�5;�v��������}|��oFe�GR����y_67l�!V7���O�8^����/�u���=�Z}T�s��g�������w               �;���ӿ��xK�[�w�4��������{~|O�j�X*Ƨ���|>��|K\x����f�U�U���Ύ{�����/�7>���               ,gB1 +ж-۞s�};�9>���Xy,��r�_}��t;�]o�w���q�g��5��|��/               X�b He����s�����=�X�K�Y�&�E'_��?�O�0               `��h �j9���?���XI������柍��������Z��               +�P�
V����|�o�ۯ�'����������o��������\���               ����C1��R�O�/x����X\����߿��vI��?�����{��O|?�O>��ͥq�	�č��               �4t(�<Q�����/�J,����Y�}�$�P��n}]<��C���~������sqʆS               ���� �T�����j���               �;�                �%��C1C��X�[���c�������XΪ�               P���s��C1�T�����%�}`�|������7               �����j�P                ,�R��PB1 +X���Ľ?�7ƧT�               ��]�v,�P�
�+]������Ͻ=���;              ��cjj*`��b V���:)�����o}"~�~/Ƨ�               X^�b @.��w���������^w=zW                ˇP@���&��k{|�Ώ������L               ��	� 4�BS!���ڸ�E���>���o�}               ,mB1 ��M��=�{O|�Ώ���E�Z               `i�h`��B\{����b����}�             ��Da"FZF�5��|  �P�
vףw�U��*Z���{ɱ/�{~�����>��#Q��             �����@[<6~c� X���j������X���gS*�bzz:`��b V��v���������Wm}ռ{WV���\�;�uq�g����z(               ؿ\.�|>��������T�����x�'b�Ν�ux��b V�����q��� �>������<V7��w�Yǟ;޳#>���G��HT��              �HR����9Z[[�P(dA�J����1<<�E`���CCC122���j���I(�Lצ��{n���+n��x��wk�5�����������^?���               XIR&�`��ڢ��%�������TٱcGDLLL,6�������q����u_�
����	����?�����Ưߘg               ��R��E_ҬY�&�����O��سgO��倥N(��T�+q���~1n}ӭ��-/�w���_r}\��K��{{<��               X*��jg���b0�����ߟ�ki,wB1 ��]ƹ?7�9������bUaռ��;鼸���������D�j�               8�*�J���dїIA�4�L����g�P@�LW��7ė��Kq��ƶ-������7��x�������ձshg               <�R)��L����K
���4B0�_:���"��ܾ��V�}X���? ?x�q��ωkο&����XUX5���O�8x���_������              `R&�_�ԃ0�������5t(�_��;}��7m���zۉo��ν,����}UM�RS����o�/�Ǘ�+n�m[�ͻ]뺸�7��_��3���              h<O���b0i����r9�篡C1 �����9?'�9����k>-��y���E����q헯���9              ���R����P�??�xxx8j�Z��r�\�K��,�,��Jܰ�����_�[�tktm�wG�#nz�Mq��������9쟱\-�Xy,              ���B0###100���Y�%�ׯ�s!���իc���%L(���������mq���ć^�hɷ̻��]o��H��w>o�۷              �cccY�ehh(���g�/�<M�T
x>r�܊	���Y���5t(flb,ƛ��rr2��U.�c||���R4][��Y*ӕ�a�񕇾����x�^��ٻ��{���$!aH�L��xEq�Zg�׹(2*��[�Z��[](�hۧ�>�`U@E�Z��@���TGpDEP�B2<�y+<���$�|N���s����Y�`��w              ���KI���ˣ��t��E�i%��u��1���9����� @�ŬX�"V��b�)Y�f�PL#��������|I�9fL䥚�_�              ��*++cٲe�t��())I?�l׌d4��ݻ�E�b ��5�kb�������c�>��T               ���"JKKcɒ%�|��Q�ŋ��K����2�{�4� ��]��[O�U$            �dG�tDL�35 ��Z�re:�RRR�~��v�\VVДu��!z��4� �0�0�?���d             ��ާĻ_�o/x;2Mn*7�=���a�F�_� h����cɒ%�|��X�lY: ����~hΎ8����
�P tT������o            @ӰK�]⮳�Q�����12E���1q��8�ǁQ��,  SUWWGii���K�)))I��-UϞ=c�]w�P �jת]���_�y��W������q��������            `��s��o��v8(ν��(YYҨ��=N����� 4����t�e�����$��_/^��$��``݊���SN	�P 딜��}��ѳc�:Ϳ�����Ϗ�e            �,��yZ��u�8a`�6�?~��Vq���Ņ] �PV�^%%%��K2j�k��@Luuu �өS�8묳�u��A���[
rb�Q�㧇�4���78I����ńY            �\�:���/|>F=2*n|��=�!�b�n{ lN����	�|���+�|R�T���';�����P k��q�w�O��ţ�<��w^�[6/            �̗��7�xC|���9��I�HzK�gH�|��ѶU� ��*--]~��L2V�^��ӦM�h߾}l��V��v�E�^����(h<B1 �O�\q�q��/�Tvj��KV��������            ��9y��c�m��3�<#^��;~AnA��_Ņ] P����X�d�ڑ�_�8L2.\(�]�vѩS�t���8��������E(��ۿ��q�w�.�w���'�{"ν�����             ����o3Ο������]TWWo�u{w��O�]�������� �Seee,[�,�/_�~�	�,^�8�]RRUUUlY999�LM��1�Ν;���t���B�r㗇�2.;�He�68��e�ӿ�4���6�	            `˙����wX��ԫ�9y������О�ƈI#b�śt̑�G��+�-X＊�����+��i� MSEEE�����/I�%��$�k�K^�&FAA���K2�L������
���hϮ{Ƹ3���������s��9�Ή�K�            �4�5���{C߸��[�}�Z��w?1^��8��3�ُ����ڵj8�q�>gnp�g%�Š;��= d����X�|y:�R�I0�H�K�	�@�H�RQXX��$�$�R��رc���-�P@���?��Ob�1cҥ�Y�fE�yrL\���QU]            @�R��4�=8���d�|���&�M�s�+�.�:���f�51fʘ:_S��6�Ƥ!��gǞ������{�Ǣ��ƕ�`j�/5A���If�ʕ4����t��s����$�Daj�����b Z�=��#Ɲ9.}ҥ.����8���c��9            4m�g���?}9&�����u^r���G���v8(��_:�ֹ���ta�=nl��i���WTU�;@�ƫ���+V|+��t����d,\�0V�^@�*((H�_j�7c0ɀ�h�3?��O�ʣ���ɖD�����+����w�            ��w���n���q�J^�����.y-�LSfO������������:}���d�'q�g��< lk#0˗/�e˖�C0�/N�WRRUU����J����0}I0I�&ӱc�����B1 �خ]v��g���������D�������            @��h���^3?�7�rs�mնֹ]�u���},��zu\5�����L�߯{��g�=��V;l�xy�/qΤsbI�� ���I�/I&y]�^򺺺:��WPP�6���$�Daj�������f�?�G�"1++V�O\����'k            ��k¬	��ܗbҐI�W��j���N��F���rp�8$N�����#7�����k�F=2*n|�� ��������˗ǲe����u2j�0@�Ib0�:u�Ν;��/5Q�$����X�b Z�7�x#�M��{-            ��㽯ދn: n<��8o���;�О�Ƈ��a��6��_�'L_��RՄ`jF�I�/���E�bժU4����h׮����7c0I&����3Z�Օ���WǵӮ����hJ�v�]����L            `㕯)�������}<���?GqAq�s���0kB�����|�� h	�����s��MG`JJJbٲeQYY@�j۶��LM&�NF�6m�"�����oư����_��"9�t��Gǐ>C���'Ǥ�&	�            �f��?L_ot��{b������Ip�?'�g��?@KPQQӧO�_|1�4�T*�����K��7�sss������"~3�71��ѱ�bU4�u�-������v            `��x�������]�x��#++�N�{{��1p����Z���Ҙ8qb̛7/�-+???ڷo��$�5#y]TTT��@s!�B$'[ξ��x�ӗ#����A:3�ǀ             Fr���oN�a}�EQ~��/Z�(���1�t~ �"1��|+S\\��0��	� 4sU�Uq닷�œ/�kVD���ʎ�z��Ü���:�u             '���ˏ�<.;��v]th�!^���8��3㹏�����z���Y}�f �f$����kh��|5'�����'Xzv�g�=;��7,�-�6            ��׹m�sНqd�#������c��3⚩�Ę)c�7�h�>����?��w|+�R\\�6
�lgee��Zv(����UW�}z=�[F�;�[����!2Q~N~���	1���8����a            ���OGb�n��F������v��J@s3e�׹�b%���/��f&���ly-:S��$�.�[��I�
h\K�,��s����H-8��g�>�8̙���Z�            ��$q����*~~��7x3�E+Ōf�)�OY�#v:"f���t�x�����X�`A|��g�YNNN�k�.~���Ԅ`:w��4.�B ��n��bH�!1���ع�Λ�^�겘����[            �8�mO��v8h�s_��R�q������
�|��ѶU���=�G���W�US��ʪ� h��|�̀�m۶k�/I&5��}@f�`��K���;�>�s�'En*w��KN�0��?s|L|ub��*            `����q�wD���;���:nz�����KcM��{fM����L����]�gS٩}��8�_��w�y��@S�駟4�T*
׆`���׆`:t��Z�
���`�٭�n1�������ܶ�&������q�q3�����            l��윸����#/�����]X�0�N����w���jv�b��c�.\�:��<4^��z��x�������/2E~~���KM&yNFQQQdee�<��P�/D�׏�ZQ�"�~� ���QRQM٪��IQ~Q�{`:3�ǀM^���Ǥ�'ş_�s�Y8'            �M׽�{L<1�q����`F�u�Y�y���YY�2.��E���Oş�9���un�����s����).}��XS�& �����X��y]J�+((X�IFM�f[Z���]9�^�Tu	�q}Z�i|Z�iи�ZprBhH�!1���h��z�֛�l^����q���ų?���            l'�~b�6�ت�V띗\�Sߘ�_��K���+���P��b��0�w�g�yF|��� h*V�\�����|+S���~��O �l�;�������튷�,k���Mq�CGeUe             �O��Vq���ŏ�8jY���C&�'�{����d�'q��98.;Ⲹ����7��M�����K^�s�=7}�i�� 	i��(((�V����xm&����� �L(����ɏv?!F���<|���s~�|�            �.��Eq�Anp޴9�⬻ϊ�6�XUqœW�+����=�j�U�s����!��O���+W 4Uߌ�t��)=��$��� ��P �t`�c�~��{� 
�7i��K�F�T��ҮK             #'{���&7��rʕq��k���j���}~�O�=���c@��Z_|�ű��c��> [NNN�k�nm�����[a���� h(B1 ��u��c��cD��g�=7i��5���fM�G�}4�8�	�            �_.�2�=8�̞���Nn<}�͇�eG\�yydge�:w�n{ 4������d$1�$
S��� 2�P@��Nš;#�����8)rS_-L����|��9>&�:1JW�            �Y�͙����/��ŎQQUW<yE<���q�;�7��ƒJ����0~I0I��&
ӡC�hժU 4B1 -Ԯ]v�a}�����G綝7i���z/�y��?k||���             2Oo�f�51fʘ�M�B���7{ńA�^G l)999Ѯ]��1�N�:�G򺨨(������hA��b��chߡ1�ǀMZki��x��c���1��iQ]]            @f���8��3㙏�i�c���8�O����Y\��D*; �1


�ᗚQ\\����lgee@s&��egeǁ=�!}���>��un�^���2�0=&̚��~�X�"            ��6u��|��XP��ѾCr�����s_��Ϻ;�v��j��[GѪ�z}�C���R�(,,L�_� L���t��1����%�h�����{���^�}��y��Wc��q1�Չ�z/            ���T��+��2�LU�U�	f|0#���^1�qq��FK�ey�辬~�|�)�梠�`m�%I&���lgee �&Ќ}�_��ё�/�}��q_�{y\���+            4-7<}C:�i�-��o;>~v�����" 2]vvvPwI襨�(~�	�Ԍ�u~~~ �q�b XkUŪ�2{J��5>���_3�$            P7�|}Puuu��>6��?- 2]AAA:~���������ڵ[)..^��ԩS��� ��P 1�Y1aք�땻�5^            ��0�ә�鲳��u��QVV-I�6m����7��H O(��Jj�����ƭ/��/|?              X��ݻ�;��I*�����h߾�� L���:D�V���"�B�r���
�����c��Ӣ��:              ���={6�PL{���$1�dԼ.**���� ���h���cH�!���W��=���g��}              �?�{���S�Fyyyd������d��$�YYY@� @�Νv��G��ˏ�<����?s|L|ub��*             ��,///���4����t�%	�$��LM&�@��O| �%;+;��7�tc<���1aքx��Ǣ��"              Z�$3{��;w�f_���`m�& S3
#+++ �E�b���{�u��u��o�}h\{����M�C��UU��X������^��}���/������uzz�[6/��������y�             @K��Zw�uW|����lQQ����?�`�P lH�����ؽh�:�ߺSݣ2���O�}��'DS��',S��$����c�.�ư��b�~ãs���^�[a������o�������o�/�              -A~~~�}����K/ŋ/�K�.]�/''�[�d��uqqq�R� �MѢC1 -�;މQ���_>��8t�Ccd��q�'En*��k��e���q��k�������t�f�cu��              hΒ���˖-����t$�]�v [�P@SYUS�LM���m�#���=��Y�R٩8b�#�ci�Ҹ��{c¬	����Fuuu             �ka��١gtl�1rR9��bu|��˘���X�bQ�|�����K��;ﯪXC&	�����0 ��� �`�K�ǍOߘ}��#���3�93ڵ�����8��d���1�I1n��h�G            l9YYYq莇Ɛ>C��^G�6E��:w��91e���s֝��'�7�wܮx�8}�ӿ�~�겈�  �A��,\�0�YX���[��q����u��f�����D�>�?���q�C��i{�#�������I��ڥ�.1���q���������Y� �             ��눝���Ǐ�}�ٷN�w�Sz���1�әq�ԫ⡷
   ��PL�� �-)���9.=�J�}ſ���c��^+;+;����             6��T^���w��m�͢}����O�)���^s�	   s��P ����Oc���q�S��a=��}�Ʃ{��s[            �8�䵉�G<��<t��wd�#㕋_��rA��9>  ��$�UUW��9S����Ǡ}ň~#b�n{o���:U1�Չ�0            P��Tn<x���-S�m��1�qqx�����嫖  �Y�b ��E+�M�ܔ�o�{�3$F�7":��Q���a�{�ظ��k��O���^�/�~���j�W            |ۯ��U��-��оC������;N���  @��`��5���Ȩ����ɥ$sr�#'���dgeǀ��7'�&�0=&̚��@��.            h��������qzu�3Ο��阘�٬   2�P �lUŪx��ӣ[a�t0���ύ�{n�z��T���q˩��#o?���<��cQQU            ��$7j���"++k�󪪫��O����z(}���DUUUl]�u�;qܮ�������:�t�i�>-������G�  ���b ج�-�c��M�>�����GƠ}E�Vm7j�ֹ����NO�E+�o<���<��Q]]            ���穱��{�w�s?�9�?��O_����#}�Ѹz�ձ[��b�a�b���)�/���{<N��xr��  4.� ��Y�͊��ø��Kc��c�~���n�zZwH�g�q�s����            �����w��_�s�Z�ʪ������c�ġq�K��N�C��ԫֹm���C#�3�<#���_  h<B1 lq��J��oM��;�g�sf�7<�w��5�            Z���o�8����f����;/�����S<{�f�}�����?����u�k��*�z_�4<�ug   �C(���W��O^c����z#����81�Ry            |ױ�[k����^P�HL��+���"^���wƸh۪�:��d����kx�  4<� EUuUL�35=�����:=~t��b�n{            ��%7l�ͨGGE��M>ƃ�x0�_�~L>9zl�c�s����SnI�4��gn
  �a	� �薔/�?�����}��cH�!q���F��            Z��n���W������f;�_��~�/�r�_b@�뜓��7�xc�r�3~  @�� ��5���Ȩ�������-����˿F*;            ��$A���/��7���QU]�Y������?��O��w:|�s�X�oN�M���W�U   C(����bU���}�mѶq־g���#k=�            �Q��������}3>��E�Y��,���������]��u޵�^��Ō�2&  �-O(���Y�g1v�ظ�����Ɛ>C            Z�$S��_��b�]Y�2N���8xb����Z�]y���&�M����  �e	� �dTUW�3=��U�           �9).(�uߢ�E[�ث+W�&� nx�zo���C��T\��  l9B1 4II4            ��6ymjݷ�b�?~eUe�4<�|�~g�:�'��I�d���]���  l~B1 d���!�j��w�_�bq|���            ��l٪e���ئc�]:w��$3��Q��4~|Џk�w��.��܂��?r�h  ��b �hWsU���Y�y��W��w            hΖ�XR�Nm;5H(&Q]]M�(*�*��/�u���##������� ��L(              C-)�=ӹm�hHI,撇.�U�b�a�j�wN�s"';'ι�����  `��             �P�W,N��Zo��}������}����/�E��)�+����9����Tn�8,*�*  �tB1              ��y�ǡ=����pP\7��hc���kV���__�A���T^�kP   �N(              ��6�ZC1�Y�QU]���O�:}�_�����Z���<-
r���	  `��              d�$�.��G﮽��y�Gc���FEeE�p���b�����w�}  �4B1              lڜiQ]]�����6j(&�g~�k�����>����9�ka�   6M�Ŭ\�2��YZ��:t�q����ҥu��f��             ���K>�7�����ξ�}���_�U�ј��⟢���N�C��  `Ӵ�P̪����G]���и�PLII��I(            ����{|���m����z���X4�[_�5V�^����T   �W��              4I槇�t����wNF�bw�zw:s����bj�E�/�,��^��ئc  �P             @���������ئh���;i��b�λĻ_��`¬	��bU�u�]���R��e�/ӣ>�
�� �yj���^S�&*�+�<�*�*��U�U�Yu��f��             �QU]_��r�w���Sq����Yw������M�Ϻ;rS�  l����zb�����8���x�^����ʿ          MWY���   �玙w�3�����z���΂w"S����Q��<�@��i  ��iѡ             ����o�_�{v��;�R٩����c�]�"�<��#q�'ǃg?�9�  l<�             �&�����T�:�U��D���Xv�aѻk��쫨�  �n�b              ����e�<���?y>=  ��'                ��b                 2�P                @��                �pB1                 N(                 �	�                 d8�                �'                ��b                 2�P@3�K�]bۢm�)�Z�5               ���h�~|Џ���               �i�                �pB1                 N(                 õ�P̨]F�n���y�6]�	�q�nP��h�.x��(]S                uբC1�S��MN�:��O�и�Ry���f��                �ѢC1                 M�P@36��c㶗n��h��               -E�ŬX�"����<���4�5k���w������Xs��M               �ikѡ���(�.����+Wи�`SYY����!C1               @�ТC1                 M�P                @��                �pB1                 N(                 �	�                 d8�                �'@Z��n���ѻk��ѾG�o�>��I�+]U��ǋ?���/~�b,Z�(               ��!Ђ%!�����}�F�m�FVVV�>WYUO�t���1�Չ��ru                [�P@�a��wn\{ܵѡu�z>���Cv<$=�3&.y�x��               �2�b Z�����0hB���	�e���������m/�<xA��X               ��%Ђ$��'G>�����k��7"�-�6N��D�               �̄b Z�Tv*&��E"15��uT�6�tנ             ���m;ǀb����V�������ͧK�K�E�+���/|?  ��K(����ῌ�w>z���}Ό'�{"��            @�P\P��;'F��u�m���.�w�rW���ߧ� �M'���a����h��]��1��ɱ�|i             '?'?v�ctl�1r�sc٪e��|>Z�Q��\S������.�����h�צΟ�^�=~q�/⒃/��~�����/��5�  l<�� ��$'x6��E���=����ļ�y�hŢHe��C��}���О���;[��z��tj�)�?���_��W             [�6E�Ĉ~#��v���g�}�����+���_��oN�q3�����\7����a��!;��߭UN������rl���k�Z�n�ݢ�����L��  �b ���Zo����9I���.�{^�'���j��� J�3��?/F5:}��6� �N�U�            l~�q�1W���t�e}������s̘�n�uq��k��u�ҮKL9%zw�Y��]v����8��c�W��%�T�)�/�^��V  � 4s��>u�'yf|0#Nwj,Z��N�%'~nz�x�G���n]v[�n��ҥ�is�            �y�تG�m��b��w��g�Ryq���1;G���X�b��'�#=v�c�-S#��<~�������9&  �aB1 ��q�W�7���zl�X����~���8���ū�]��sNr�H(            6�m����/x:��)�n�7��d����b����>���g�}bK�a����!Nz  ���{������˵�Isk�
��B��r�# �P��eDgG8�Ł3�=��3�KE��((

3xA��P�S(��M���ٹ�$��~Wz�씴�ms�|��+����<OX������2B1 cXaAa;�؜��ޞ8��s�*3`m����_�]��S��9?�]�            �?�E�q�'���H̀Cv?$�;庸��Wg_��e^|�}_����ύS�95~���  �P���=�6U�sv۳��������{�w���'�șG���Q\X��L             ��ړ���]���]�~�۱�uu����{�X�9�-y(�\�d�k_�]�QV\��'ǾS���>1�������Ӿ"  [H(`K~�2��?����'�V�P̄�	1kҬxm�k            l�ݪw�+��2��-)*�O�����?��:?�9+�W���>n^x�;�b���8<���/��sN�$vs̬c�7	  `x�b ư�����ؽ1�Z�T����k9�V9M(            ���#.�TIj��m[�,�'}��X׾.:3�1�bJ̝67Θ{F6㰜_wּ�bEӊl4�o=���8��ψ�tӰ��'W<�������+�}%


r�w��  ��ê˪s�/\�0zz{�v�7[ތ����^5}��            0|Il�C.r�������7������y���>N�sr�t�M���z���]���?�k^Y�J�������zK}��_͆g�?�����������  �;��jR59�W�����V�����{             �神G��HB+���'㖅���u�{��8���C�=s��ٴ_TX��9e�u?q�'�*3 �ל���1���fS&N�y�̋V�  �;ס����x���a�_^^�����o�9��vD��q��.�ι��є�{5v4n��             �IsNr��'~8�H̀�F�g�'���l f(��v<������L|����mݖs~�G
�  �0��PL_���c����ع�簷w��툴C1�'��O���~��������T             �f�n�s�o�����-��ӫ��[��5.9��!���?�|��Ż���zR��A��v�/  ��ס             ���������_g#,[�gO�l����_�?�+����H�5�A��&�  ���              �`�*c��=r�������>�����{cT�V��l^6n�|yf�39C15��   �g\�b��<+
V����� v�e�ˢ��7F����             ��Tm�=�����n�/��.��f6h�ʺW"���^uYu   �3�C1��n���T�V�s-�[K2K            `��,�̹�����/ަk���圡��ts��P׫N	�  �p��P             �HW5�*�~{W{���lӵ�;s\Z�Z#�Z:[r�W�	�  �p	�              �`'L̹��ն��n��}�Ξ�ȧtO:�~q��� �p��3             �VXP�s�+ӵ�����}���~   #�P                �'03�����z����s����ǔ�S"ߞ]�l���m               �P�8t،òkG8a��+�n}�V�               ��                �N(                `��                �b                 F8�                �N(`��tS�E�7               �B1 c����.               `t�             �f�̈%W/٦kԖ��ܿ�K��}O�|)-.  `��              �B%E%1{���r���  F�               �B����aÆ����O�4)R�T ��"               ����O>�d<��c�����YYYY6S[[�i�������� ��5�C1Vu�u�>����`�ګb��c�1�=��H���              �KWWW���?��˗�wvvF}}}v�����������۠LIII ���P̹������]v�%���S�g�}f�fi�K���              �G���2�Nz{{���!�r�����I^WTT ��P               ��?˖-�n�okkˮ+V����f�1ɪ��y�q�
��O(             `[ټ2~��c,��t�h��d�G�i����5k�d��J"1���Q[[�)��.++ ��             �l��E�;> �</��b����������)��.]:h^QQ�)�րL򹲲2 =�u(���!{�}~�@`�������?�#Q�/              ����z�V7n̮7�|sЬ��8������l��L�2%JJJ��c\�b�2Z�����?��+y��ed)+.�y�̋�����Q^R}�}�a�Xָ,^]�jt�t             �H�+�2d2�hjjʮ�K��mVPP��՛�1IH��eee��5�C1 l�T��zI�2�8jϣ"U������xj�Sq�swĭ�����             ������M477g�o�1h�J�6�c�USS�)&�'� �K(���:�;�����ˣ��tX_��w��Gg�WN�J|���ė��r�u���y             F��������.�NgW}}��Yqq���1�z�q2`���'�8�[�n1�xB�YSGS4���z�#�8"n����Y;s��Q^RWU��������O�x2              v4��-��dbÆٕK*���I�[�2�qAAA 0�P�W\X/\�BԦjsΏ���xh�Cy��I{�����̆^�a֤Y����1ι������            �h��zU���l���U��X�N�����~Ь��8*++�ј�S�F]]ݦ�Luuu�x%0ƽw�{��ļ���xx��y��>S��_]�EbT�V�]�+N��	���'            `�ڐڐ][�+� �E&������Z�t��fEEEQUU���$񘚚��q�&O�&L��L(`�;}��C�n|�������}jR5q��ݓ��=�JRq�E�Ł���h�l              Ɨ���!#2�T*�)��$$�e�

`4��Θ{F��������[�v��O�>���;����3��o�����              ��J���U__?hV\\����hL�I�1A��S�f� #�S�a�V��M�/���go�tO:/�I1���a�ۜn�^{ �[�\4ll����V9-��6?N���(-*���_z��G���5              `82�L455e�ҥK�S�TL�2%�ykD&�ʔ���H 0���C��|�μ��+�}%J�J6{N�����M��]����Ԧj��]WՐ�K�2�9���3            �X��{��-��q1m⴨��������?��7[ތ��ǂeb��E �E:��+Vd��J"2�d%!�$ 3p\PP ;�P�v����߰qC�i��r�i���C|h��,oZ���i��ڗ7{^S�)���ڸ������C6���/�+�2ں�            ����uL|������yL�0qX_�F��~�]��h�h ���L����͊�����*�I�1I8f (SWW����/B1 cؑ{�s��E�D�/��{\x���
�P�=�8��������Z�ra|�G��?s�JR����N�{z����            l?�U�7�sS��ߙ[���&͊�O�>�x�q����1��� ƒ���hjjʮ�K���R�M�d%!�$(3eʔ����-!0��{��s�?���y�����f���{m����-��c���xC�A�$?X�           `<9|����圭jY�y�7y��������cw�����t�������k���iq�-�EKgK �&���[+�NgW}}���@D&	�|�TUUEAAA ��P�U���_�'�-|sa^��=�]r��p�{������C߈K��4v��}�콳�            0�|崯�I{��s��w�c^�u��c��KⲼ]��9'ǃ�=��t�X0����fc1}}}����LQQQ6�րLr������K`���fM��s���-�[��{$?�ٜ�.�ntf:���=q�S7�5']3h6�vf�R�K�i[            0�U�U�~��������^�{��䎼Fb��m~��_�i�~Z����hPPP�T*6n������FSSSv-]�t�| "3�8NVEEE c�P�5{�����?}��)Vn.����x��|�۞�-g(&1w�\�            ƅ���E�9gI$&���Cr����Ɣ�Sb{I�Y�x���� �Ŵi�r�:`gimmͮ�˗�Gee妈LMMML�:5�L����QXX��$0F�Z�k��5���l.��ʧbY�m�ǋk^�խ�cת��<s�̉_0            `�;}��s�'���;�~'o�����]����S��_<�Xټ2 F�3f�0jd2�hjjʮ��s[TT���$�$$3�^���0r	� �Q�*s�7t4���uu�w��C�\��������:qj            �xp��cr�/|sa��ᵼܣ&U����9�s_�x�����`ق�/���tf����>g�vT�U��e�e�{}�W���`�����~8`���������%�J�- SSS�)"���� �Q�9����y��!����#K�|yi�Kq�>�گ�P            0�M*�{M�+�����}�p�br��͞��}]��/�.~��׃fk����_��x�?b��)q�Y7�G�t�k]t�Eq�o���/�؞�M�ӧO������,�NgW�?륥��2�e���ؾ�b ƨ�	�C1I�7�q�f�O,"�%��Q.�*            ƺ��8<


rΒ(K>����f�y���8�{�Œ�%�x�����[/�W׿_:�K9�I���/�o?�� N:餸�[ƫ���X�vmv�J��ј)S�d�[�2eeel;��1���?���҉y�����Yָ,��֮֜�UeU            c�{�s��/�����r���u\̬�9�<ӗ��z��"1ou���^w�͇��P0j̞=;�͛/��R ����쪯�4+//[8�Ǖ��CF���Z:[r�WN�����qؐ��W=���՞s?_�,            0�͝:7��c���=.>������c��[u�+�2>8�1�|Ҡ�{g�7�>���� �:�hhh�5k�0|ٵjժA��������������������� �B1 cTK:w(fת]���3jf�nջ9f�3�OE�E9��2]            c��ɳs�/\�0o�8y��CΒ��|���n��:�k~-�v��͊���=�^{  F�$Xq�����+V�`����FSSSv-]��m��������d�1����T*0�� �Q͝�9����m���3����/o�%򩢴"�~kWk            �X7kҬ���zϻ&�k��X��E�ě-on�=n}�����_��A�Cv?D(U***�c�X,X� {����`��������Z�l٠yYY٠���quuu64c�P���}}����3�6UM馭�����r����-{,�i�ĩ9�[;�b            ۪ʪ���.���5/����>f��_<�m�Ǫ�U����|o�>S�	�Ѧ��(�=��8�#b�ҥ�|��hjj�����J��lI����>��V����l
��mP��Xr��g\����ꎍ�.%7�������n�s;������I���yg�-o��k`���=���h�l�|�Q3#�P            c����9�7vo�tO~"��:�����ro^�����s�bfO� �Մ	b�ܹ��V�L&��ڲ����hooϮ�8�knn���� �����hhhȮ\R�ԦpL����@L&9Nޗ#͸Ť�ұ�mðϟ<yr ;W����܎H};�6��Es�9jR5�fy�G�:3����=��?���ȷ���˚�            �e�9�;�v�#�8b��S+���������/�ܯM��XS\\�)>1{�� V�hmm;w6�<�IB2I`&9���	`�I���U__?h�<Õ���g8��$��x�ԩ��Daaa��0�C1 cY__<��#q�~g����ǡ3��+n�u/;���x�ȧ�8p�s��[            0��iJ7����N�w��#K�|Y�>����˪`�)**��J�H2�J�2I@f�u����`��d2����K��m�Db���Ed^���l/B1 c��^�]�PL_��Yߊ�w\d�2þތ�q��9O*���z_�Ӽ]���	sΆ��            �C�b
����w�E�ECΟ\�d�Ks�9�~eYe 0X*�ʮ�ӧ�'!���L�inn�F-���J^����_}}}CFd�s;�IV�I2���{�P�v��wƷ��v����{?8��_}jX�O�27�sS���yί��Ut�vG>���	9�:b��            cYg�3�~���U����Ο^�t�K[W[���	U���L�2%fϞ=h��d���$f��d��L���dOH��$┬���A���⨬��Fc�xL��$�rIII���P�/{~%�HN�=5.����<��h<��_�vg���ǎ��}]���q�A����OƤ�Iqٝ�Ś�5C^���:���3枱�����E������f�3            c]KgK��ʲ��b�qؐ�Ǝ�X޴<�;�{�J�J��,;ӗ	 �'	R(r�dz{{���cSLf ��Nֆ���;��IN��ҥK͓���s���S�F]]]6*SVV0�C1�}��|W�/�����]�]��}���Ǉ���(,(�9?{��ㄽN�;_�3�~��XҰ$ֶ������=iv�����#>uu��ςe��7���>�rZ�4礜���<            0�5��s�O.���%�I�e[�g�{����ͿD>���~ssg�S$`'(**�����>}z�s�����E{{�ۢ2�����9����,y�U__?h������l@fภ� ��u(`<xf�3q���}b�s�(L2��9����]�v���%�\�b            �
�$��e����?m��w��%f��r��P��҉9��:���)	S$k��L&���I�1�����{����� ���"2I����*�I�1I8f (SWW����� 0\yϕq��'Ō�����y�7�В��~݋�8�~�'O�|2            `��ؽ1��MQ��4;|�÷)sҜ�6;xi~����ܑ�֮� `t*..���={���[C2�����ښ��$Q�d���%����6����g*YK�.4O�O�j���L�x��!04v4�G~������GyIy^���eU|��OF���1��9g�-{,�2]            �������=��ށ��7��V_����r���Ă7D>�Q�G����O �Mo�%�No
\$+	�$q�dmذ!����6�s�����A��9����>�S�N����M����(,,F��q����y��w\rG�JRy�f�'�Ьk_�v�qW9��Ż            Ƌ�V>�3s،�bߩ��+�^��kVN����=m��3������ȧ�w�?��k^ ƯT*�]ӧO�9ooo��cZZZ6����^ggg [/��l
5-]��m��������Fc��sϘ;wnL�<9�y�b Ƒ߾��8���㗗�2���#�����q֏����)��L���ќ�������#            `�x�����|a�~AAA�p�q�����k~���gc1C���{#��~P���� e�ĉٵ���'���x�[?������`<��퍆���z������:(N>��(//v<��q��+�~����i_�O��(-*ݢ�OB-�={[\��bU˪��=^s�5QTX�s���ǣ��>            `�����cc�ƨ(�4;k�Yq�����1��U�U�U�_��s~���#����g��䜽�� ��UVV�]ӦM�9�d2o�$!��5�Ib�;���g�y&�-[\pAL�2%ر�b ơ�Ζ����!����㓇2�9�������,iX��z_|g�w�5/m��mﺽゃ/r~��w            �'I$����0����4��M��k�㵊��sn�ݫw�+�=�2��Q���9�`{*..�ɓ'g�P��t455mZ���ـLr���]]]�?ɳq�-�ĥ�^UUU��#0��l^�����\>9��u��5iV���g�b���x��X޴|�|OI���o9�����            �77>r㐡��������o��������͙2'�}����}N��~��'�og�;+�~[W[,Z�( `gJ�R�5}����7Fsss���FKKK�8	e$��JB30�$1��n�-�)((v� �:��%g�δ�}]v            ��S+��߼��8c�9��/���+���q߫��3�����k���*��1����gŅ�k�-oƏ����~���/:����o,�L_& `$���Ȯ�v�-�<��d�I<���1��۳+9N���L�XS__.��;,�1�b              F�+��8q����l�s&O������������ȧ$R��=s�^�s�5 �Cqqq���f��ٳ�{{{���%��h��~nmm͞��C=|p۟P             �(�x���+�;��v��S+��?��_��C/r���
 뒀ƤI��k(�t:�������=���6�nll������ _6n��/����/���b              F��.�n����|&��m�h������ۓ��V�UŹ��s֜n��i ��T*�]ӧO�9OB2�����Ғ�sGGG�βh�"��D(             `��]����~|�=����ںڲ��e��"�>���GuYu��=���{� ƪ��̮��s��d���-������=Z[[������^�����V�X�B1              �Ho_o\v�e�\�s�3��[}�$s��=3^\�b�[UYU�ӱ�4�����  ?������6�r���͆d�xL��Ǽu%��I����3���b����/�L(             `���ߏ߽����/����ams�9���oƷ�V�v�n�������T>)笭�-��� �EEEQSS�]CI��ـL���۳a��׍���e�ƍB1;�P             �(��iy|��O�U��*>��ǉ{���~H̨������խ��%�����^��l,f{I����}"��M9�w�xwtf�� F�T*�]ӧO�9OB2---���ܜ]���$��5�BB�1�	�              �r����w|7�e�eQUV�������;��I��c�� `����.9�L&��ڢ��)��ۣ��5�ill��%1���� �޸�|�]��9Us�}������u�ng�������?bcF            �~:3����  ;Jqqq���f�P��t63����@\fÆ������u(fZٴ�=���ϯ+�`�)�٢�v$*.���              ƩT*�]ӧO�9�$����hnn��I�2ɂ�L� `��������ڻ�c]��               Ɔ���P2�L6��c�!���L��������b ư�O�>.?���n}�ָ��              0>Gmmmv͞={м��7Z[[���=�y �De��Lr���0Z��PLWOWtww���,�\�s�%��H���               �WQQѦ��P��t�����Օ=NV�I�2�}��u(�uck$�USS�Ε�G5)��fB1               ;G*��+V�m���2�M����QRR���===و̆�!�丽�=;��a\�b                ߒ LKKKv��^{�uuu1{��(**ʮ���������l4&��$_�~��lL���YH��F(                ���_2�Lv(((�����>}z��~ِLqqq���Fwww���l@�7ވU�Ve�4�-�b                `�mL&	ɔ���̙3�+���7n̮������_|1��0B1              ����:c�����:�  F�	&dפI�6�-Z�(z{{�C(`�џ-y(ƢM+            ƃ��c�n�c$��tEGOG�������cm���������0�����k  @(`{z���            �^��84����2}�Xټ2��.��6x�xb��}   ��b              �*Ņ�1kҬ�:{���S���ts���m�����˛	   ?�b              ț�TM|�=�ͮ߾�۸�w�ĳ��  �m�b              �.N�{z���)q�o���_���'  ��#             �vS\Xמtm��Qq���Ds�9  �-'             �vw�^'ă�=�}�h�l	  "������7`8�b              �!�~P�������L  �wS�N��+W�P             ��p��8�'�HP[^�Q^Ruu1w�ܘ7m^�3u�(-*�5�������k�?\  ��ĉ�K(             `k�h��_�?F����8�]��G�4>����&U���9隸�����/ �xV^^0\B1              l��ޞ�������;/�ˏ�<�t򗢪�*��Ņ���ӿg���  �
�K(             ����tƿ>��q�w�ݟ�;�����}p�Ɯ)s����  �΄b �ٓgg(�G��{��1�jzL(�5��(,(����H>�:��+��ZWŪ�U��iE<���x��             Ƈ��D��t|,�����}�

�3G~&���   ޙP CJj����8e�)q،òA�mєn��V>�_������+^��z             cWcGc�s�9����Ң�A�s<G(  �I(���8ab\t�Eq�Q�����kצj�љd��3�O<W�\|��ŭO��7            0�,Z�(���w������ڙ1o�y�Қ�  �<� �&O�<������T��继�;~p��3n��>�ո����;            ���[�|+�p����p�쨙G	�  �0� ��u|��y�����r��Tm|�_�O���W��CK
            `�Xټ2��.��6�,�  0�P�8VPP����g~#�w����+���������r߿D__             c�_�c�(�>S�	  ����*  ;EQaQ���?����I���K�|)�Ý�~qd�2            �~���h\�+��^�{   �L(`*((���q�!�Hu�A�G\�󋢯�/            ��mu����*�  �΄b ơkN�f�"1K��ӫ��V�˚�Ś�5���m]m���d�)),��&Ɣ�Sb��i1kҬ�������o����h��������s             �[�^�\�K�  xg�:���6d}2��'�s�������nG���{�S�ןz���l�c�ӿ�4~����F��t�$s�>��E�\G�y���暓��'V<�}��            �^s�bJ�J���x�/�  rס��޾�����������-y����܎H;1��ux����p����������w}��楼�?	�|���g�~���>���w����'�����ܯύ���             F�$3����   6o\�b ƛ�O�:f����9K���~�X�l�v�^�]�����柾7���g�>C��{��q͉��տ�:            ��ir���]�.�  ��q���.���/n��{_�7���y���;ʟW�9�׃��o���?{�������1ִ�	            `�����s��{ǽ�	  F�q�y��h.h��e�e�\k���b��1������^~��Q^R>�����#�ӻ㿿���8��s���q\|��9ϙP<!��迏k�6            ��g��Y9��[�  xg�:�x��[t~o�7���ޗ�-SZT�;�sC�����q��H̀޾���/?�{�%g]|�73{�lvs�$�%\BJ�R.���@Т�
U+ڣ�ZK{<mEO߾�}{U(��K�*o+r{=h[���P�\� �����wf�}�ξ`f�&l��3�Ϝ������>τ���r�|w��e�C�V�O�����[����            �.'/?����=�  ���:P/N;��X2wIŽ�сR$��+#��8������>�v�_4gQ��u���            ��rʊS*��ݴ6  �W'P���'�����Y<����z7���~q��9�Pq�G}@(            f�c�;&�/Z^q��  ��b j\:���W�]qoKߖ�l�eQm��������Q�����z�Yєi���H             �ß��O*��Ÿ뙻  xuB1 5�}���sVܻ�Ǘ���@T�$��;�_zϗv؛�<7�����{��            T�3^F����W�{d�#�|��  �:��w��*�'��k�6���y���_��Wјi�a��U(            f�7t�!�q�7&�����-  ����qo:�M��{�xf�3Q�^̽w<sG������r�[�o�o            @�z���U��,�.��?<6_��  L�P@�[չ������~T�۟��b(��            P�������;>�un�R�I���+K�p  ����N�ce�ʊ{w>sgT�;������Eˣ)�#��             fVkSk�~�����N���I����������
 �zW(�J(��-��,��ي{k7��j�<�b��C5�!�+���7?            P�^xp�{Թ3�4J��z^v^�5��ܦ��p��R &y~�ޮ��M��s/ @�
�*������+�o��z7E�������لb            ��.>4����;jŕ�\�x� @���@�T	� ԰��Ί����l1Y(fi��             f���)~��	  ~a۶mS%PÖ�]Rq}S輦-&{�K�
�            �lrُ.������B>  ���������a��,���R�K1[l�m������            �./�^�߹�w�Go  `�	� ԰����냣�1[L�\'��            աw�7.����;�.��  xm�b jXSCS����p��c��ksCs             �e4??Z�����k�3���  �B1 5�)S9�/�c�-�V\oih	            `f�s�5���<�u?��p<��X����{l�c��?ۥ���v�o��  �oB1 5�1�Xq�X,�l7ٟ            j�mO���0�A�H��G�ݗO�#����h  @]�bj=(��v�x`f�ӲOt���짽?�|q�~�            ��h~4��  �ou���bռUS>���3��uz��z���.����	               �O�X����(�a��:                �%�N����|���D___lݺ5�l�2���r1��                ؉$ ��dJ��I�/I&��ݱiӦ����a��               �n�R�hii����hnn.�`��Klٲ%�n�Z
���00S�:ӝ뎞��T���0���g��j�/�              ��/���ҥK#�����XEwwwlܸ1�o�^zժ�C1�c�1:::��80�
��.�n�QR�              `z%񗁁���닮���H"0��d���K1220[�u(�^���q�!'�l�O�>              ��`z{{K�\.W�'!��۷��zzz�P(�*��:��mii               T�������+E_��K�I�ג��b1�^	�                ��F.�+�_�!�$ ��r��P                �Y�)�_�A���m۶���p �O(               ������Kwww�����/�}2�k�1��#               P����J!�$ ��墷���پ}�D�P(T���5�����                Ը��`��K�I�ג��b1`w̙3'jA*��G��a��P|�oE-�wý              �B)����[�/��������l���D-�`�\u�U�              �nI襫��4r�\���M<޶m[̄8 	�{�P               �����Kww����陸OFrT��+W{�P               �466V
�tuuE.�����Rf���$S(f����8�#��C(               �5*�^��K2������Ԣ�;.�����C(               `'��K|��흈���0�}��z���'�|r���                umpp0���&F.������|۶m1<<���N��}�{_477{�P               P���|���Fwww��������H��&�Ĝ}�ٱ|��`��               f������Ꚉ���0�����b1�׮��-�����!��}B1               @����$������9�L&���8����㏏���`f�                3fpp0���"��Eooo) �<NF___i {VCCC���łb��x���Hϛ7/��t0�b               �=��)�$��_���m�bxx8�=/�͖�/�1��R�<O�RAu�               vK>�������K2���c���d>::����d����~I0I�����舦��`v�               *����r�������0�b1��#��N�_���`�(Ly�J���%P�>����5�]{7F=;zߣ��e�Ǖ�\              ���!�$���_���5!���1�ŋ�F9
�aZZZ��%P�>t���S/��_�����E��D=Y6Y|�����~�cq��
�              ukpp�|��r���[
�$��#������hkk���̟?"�dɒ�>T�o@���8'���A|��/ƕw_�Q��m�7>���ƅo�0��             �֕C0�a���J�^z)FFF�����D�%I&��T*`W�u(ftd4RS�&0��oDj;v2��]_~ϗ��~>.���q�Kc����%-<(.:���~;���              ��|����r�%��ݱ}���Z2`��d2���^
�$�$�R��tttDSSS�t��P�@�@l�MU��fVR0ܺu�۪T���v�vğ��OKA�����+?�J<�환��t����o�t�{Թ�Ig             `6���$��������0�b1�����P
�,Y��t��`��Dy�J����� ԣ������>x��mO�W�}E����1��������ѿ���8zߣ             �Z�<��_��K2O֒!3/�͖�/���L2��� Ԡ�}�sq�{/�e�MzL:��SW�Z��6���^7<zC���]�/䣚�i�g���x���իV�O�}����uI              �)�\.�{�R ����IF2
`f544��/I����d>o޼�>���Ԡ��)������}!.:�h�4���ζ���[>U/�^�������w�g���	���?޾�����q��gN9��6��˹Ɜ�P,             �t[�n]�z뭥H0�Z[['�/�L�q[[[@���P̷G�M�SuZ������9��kc6(����������K�{I���wN���]�x�'J#��<�����S?����I<��xz���_inh�UKWő�'|b�|��qȢCv�<c�����������             �n�b1�����ޑN�c޼y����"���P�:�]�ޣ��/W�E�����/�<N���8e�)��g�y�p�	S��t*��wLi������n�il��{7�=/��ͱ}`{)"�=�]�O��!�m�mєi��sƾ���~���e���G���+�!��oI�T�?z}|�?�Ol}"              ��[n�%x�� �Wss�+�/�(?N"1I,�]]�b ��mO�o��q��S�W�u��ѻu�9�s��eǗF5��� ��;<�*             `Ϻ��{Eb`7�R�hkk{E�<OFkkk ;'Pg��ʱ_:6NYqJ|����Y���M�X������[�w��;              �������~��2�L���O�`�ϟ?���舦�� v�P@JB+I0&�-;.��?����h�4F5��+�2�~��ǆ�             ���v�m122P���D&�L2okk�T*��!P����8����wo����Q���x�Ao�j�Dmn{���_��!�G�             `o��{,�^�c0�dɒ���(�`ZZZ�B1 �tv�w_Q�:W���`����_��W�z�o$?k�]���w�����ػ1              fJ��MMM��$����O�g2� ��P ;x|������|it�uƻ^��8����W��j��X1��+��c�����I����>uk�s             P֭[0�d��W�`�!��<�J0�� �S��6�5�]S��q��������C:�X�? ��wz���Xߵ>�m_��œ[�����?��p�             @5z��M&�)_�!�r�<����-B1 쒮���ޓ�+�_���--1/;/���͏���p�����@i             0��r������mmm�dɒX�xq)S�̛7/��t �C(�i�?�_��             @-�����=!�J�B0I���I���l6 eB1   P�F�����   �UŦb        �����^�L&�����������舦�� �
�   �QC��            {V6����$#��$Q��<�J�k%               �*���b��ť L)Ga��---��	�                u�����)�_^�Y�dIi`&�W               ��lv"���$�Da��T* �J(               �	�L&���K�$ ��_�Q����hjj
��J(               �5���D�%I&��T* j�P               PU&��,^�8�����u(�#~$V�]1��W,�������zK�f��?���`              @�jhh(_�L�IB0�(L�ill ^��C1��=$�w���������v���5���b              f�T*����R��y�<�� �k�:               ;���\������2�L���ǂ&0�<�-*��`��               �$�H̜9s���?�QKKK) ��`��d��$�N�����C1�c�1666����| 3+y���C-             `6��쌧�~:jU6����$��a�d��r �yu���uGw�{��'53`fEw��_��(_�             �M>��Y�ihhxE��)�d���_k               ؉��:*n������Q����+�/��ϟ�$�T* �nB1               �mmmq�G��?<c�!�NG{{{)�R�$#�'!���� ��	�               ��8���㩧��\.�Ǯ���P�Ҽ< S�,Y���@��.                �"���?����7�����}�$�`�L9S���� LF(               �`����.� n��X�~}�c2�L)��`��� L2/���� ��!               S�x����G?�7o�6���h̙3g"3o޼H�R �M(               vQgggi ��"                P�b                 ��P                @��                �rB1                 UN(                ��	�                 T9�                �*'                P�b                 ��P                @��                �rB1                 UN(                ��	�                 T9���{o��X�juԢ�������"               �� ԰Ö��<5jі�-               �B(                ���u(&ד�-�-S>���=�����[�L�u[��               �K�:�����Д�	`f�������_�UI(               �Eu�                ��b                 �\]�b67E!U����o����m��fc㷽������=���               �zQס��|����?�3�������\����                f���                 �B1                @MH�RQ,+���̈́b                ���������c6�                jB{{{G�P�a��av�Vf��                ��p*���_^lll�d�lْllhh(,Z�h���}��NX(���	�                 ���Yg���QG�b                 ��P                0�
��/}�K�]��T*U�/444������L&������;���n��'>1UH(                �y�b�|�i�&c��X>>�1>~?�����񥆆��������yST	�                �q�|>5>�Oߕ���u�e��477��3gΟ������s�`�H��q�>G�qˎ�%s�Ģ9�bn��͏�������gc����E��               �i���M�㔁��{���u��������ߙx.B1 �Q��8%~�����<5:Z;^��ޡ޸�����{��5Ϯ	               �i�B!��������zfΜ9g�w�y���� �q�����s.���]�������q.��?����M��'�>             �t:]�T*  f�$ʒ�������[>00���k���o��o��޺�P@x�o��Ms+�=����нaZ��D^��D�1���sڡ�Ń�`\xÅ�/��K             05�������L&  f�$3<<CCC�8K���󩮮����ꪓ����|����k
� Ը9�s��o������7�#���i�ޅo�0.��˧�.�<�k~��X�]_���            ���v͝;7 `6K�ӑ�f���)r�\f�j���w��������j��?���{�ZB1 5�+�Q1������͏M۵N;������N[$�,9�ߝ�w�B��G�             T& ԚL&mmm����b1����P���}��_=��h����P@�;��gN�w�]�N�u�/Z���7�!�g�Z�X�U�*��po��Z             �RKK�H P���t���F.��j544�p���rO]��C1��G6�ݥす��qA�e�b6{n�(�ީ�%q�3��yv��q��n��k�ՙ�bOjoi��~�X�ϫ            �WJB1  ������)
Q����V\}�՗|�c�̞8]�b>��ӱjު)�����z�~�տ2�#!�wA���k-_�<���Ž}�_#_�O�u�z�[�}G�oJ��d�O�;?�N<���ֿ-2�L�ӾO����>+;vG;��J�[��             �J� �e���1<<լ���S7�x��<�s�M���:P�N8��I�n\{�]�����-?�o�0�x�����z�[q�_\
�\�k�Eg��q��N�H(            �eDb �z��d�����tWW�WƧ��s� ԰��Y�}]<��r�C'|�N����YW�]�]�z��!�z殸�w��V�W�]
�l��               PM���W��Ը�t�W(���p@�P�͏��o*�r����s�t?����s��){1�b����~��Xڶt���tC)s��W             �B!  j�l��gxx���k�}�����<o]�bzr=ћ������̬����������v�UKWU\_��i9��б��1���3��o�.�{C���ܿ.�>���g��L�            ��666V��;���  ������|����l6��P(�7��1~��*244��!3}F�Fbddd��'� 3+�����%?h�K�.���s+������r�7t�!��_6���Mk��G����_s�5q�I�����|ЛK��bo��            �v�/k�f� P��HL�(K�R����'�I��b1u�W��N�?><<|����1�FFF���s�u(��-_�������Xߵ~Z�q��'�t��_�ba�ϟ|m������^GkG��xv��            �/B1MMM��d �����t?�J����#����}|�{����J
;~�=9g2~��c4�ו�{���������.8���b�� Ԩ�\q��M�N�5NZ~Ҥ{��Ѹ���_�5�{����:yc�a�%�	�             �����}}}���& Ԍ��8/����|�#W}�������ȵ��{A�<��866V��v2���7��B1 5j��%׷�o��k�,s�3wƶ�m���u?W��,_�|���V             �_�P�����f����\�x �Ile``��=ή:�3����555�c����Ò�J#��ښ�-��k� Ԩ��s+�o������}���t��g��v�ڊ��E��            �W*��T�>��N�c �Y#�^&	Ì����Ź�;x��7?0>}G̀���t�O(�F�6�V\�잖����;ݿ�;c��t�O�=�޳�z{s{             Ժ��P�yqMP_2�L�츝F~�����'f�����6�- �=o�x���t��]v��T*������H(f��+��|B1 5j�PL�����'?\N&_������e������-B1            @��銿��_�eava<v�c;=fӦM�q�Ƙ~����Ԫ����Q����^���<�P@���>�i��e�O����'��?�K�p_����               �ɤ�駊��L]~�뮻���s��i P�z�z*������J*��c�?v���^x(��dљ����              �6���=��df������e��OO�Ʉb j�d��������%���sN�����tj�4W\�,                ��n���)�O�3�
� v�{����:���}�'�t�C1s��T\��               ��������o�y��t�L\?�N8]���Q�z7U\�l������<���>e�)���Ž��O�>�{�z               ^E��	�
���\B1 5��-�O�w��ĥk.ݭ�fҙx���=��=��)�b���+��uv               �L*��T,���k�O׹�b jԦ�M��wc�۾�{�s�n�b�v�ۢ��c��;��3���K������               v�P(lJ�R3u���u"���ç���y;��p�	q����ۏ{�����|j���{�{1��2M��sUŽ����               �W�=�מ3]'��a��������߮�۸�;�{p��g��wL�>|�����Ǐ��(��qˎ+�b~Y�X�'�>               �3�t�?���i��	� ԰o?����bn���Vt��o_��8���cpt�U����W��ՑIg&=�_�ט�7�SV�Rq}c����               ؙb��?���������?����{o����'|b<xу���>?Z��I�s�>G��>��8zߣ'=&	�|����t;��*���ܽ            ��c�ރ���D�  �*D\jAQD�hA�^�`��n���[w�;���ә�gw��O�Ut��p��#��h�(JѕZQ��E֘r!�<�sH�ےh~O~��o~�����.O2��� �'�d2���-@����M�dƒ�[Է��	b�_�����M<���QY]��vEYIY�:.�~fn�w�y�+��c�����iצn}���3�����3o=               �	2�̝G���v׍�b z���[㟞�������c�M=vj�y(��lܰ��nW�vu�s�z�W               ���K/}�����	� ��?>��q�c���������iצn�g&��ŧ.nw�vomlܱ1                -�b R`_v_,\�0����b��Q�z�ׯ�>�۹�΍1Cƴ;��[OE.�               H���x��8�����%���A����־�/�<�Z���}{�;�{�Շ               �D( E6��g�rfܳ�8w���u�u[����̏��ދ�6k̬������5�4���V               ��P@��س#�.�v������:�K׿_�~|����mkn����O�[߫#On~2v7�               H�T�b��l�߿���[ZZ8���oi_>���_�;��_�ta,8yA�3���1Սձ����7~�m�/��?�w��'3���p~�++               �&ա�����Q�������8�v��;vt~�&R.�%����X��j@�3xL���G&��?������5.s$lؾ!�|gH��{��               �M�C1 ��=M{╝��whjij;              ���                 $�P                @¥:�D�����Y�fύk�ѳ!�!�ny;
����                �T�b�˾ץ�s8����Q��               �4Iu(               ��Z�"��G&�	 �VB1               	Ӹ�1�ox?*�* ��P              @���}�_ @+� ��~C�؁�Fi��X:0z���|>r�\�6�F���رgGT7V             �u��xk,>yq�?8  �b �X�!��Ǟ�GO�ӎ;-�������E};u}����Z�5^��j���X�m}��\�-�             t�~_}\��5��G���4 ��� 8HI�������K')�?���_����կ�_L���v�޳U}s}��ݪX��X�ʊؗ�             ��^��R|���O��$�� �^B1 ��!��ķ>��Xr撨(��ԞSVR�,h;w]�+�|����3?���5             ���﬎y��Ž��� @:	� }z��o�������m��I�ˇ�w��N\7뺸a����K�%�             �G6�l�?�_������b��� ��P@ʍ8*X�@�=���C���.�-��zE\yϕ�}��              >���㮍w��c�����F�޺(�]ک����G���q4T5U px�b R�1g�#_}$�����=vv���^��~zY�ݲ6             ��m�� @�� �Ԭ1��_���1�t@$MEYE<q�q�ݗ��7W               ��P@
M1)�mɿEyI�!]_�\[k��κ�Q�X�M������2�L*C���#��A�GYIY��ѿ�<���b�m�b㎍               i&�2K�C�P�"1�Օ����/��elؾ������$�����FM�Ϗ�|\��℡'t���X̊?]�8=j��               ��P@��z٭q�?q]K�%��p������r�!?�5(��o����`�ج1�bəKbѴEQԻ�c�7t\ܾ����+               �J( Ef���O]���{�����]�����{<�并�����ޅߋS|���L�J���]����               i$��L&n�얶�ٻo\��u��zD��ͪ7cᲅ�hڢX�pi���u����7�)7��|.                m�b R���BL=vj��{k㒻/�g+��#������/��_bXٰv�L19.�xq<�ڣ               i��P�e�.�1��tz��c'pt}���i�9-
��o�M��#���Ϲ�ù������,8*�����/���B<��D������s�V(              �TJu(fڠi1i�N�1pD G�	e'���ΎBv����x(f��q����p���|3V��:���������=��iw~���1q��شkS               @��:���ry�s�����/�����{�˧|9.�tI��s�}�               i"��,lw<��Ƿ�V��$�~���œ��{�>h�5z#              @ڤ:��e#��uz}�B
�F���+�6��qd����8uԩ��=��ظcc$���q���c�i���8|b�4:ޭ}7                -R���S���N�/++��jll������$j�TI��ΎL&��ܝ��Iu׺��Ŵ�5fV<�               �"ա�48{��펿_�~<�'"���|6�To�1C�47���B1               ��P@7mԴvǟx�hɵDR���x�w��_�����:�L               �S	� �p���l�����H���|��P�I'               ��P@6�t@�,��܋�I��;�;(F������               H���!'D&�9h|v����t[j�D}s}���47���B1               ��P@6�|x���Լ���"���|l���FM;h���               =�P@6�|D��;��B�s���C1eB1               ��P@6�lX���ս�bg��v�+�*               �B(�+/)ow���.
EG���g              ��H(�+�]��xsKs���M펗�)	               H����P̾�(EmJ�J               �B(�+�S��x.��B�?p���               �DB1 =X&����W�W               @Z�                 $�P                @�	�                 $�P                @�	�                 $�P                @�	� �Љ�N��O�<
���               �N( �.�xQ�	               ��.سgOlܸ���KJJbȐ!1t���ݻw                 
��.����u��}�L&�w\L�<9F�                 �K(�������1�                ��"s�&L��N:)JJJ                ���:�X�U{��ڱc��ԩS�"1�L&�#���!��m�&F>                �$ա����������KJJbʔ)q�YgEEEE G^sss[,��	�                ]��PLWd2����c���P(nXuC�����'�o�               H��N������ǖ-[��K/���� H�����               (l��T8J3�]����E������+�F�Њ ���LCTe
;|�=p                tE�C1?o���]X�����X�pi\9�� ���[��盞               �4Iu(�p�5�Ţ{�3o??��Qڧ4                 >B1��_���Y~��4bR                 t7��n�iצ�y�̸c��hڢ                 �NB1ݤ��.����X��Uq��ۣ_Q�                 �B1�l��e��������1iĤ                 8\B1��M�6ř��w,�#�:��                 8B1�����X|��x������Dߢ�                p(�b>e���c��u����1�bB                 t�P����W���O���q�iW                @W�!���q���ē��l��/�                 �!s�-[�,^��B,�zy�<��                 �$B1G����z̸eF�<��X2cI                 |���d���q���6�T����ѿ�                 �G(�([�~Y����X~��8y��                �Ǆb���x=f�2#�����7��f                 �wB1	�w����G�&^��R��EYIY                 ��I�e�źw���k�ǔ�S                 ա��^�ѧW��k���͍�Ǎ�Y��#%�J��OQ��lC���                ��UR��o���4pR$֮�����ԩS�O�T���\y��q�G!�ڋ_���w               @g��$�֭[���&�8�8p`                 �#S ����駟�ɓ'Ǹq�                H����fc�ƍQ]]ӦM�>}��                 -R]�k�����QH~�������cΜ91x����inn����ڷ,��               @W�:Ӵ�)����д��C=3f̈ɓ'�IKKKA���.��               @W�:SȲ�l�]�6v��s�̉���                 z&��WYY���1o޼:th                 =�PL�{��x�Gbƌ1y��                 z��"���ڵkc�Ν1gΜ(..                �g��a*++���*�Ν                >�����.V�\3gΌ�'                P؄bz�l6k֬�m۶�9����                &��n˖-���Ƽy󢢢"                ��#�����r�ʘ1cFL�<9                ��"��l6֮];v�9s�DIII                 �A(��ZC*555��UUU��͛c���1jԨ                 �O(��r�\444D�~ΥK�Ƽy�b��ّ�d                H.����f��jժضm[,\�0���                H&���{��"��Ǽy�b���                $�PQ__+W��.� F�                @���&��Eee�P                $�P                @�	�                 $�P                @�	�                 $�P��e2�(..                �����>}��ȑ#                 i�b                 N(                 �R���r��f�������o              �4Ju(���.�Uo>4r�Ȁ�����m�
|��               �KR�                (B1                 	'                �p�ŬiY2���Jc��������A��(d�               ��Hu(�����GNϞ�t�s�c{��                H�T�b                 
�P                @�	�                 $�P                @�	�                 $�P                @�	�                 $�P                @�	�                 $�P                @�	�                 $�P                @�	�                 $�P                @�	�                 $�P                @�	�                 $\�C1s+�ƨ����:3 ���db�����h�5               @g�:3g؜�4pR�1��$�䁓��QG!{tǣB1               @��:                P�b                 .ա����H�               �T�b�j��jU�c�9& ������m6�       ���+N�(�p<��Sq���"       ��Iu(        ����cXٰ��1��        �I(                 �b                 N(                 �b                 N(                 �b                 N(                 �b                 N(                 �b                 N(                 �b                 N(                 �b                 N(                 �b                 N(                 �b�0�x㍱{��H�g+��6<�c��㢡u�sƏ                i#�骫�
"z��W<���PL��~q��s               ��#                �pB1                 	'                �pB1                 	'                �p����5�j�566t�\DM�=v�|                tI�C1���Ş�=������S>��={챃�                ]��P                @!�                H�T�b��ث1�оt�l&�{��                ]��P̊}+��4�o�/8��|�� ~���                ��:                P�b                 N(                 �b                 N(                 �b                 N(                 �b                 N(                 �b                 N(            �����o����߹�>�9�/q(�H�D�Vh*�Ũ��a5�Q��J(h6�:,�/�RUQeӑʂJH��ĂQ;�tjK��R4�����v��>�3�}3�$��㜘�������^?'�mE��5    ��                H�P                @�b                 '                �8�                ��	�                 $N(                 qB1                 ��                H�P                @�b                 '                �8�                ��	�                 $N(                 qB1                 ��                H�P                @�b                 '                �8�                ��	�                 $N(                 qB1                 ��a͛�o����tp����bk���]�˙_                ��Pk�8�F>ܢ���8��;��               @b�bȍ�Gb�4@�?�ؚv�gd��z��ڼ                �P��?������
�_bG�t;Q�'�V                M�                 qB1                 ��                H�P                @�b                 '                �8�                ��	�                 $N(                 qB1                 ��                H�P                @�b                 '                �8�                ��	�                 $N(                 qB1                 ��                H�P                @�b                 '                �8�                ��	�                 $N(                 qB1                 ��                H�P                @�b                 '                �8�                ��	�                 $N(                 qB1                 ��                H�P                @�b                 '                �8�                ��	�                 $N(                 qB1                 ��                H�P                @�b                 '                �8�                ��	�                 $N(                 qB1                 ��                H�P                @�b                 '                �8�                ��	�                 $N(                 qB1                 ��                H�P                @�b                 '                �8�                ��	�                 $N(                 qB1                 ��                H�P                @�b                 '                �8�                ��	�                 $N(                 qB1                 ��                H�P                @�b                 '                �8�                ��	�                 $N(                 qB1                 ��                H�P                @�b                 '                �8�                ��	�                 $N(                 qB1                 ��                H�P                @�b                 '                �8�                ��	�                 $N(                 qB1                 ��       �M��X���r��lD�݌+�+       �LB1        �	���oƫ�?��lďN�(���       ؙ�b                 '                �8�                ��	�                 $N(                 qB1                l��阪L������:����b����                6�w��n<��#�����n��l6��j�0��F#߳�ެ��l����r�r,�c����y���G��uR'               ��+
144�O�Z����"1YH&�z���Y@&��~��ɑ�b�����4�^;��\h]��q�}q�v�׻���                ��,(322������e�V����fee%�B����_.�czh:�c��>��Rg)�\l�@�\�\,4b���Y�b                ؒ�����p>�y��`����y8&�W�w��u�Q+��9X9���P�Bs!��y@&�ݜ�K�Ky�I(               �m�X,F�Z�grrr��,���bV2�,//G�ټ�3F��q�r8��tW�l�l�����\>�?�(�                6���(Ky��Bq��/
���t:7�c��L�w�ݛ>�Z�����|���]�����\�Z8����1ߜ�F��Y�b                �4O���|2��ɘ��;F�=�=���7�T������[�w�sS�2�R)j�Z>�k47�c�^��VkCg�G����|V���b�b�Y���6f�R�R���b                �\|X�0�w����)���/ľ]�b����Wۗ����v��r���Ǒ��|��n���1����F�k���|�=���Jw%��1S��'��,4�;�P                �jw�1�4�ϯ����犅b�Q�#��S�'��'�������;��o�r��Z-����n����xL6�fs�gT��8\9�Ϫz�gg�h�l}6��6�F���?�                ��,�rv�l>�9���*��C����C����/����^�x���x>�:�N�����c��L�^���b%�T��vF��[�c�>��c�=�V�l/B1                l;�n+����|��Eb��7�̣1G&��ǿw���{(�JQ���Y�n��h���R��ng�m��B)��+���W~F�s���i�ğW��5ދ��B����K(               ���i�;����z��Z�92y$ߏN�C㇢Z���r��w��gU�^_��d���Jt�ݍ�Q(ǽ�{����׮�ѭ�lcv-3S��K�K��!               ����Z��^�m>���b����<�O�Ǧ��Tej�gW*�|��ٓ���W����1Y4&��v�����J��g�rg9�s�~���k�řƙ�o�G���#       ����P(Ķ�����.��W��Y�ta)�{� ���Q,��+�W�P������_g       ��n��Wf������=���7Ƭ�c���N���gī��u:��pL�^��1�t����hi4�T��s���b��gb�1���Xh.���ϏP        ��D剘�M�vs�̙x���o�9/f�_".^���W�X�/��O?;M�Ўg��      @J.�\�s�s�X{�v�c2�R)j�Z>�[��\�z5�d��D]����ڗ�YU��c�9�d�"2��`��                �-��x�������<"sh���ϮV��LMM���HL�^h<�R�����|V-w��Z��k�d���>��t�x��'���P                �����N�S��=�����xp���5�k��
���c:�N�YZZ�'���vo���h�=�Mvf�\��'O�ۿ��c����_;q��!             �⾱����|�
�Bz�  �AZj.�O�秛v�ʕ�8}�t��9��/�q`�@<0�@�>���]Ã�d����R���J�&k���������`>�]>�ng��.����=|��?��ɦX,��s�=w��l�z���{���	r�N���K/���5B1        ���*M�v�����������4�+   �s�������w  ؞�������,7�j��^[[ɹ8w�3^r�?�穉����N���oś�F(       �u��Vblx,����р��������,�n=        �                ��	�                �c�J�����L�v����               `Ǫ�j���l�F�Qx��go��                ��	�                 $N(                 qB1                 ��                H�P                @�b                 'C�{�}/~���܊n�                �P����                H�P                @�b                 '                �8�                ��	�                 $N(                 qB1                 ��!�Jz�W�O-                �EB1D�����;�P               �-�                H�P                @�b                 '       ���K�(�J���ŀ�
�m���YJ���o      �O"       ��M�O�de2������ԍ���������,�n#        �                ��	�                 $N(                 qB1D�o`�|^      l;'�x2Fˣ��\�����]�]<�gb�iw�       Ő�       �uy룷b[�( y���W�*       ��I(                 qB1                 ��                H�P                @�b                 '                �8�                ��	�                 $N(                 qB1                 ��                H�P                @�b                 '                �8�                ��	�                 $N(        `��N       �s	�        �n��F�.�����������=v������ ~���b'i�Zq�y*       `��       `ݎ���Do"��������x���}8N�:�f3v�v��B(       �b         ���z(���/��B�;w.    ���Ft:�   �Ai��7}�P        ��w��8q�D���+���    ��Rs)�F   �������F(       �u+��1�_�M�&��}��Gc������/G�� �_��L��\���}�(U@����أ"(F��u��$�S<����x4&�$�ģ�E%�1���B�PD@@iK�]�|�|����.�����\�{��<�����      sy�        ��z���)�Sd�u��4V��Ot��-&M�˖-�LSZU1'       `�'        ���	'����J���       d�        �������;�s�=���       d�        �ҽ{�hݺu<��S���Gc�����       �K(         �������'���^z)��m�F���       �_B1         (777�=���޽{<��CQZZ       @�%        ��z���:u���?>��        '�        �WTT�{n<�����/       ���         lrsscذa��.���?�ׯ       ���        ؎���;:u��ƍ����       �8�         lg�����΋��~:^xᅨ��       �a�        �egg�����k׮��C����       h��b         �c�z���.�(����?~        �P        �v�U�Vq�y�ų�>�'O����        �         ";;;�8��޽{<��QZZ��K~~~        _%        ��H�bF��&M�ŋ       �0�         �͚5��;.fΜ3f̈���        �-�         j��Ύ~��E�bʔ)�nݺ        ��         ��ܹs�x�1iҤX�xq        ۆP         լY�6lX̘1#y���       `��        �keeeE�~��cǎ1y��X�n]        [�P         �֩S�8餓bʔ)�`��        ��         6I�&MbȐ!1cƌ䭺�:       ��%        �&��ʊ~��Eǎc��ɱnݺ        �P         ��S�Nq��''c1,       �~�         �E
c�С��o��/�UUU       �-�        j�U�VѪ�Ud�f͚������ڵK�b֯__'kT               �&��ˏ����4���Fu%�<xpL�6-�,Y���U�T                @+((�A����o��vTWW       �e�b         �sYYY��{D۶m��^����       ���b        ��wKލ��>�L3�� ��;��~hLxaB|���M�YUY        B1        l����ia ��ia�8���⦩7�'�06Tn       `��         Pﲲ���.��#�-�(       ���        `��e@̼lf����1���       ԎP         [U��V���⦩7ŏ&�(�+�       �8�         ���������c����ȱ#c��y       �'        �6��̾lv������       HM(        �m�ea�w����߈?��(�,       ૄb         �沲�⒃/���#�s��       �	�         �`�۩_����8��1nָ        ��         �gĆ�       �/�         �����x`�q����럾       �W	�         ��,*Y��|{���M�lݲ        R�        `�+�,���k��?��bM������       HM(        ��.?'?��G�&��nY�2       ��b                 8�                �N(                ���                h��b        ����m#/+/2Myvy,���v�g7�9j�����UK       �wB1        �ڈ�QT]�擜O��/>�m�ov��;��񊬊����       ��P                @'                ��	�                 4pB1        �ZQ��h��>2�ڵkض�5k��׼��U�E|       ���       �����0�02M~~~ �Vnnn���T       B1                 �P                @'         �Ԧi��ܪst-�Zt���(jRY_|TUWŪ�UQQU�W/��+���Uc��       [J(         RHD`uG�~d�۩_��y��ز�&�����\83�/�O��T�2�����       �B1         �O�qH����ql�c�M�6[�^�V����z?=���lݲx������o���       ԆP         ۽���oT\~��ѳ]�zݫmӶqv�����������o�}QU]       ��P         ۵������]�����{��a�{��d��G/�g>x&        �         �K�
[�u�]�p��~(�Wǽ�������>|a�.[       �τb         ���n�;&��=����dT�Q���㸿|�A       ���b         خ��Q��YF��V�������/ǉw���|       @�P         ۍ#v="�h�n�}+�*��eƻKߍOK>�ū���cu���,/'/��7���M�C�ѱe��ٮg�h�#r�s6i�6M�����{�mpL�75       @(        ������o��u$���:^���x��'bʜ)1}��(�(��}����?����sh��ZݯY~�x����[�Y�f       �7�         2��v��g���Ϳ�����-So������x��[�wiEi��ы��5O_=���s�?7�s�w��I�F�۪�U<t�C��w�b���      ��K(        ��7�1ѥ��F�)�(��\�={]�)[So���e��"~=��q�7����,�r�Ҟ���1�~�� ��m�G��mR��Z�V2"��z��M��8^]]3�      2�P         mdߑ1�琍�3{��8��S���ޏ����$��������z0z������'�9!&�9!���ڡ�&�?���=6�z3nԸ�ӡO����QpyA      �لb         �X����ύ�3���q�}gǺ�b[xk�[1��3��z������x�'c���      ��G(        ��u����N�vJ;�o�}q�}gEEUElKk���Iw��F�������m�G����[�̗�Z_y�=�G��(~��       �B1         d��윸蠋��_���(W��#1_*�,��ƞ�_�|�2 �9?8�����U�Af���F��=6z�^       ��         2�q����m�������)cN����hHJ+Jc��#����՘'�!����A��ӡO����k�;r�#�kQט�r~       �O(        ��t�>���]��U�`Ղh�>Z�Q����o��M��){�"��F]�󲳲��g�5O_      @��         ��İ��R��,�?���h�����C.��-�ט��񑗓*7�'?'?����Z�_<�8~��/���:      ��&        @��S�hY�2��o����h�J+J��7�5�\Sc֦i��۩o���kA���ر���>�{��qh�C�ٹ�      �لb         �8�|`�����q����1�g�=���?������(�����&ߧx@�P�v�ꧮNƢ�UUuU      ���b         �8�w�������Gc���b֢Y�o�}k�vd��-;�1=�I9[�ny4�o�5f'�sr\4�()-	2����      �/�        j-?/?���#�����m��䤼�TUVm�z��k��/|�B4&/|�B�P�.mw	2���ώ���o�g�=ѹU������yM��}N����       2�P        �֪E�hY�22MӦMض


�e˚ח����Z�[�n)�O[0-�W翚�x�6݃̓Ť3f����2u(&�x@�P      d8�         2Jana��l����}�I��ۮy�(�-���� 3|c�oD�v=S��Y�NL�dZ�ʞKV/��-��8g�΃�W�^�s     ��$        @Fi��,�l���ј|���ǳ�����PL�(X�v6f���U1n������S�wN�s���/       3	�         �Q6�Y�~U4&%e%igM���/>h���S�95嬪�*�N�?�뵻҆bF�?y�'ɠu�EA���ʎU�����5�,l9Y9��|Ml��      �/�        j�o�"�s�#Ӕ�/`�zj�Sq��j�����
rR����Ҋ�hL֕�K>��¼� 3���)�I*��L���ϟg,�o.~3�t�S�܎-;�1=����~�^g�摗��r���$�6u��I*+֯��Х�K���8r�#����mvNFb��lݲxk�[ɯ��o?�}��V�l��$a�f;Đ�C������m{D���rN��:o��x����?���k����      uG(       �Z[\�82R��F@FZU�*毝_'k�U��?%b+��C]�,�S���$��<i|�����6�Ʊ����y��<�����ypԃ�M*��KV/���^���ث�^5�WTUDޏSk6W"
��c~��>>r�sҞ׶i�8��!�ۥ_�������q��[�J�j������W�G��#Y[�]����,��������s^�[=��Lގ�����}��r{��ҭQRZ      l�         2����ig��Ū�U�X4/h�v�~C�ϓ�c�v����r��lM<���5��3����_����h׼],]�4�z�9���!������b�٩�Nqð�.���F��yS#$b/:�Oq�.�n�:=���_�U�����"n{��F�     hh�b         �(+֭�ʪʔч�M[7�PL��mRO|~+ׯ��ő���r�����5�Z�i<���qL�cj��r���Έ��1ظ�M��c�~,�v���������L��</�L�ٿ�o�o�.
r�l��MZ�O�c����1r���|��     ���         �TTU��5K�cˎ5f���%�-��ŮmwMy|����ϓ�-3:��Yi���5����D|F(f�vl�c<��g�w��u�f~N~�9�Ψ���{g��M"X����|i����ݾ�\�J|���lT�b     ��B(        �����R�b��q�����h,v�q���篜4~G�~T��j������ٹϦ�����[�*]�
[՘��q��e@���kAMM�ģŏ�*SU]s�͍OK>�E%��y~��ܪs�h�#�s����1⎘�lN46�{]�#1����d᪅QZQ훷O>/EM������nʿM��o98�Z      ԞP         ��O_�A;�q��nĭ/��E��!a���A�7z�贳���&#%�߰>��@���y)����bҸ���ׂ��d�'q�s7Ľ3���|Vc�����8$.>��8��	_��ĝ#��>{/�s�?<�_{���<���N�3%��W����3�=#�3�;Ѧi�����f�x���[����      �v�b         �83�Ly��]��$�He֢YA�ֶi�8~�����L�k$�I���ȸ��ˢ��4�_C{��`���2����c?�u֥=���2KI܎��ȸ����C��3OSv�q�hv�a��u��Z�p������|7�%�ĕ��2n|���É���==���k�\?���      �v�b         �8��}6��E]c���Ō�3��KD:��r�������Έ�܂���?~9��콯]c꼩1w��إ�.5f�����:1�y_�����Ǎ�߸�s�z���k6i�g>x&�q�7b���~%���8ަ{��[�I^���9�ω�o98�^\�5��[g�sF,\�0~t؏Ҟw����c�ƽ      ����(         ���~�_9?��W��wz�Ō�;2��E%��ݥ��[��ⴳ1���j����3mL\=����G����s����������ɑ�/}��������w��-����nߌ�v?*��ӒO��ێޤH�?����c�f;D�ԯ�DL�C~�|�      �zB1         d��^(���k?g�9��'k��FC�4�i��7*��7	�};�};�M9+�(�q���z����?;�g���UcvĮGD�������.;+;���K|�A\2�-�c�q�߯��N�)��8�?6:?��s��m������/�����Jyΐ�C�'�      '        @F���)�m�����q�ԛ��:w�sc�f;��=0���q=pt��co?��-��Z������8��,G9��Yq�����.����i�=zY�W�o�>��?�y�{w�;���윌	�3������Om�>*7�E.�g.x&�9�kޅ_      l�P         ������E�c�N�Ԙ]~���_��W�-_M���Ǘ����/~�b�x������v>f��M^�iw��$$�H�x�Q]]۳S�95�,q�Hz�BeUe�������GCw�~gDVVV�Y��r�㩯C�c�����#��yL��Ⱦ#�	�DEUE      4V����z��X�n]�]�6��į_�֬Y���ӟ7��xB1         d�?������q|�V;��q�?�����#��N-;���<�横�
���m��I9�l�g�ĻOl��_7�xS4�kZcֽM�8l��bʜ)�=�sH���c�t��oM��떧�:7C{M;{�����e��~�8W�PL��u`�4�      ��6lؐ�|z�2��ϡ�T��+WFUU�~?W(        ��uό{⪣��n��՘��ƃ�?�͎��o��q�����-]�4Z�q+P�vv߬�bC�M^���$&�9!N����{nϡ�D,g�6;��UVUƃ�����+���7�s�?7�-�a�t�N��xN£o=+ׯ��&E)�G�v�P     P'6'�R^^��-_�<2�         2VYEY\���qǈ;j�
r��3���6��m�0�0Ɯ6&��R�vҵ��lM�xu)ꒌa�3fژ�^����J�9i��{�|/�����?��%o��Ջ�|�g>x�A�b��w�f���>Q�{�V���9�c�^�S���i�      ����^�<?q�L%        @F3}L|w�wS�"z��>��q��gEuuul+YYY�S�{u�+����ދ?�������gENvN��[�ߊ��o�ړ�L���F�V�k̚�5��}G�m/�ۣ=��v6{��zٳ�֭+}:�I;[�zI,*YT/��\83m(&�     2���^JJJ���"�I(        ��VYU�~��1���#7������wf�Y6'�~���V~z�O���H9Kl���w���,h�1�s���v�m������ď�q��9��nC1���%�l֢Y�����6�KFz�mz���X8���M�b��Z�5RJ��    ��csc/�V���J�޿�	�         ��^���h{U����I9���c[����߿�����c[�~eи���u�]Sξ��l���ݕ6s`��W�^�Βwb{ӡe�����}T/{&���ϋ��{GCԱeǴ�����۾��~�Y"Ӿy�XT�(     ���.�RVV�?�t���+WFUUU�p�        Pk'�����4K���_| �N�ܾ1�`t��������:٣��$*!��W<�8�lҜI�p��-���%oǴO�E�.��>�?�:$��vl�c�YIY�]V�����mӶig�y����d�f;�  ۅ�8?����ǧ-��M�.   �_���|yKzIKܗ�!       @���jE�E�i!
`�j��G�/>�UEVE@c׼�y���Ii�c������L�6sV���'O�$6Tn_���$�I�Y}FQV����j[='_�)�+ ���~���S�9������    3m,�R^^������\�2����b          ��Ⱦ#���T1�G�x����o�}q���#?��`ھE�8f�cb��c{��������o}W������ܔU�EyeyگIa�P     ��b/�[��KIIITT���         �z4z�贳-b��/V�ow����ʴ��Ed�TC��TT�3za^�=�����K;�P�!     �����~%���˸˺u�|���Kb�~����@(       �Z��Ϗ&�M"��m���F�&5�/�������;�t= �a��E�b��ű�(ݐ�"Ҳ�e��۪I�h��*���Z��s�X;+++��    ��S^^S�NM��͛K�.h�b        ��VmZE��v�iJJJض�5k��ռ��V�F�
h��=��clm�ٹq�~��o��m4t9�9u���ҕig�����ʖZ�>���^���Y���?�    �媪��'��{�'֬YSo���.1r���s�=�y���������ˋ�����_�bE4m�4��������:�����?N���H<Ɯ������I|߸>�JD�JK�>X�nݺؚ��:g}����?.����c/���>2t�й��#         PQ�Q�FECS<��Q�bZ7i]'�|Z�i�Y���th�!�OW�N:��Xo�vj�i��E%�     ��ʕ+��k��w�}����ҥK\y��P��~`@nnn�y"��X#�IHcnH?� ��V(���J<��Y�E����������M�����������8q�3_�~�o}��>_(         ��9�^���O�>1���xu���t��ʲ���yM���iڦN��d�'ig{w�;�C�퓷�jc�I�N}�m߾�ӯ����c���     �k�ҥq�UWŢE�&?�������j��kGfggO�8q����/
�         �Ѿ=�۱ێ����)[���˨�����Т�E��a��߈���G�fm�I^��KV/�9��$�/|�B�1��GCU<�x�C1%�%ig��x]JDV
r�d����v�O�}�>�׺u��%o����n�,�Y�-_[����yߴ��}�     ��lذ!~��_�k$�.�SN9%�����D���>�h��?�'_         ��T�[7~�ƴ��L�M�Fb���/~z�OcH�!����o�[�a}<��#qó7Č�3�ƫ]�vq\����=��1�������5<���)g#�����,����U����Z7muiP�Au��럾�v�����Gyeyԥ������?'9�9���c��u��A;�v6kѬ     ��u���ܹs�m��;,N>�d���/^wWL�8qްa�n�         c�cp�H̚�5q�s7�˾���m'ߖ�qlʛE��5���==N�{Z��16.�pI�X�"h|��wf��䥜UVU�M/��J��'Z&,\�0.?��d��_5)����μ��땔����j�+���\ԕ��ue���lu�kA����ķ'F]�ψh��Zs>���k��i��V硘�:����J;���     6��駟���sss�?�adgglC��0a�?�b         �X'�}R�٭/��������R�%�h���w��H�eF���rh��c���o�K�ⴳ)s��{$&a���1iΤ8z��S΋oR(f��yig{w�;�JAnA2TRW*�*�ٹ�ư��R�{�e(&�w�{FC���O��$���{�{QVQVg���?*�,�5�2gJ     ��x�������ֿ���I�&�X������b         �H�9�q��ǧ��-_�?w}��٢�E<u�Sѳ]�:Y�kQ�x����?��
��]F�}���Q�8˖J�.sĮGD������j�g���cp2pT]][��}O��-;F]�����������6��:���C.������w}'�u��q�����So���ڷh��x�S�=+֯     �T�@̫��Z�{z��B1         d����
[����5.>[�Y����S�Rg��/5)�'�{"���/�,
��1J+J��7�j��7�?n�c4ɫ�S.�������O]]�����(�,OF��U��=��n�K�^ڢǛ��l�Ϣ�MxsB�.[��9���s��~��=m���e@��7*��?|>�-�;��9�����<�u|���-���C��z�p�;     6�;�k׮���;u�-[�h ��         ���%�O��{��u�߈�#��}N��СE�������?���AÕ����;2�����U�����))-��oOL��<���q���DUu�׮����Z8+v�r�ӣ�o�E�7[�Z�5�Z�y���;⒃/I9�ψ��;������=
s��$<�A�k~�s7�M'ޔr����|��q�=�m�ugH�!��Y:s�͍G�x$     `s,]��^�?���#+++���         #�㐔�篜��|��W��V�&��V̋%��$�שU�d���G�zD��ߙ�������(jR�v~ό{bkK�.ӽM�8l��b�ɵZk҆b����8�ߙ1v��M~�9�9qˉ���G}IDQ�;�h�״�,���z0���1}��M^;���;��e@4&}��q���N�vJ9O��^�����Z�΃b���7��D����"     `s�\��^��ܹs@C"        @�)�-���r��fTUW��~����=v�c��,]�4��tm�?��d$�u)�y\~��c�Ӯ��!�L�C冠a=pt�ي�+�w������#��[m��I9/P\�P��c�Q������;N�#J7��������%"%>��1��ШO���$����ꨫR�[������~��:oj��mݤu�v�mqB���Y�a}\2�x��Ҟs���$�V�=zY�W��z��5-�uM��ҋ�c��	     �\���wכ�y���P         g@�Q�[�rv����|��q�F�͊!��ū��'7<wC2��_#�+��ul��A�}G���c��g�6;���v����U��֖�{<8�����R·�=<����bU骯]+�ZMĊq�T�F=�f���=��x��Ү�g�=�~g�E]M�|e���W�Ua��ٮgԥD�)tٻ��)�횷�g��l�<�����ߤ�;�������?��ѩe����mXo/~;�w���o<�μ7N�����$�q������b���"����_��s�1%�%1z�訮�     h�����         2N�}R_�zI����:�+��S���D��;��hp�K���,��9<��cq��G�<g��B1�9��I�Cҹwƽ��$B �B1M�&D��|[����?IF@��7K9O�azdߑ�������5��Yk��F�fm�C�ɀJע�)�b��8m�i��E]K�zN���x�{/E�)���΍K�4�;�1eΔx�㗓��OW-ZFǖ�1�c�8&oJ�'�I��m�F�I8�����t��ĵ���L~-'ϙ|�A򺶺lu2��S�N1h�A�o�}��M�U�q��g��      ԞP         g�v{�<��TWW��^g�w�F翜��dd���+��{ψ���hUت����D����D ���g��'^��|l+/|�B�_9?m��x@q�C1���	��_N��מ����'o�UZQߺ�[��򏢾����8��Sc�艑������������mS�7������{�m�0ЦJD|���Q1�;S�w��=�]�v��檪�����	oN  �*�Ϡ�����,��i�|	�ٻ8;�o��3{&�e��&��"�5)!�j�P"�S����E���M��.��Ւ�U���Q$��Z��ElY%Dd_g�Y��y��Й��d�̼���{9�}��u͙��q]��  ꆠ         ��AU��������N��*kɋ�~���j���-����7�O��i�ZzZz���x`�A�1����ծW��dxH2 ��$��{����?��~H�CR!o}�V�ֻ뵻bP�A��#�_k��e��;el*Ԧ�=��Sq�'��	S#73���}�'�Ϋ�@���j˪8������L���¦m���Ί��z,  ���A�ƺ����lʬ)1�O   ��b         hrvXi��sku;�:��5����Gc}���Z;0s�W�O�Q��}�ח�42�t����q_4��>T�t�s����������Ćm�c���D�.���5c��1{ŧ�e'  ��IDAT�/O��D��}D���ѿC�]Z+s�?�K�$J�Jbw�f�8��G��'?����ȩ���_�|����+�[�^      �s�         ��tiݥ��Ek��vF��D����o>��k'f�~��8�K�W���y���hۢm���)U��\�f�Y1'ڼ���܏���.�+��}��qœWDqiq��K���0�xn�sqǩw�~]���>ĝ/��<uM�y}{�����: ���ÿ���5^㭏�J�<��3�$�n�s�����8��������J��s���3      �<A1         4)�陑��S�?P���ku[_��*k�e���{O����L�4(���A�|��s�9U���݀�]q���F�}��'�R6�n�њ/-})���Ձ_��<+�xL��m_���򲘱|F<2{�ݱz��J�}���G�m*��v��֢�q�߮�[��5�=��8m�i1���HOK�rΚ�k��w��?���ۻ�t�n{�xx�Õ��h�G;������*}M��im[�vq|��o��O\c�M}��h��f���2����pz<0��xu٫b      j��         ���٭+��V�-�jӡ=�����oņ�������U��.�]�x�ܼ2�Ι���?|=�j[2$��l�D"���]Zu�-;DǼ��1������O��ز}����AK5��`m�칟�Z2e�=����zG��V�z2P&�Ϊwbنe_~�����Zm���$)�s�?�L��DZ�j�+�����:E^v^jLIYI�+X���.Z�(6m�      �>A1         4)�s*�),.���d�eľ]�����Wwy�@���f�FVzV�46� ��k���j㶍u���++/��k�      �OP         MJ2Ƞ2�i鵺����+Zd���^A1k�VYkӢM�޲:       h�         Фl޾������H$Q^^^+��m��3����m�Gaqa��4��[�  hB�����<sr���<?   ��#(        �&���������̍�E[ke;C�W�w����
�)*-
   ��k�O��i    TEP         MJqiql+�99j=�{���]+��{D���+f��cW%�h�Ӻ�ږ�[      ��CP         M���ӪbP��.�k%(�m���_�����\>3jC��֑�V��~[��       ͇�        ��}���.�]45�[��a�h�"ڵ�����l�N��|��أ����<0���U�����DZ�������]n培�J�EQiQ       �|�       �����R��I$4�����>_>��٩��YC�Z����O�˟�<v���������6�n׻��e�       ͋�         ���͍38�B�^{��u�/欘��k��m�}�*�ɐ��6}����Vڿx��       �y        @�����TY��+bܔq;�����~�d�TY�ǢDm�*(fɺ%      @�"(       �j{a����M��u+hX��,�gV>S�{���Z��e�FAqA�f�V��<6��sG<����ۧ}�����p����2l�a��/\�0       h^�        Pm,����FeE l��Y��ſ���
�������>�B-�H��g�����.���99��)���lò��¿Gm�q`*��23��      �nĚ5kvjnfff���UY_�vm�l�2u��S����re��M�V�"==�^�������m۶Tk
�         �$�a�*�I�ҺK<��g�?��-{���вC��ܿ�A=��)3�DYyYԆ1��T�_RV�>�      @�J�������ܴ��(..���\7Y�lPL��n���S�>$�uv����u��g������         �$=:���p�ѭM�J�}���^����+��I3'�k�_�pr`��=��C����4�[��p{��Uk�_UP̛+ߌ�E[      ��EP         MRqiq�0�����;����va��޲:�mX����V٭�k뮩0����s?O�Ԇ���ƐnC*����+      @�#(        �&����>.<��ط˾_8�c^�T�m�(n~��-zA�����       ��        @�U\Zg���x�ۯDNFN�m��?�[�o���r3s���ί���d{L[0-       h~�         Ф�Y1'&�iB�����H������o�s������zv��mWi�م��֢�      @�#(        �&oꜩ������'2�3ke������+��/�:jӡ=�Y̪�v��       ͓�         ��?���X�vqL>cr���o��Z�eu������[�Em�x��       �'(        �f���_��?va|���E��]k4C���+����~S�9       �A1         4+�Ņ�_�������~G�1��/��r���?�����u�bنe�ܢ�b������gck��       ��&(        �f���4�~��T�Tˬ����i��X�um���   Ԧ����q��W�/.+   �         ���E[S   �JAqA�   Ԕ�                �FNP                @#'(            �j�ݮw��mW�m��X�ni    uCP            @=9e�S���W���b��ɱ;����Ψ�?e֔��	   �A1             �䘁���^P������rP�y�i/��`Z,^�8   �ݛ�        �m���"�GS�%}K,��4��i�「*��~�[27   �/�˓-�ZV�?}��b   �	       @���m��FS�<m��h`���ű��V�/I��      �               �n(;;�N�߾}{@c"(               ��N~~~���z���DP         MNFZF��u�h�毜�J�      4g]�v����y�8���A1        T[�N�Kf�hj�o�@�jݺut�޽B���mKj�^~n~̼df4U�~:(�]�n      @s֯_���Ϗ������o��F���EZZZ@c (       �jK�����M����%�J?_�M�3      �����vX<���u�~yyy,_�<z����               �ni�ر1mڴؾ}{����_�"n��ր����v��                vK�ڵ�1c��}��W'�Z�*f͚x`@CI$�w�q               �n���O�w�}7�R~��ǭ���:u
h �dgg��|"(               ��VZZZ\z�q�7�ܹs�d�����n�=��3��QZZz��ѣ7&� (               ��Znnn\{�����6�z�(//���KJJ��.��.�(9�HOO�C�?i����]9r��m�v
�        ���X�1F�ft4U�7,      ��222�[��Vy�1y��?~���q�q�}��\����H$�d�'�O޷�>����{QP         MNQiQL[0-      ��gРAq�7�ʕ+��W_���?>���زe˿ZII�N��~���馛R�۶m����.]���j>���{�g�k,[�,���S!3YYY����ڧ�EcѪU���̬�u�>���g%_˺�VAAAlݺ��g���Q�>�f���{t��'?i+�����p'�                ��t��9N:�Jk��ũ��͛7�BD>"�lɾ�jɾ��Omذ!f̘�3z��EP                �Jfff���ZM�V�Ԕ�                ����)**J�/
�Y�n]м	�         ����=Z������{cŖ     �jWBf�*��l�*df���Q^^���          �B��Nq�~GF��'��)()�[߸5     ���l�L2`��1�(���֒�

���0h�         �����
�v�I}N����M�8    ��S2`�m۶��3�A3�(�����3���7FiiiP;�    �f�/_{�ݳ��[��gN�����1�w����O�5%毜�Sk���'���E%E��hk����-�j˪�x�Ǳz��X�~ٿjm��qT���5�����ݯ���{��q����=��'�����o�uN��+��?8��x���   �ҳRA ;�UV�8�ױ��     ��d�L~~~���Ά�����#(     ���<;�qp������z�i��>.yY��W�u��b&��w�?�ʲ�R�+o�|3^\�b�%�d�����w�~V2�fꜩ�y���|~��-隧�٩�����n���  @�1=��v9�`g�0>Y�H���     P}�2���A37n����hJ�      �P��=RmT�QqɈKR}�P���=S�N�y͋ƦeV���ظ����|[�D"�zN   @c2��� �}��!�ĬU�     �?�4��!3ɾ���FP     @-ػ�ީv��b������<��@�6�D�M���������   h,w_j�� �U��     ��]	�ٶm��d��?�炂����{�Lrn]     P���L9cJ�x�qœW�_�c���7�n��^ã_�~�p��:�N2�   ���@m8���5�k�ز"     ��-'''�ڷo_���ũ��dx̦M��.���mÆ��#��h]A1      ud϶{�c�y�7��Ώk4��$��p�������l��[�i�O   h,:��#���ڐ�H�S��w̹#  j[ˬ�ѧ}�]Z#��+���i������    ��������V����     �X�vQL_0���f�FvFv���j��֦[tn�92�j~xeD�1�qΟΉG�?i��	q���FYyY����I��
   �Ř~c"3-3 jK2(�w�~EeE P�F��._T'k�~��   ���      ����3�?_�Ss��1�:����#���QFE�6ݫ5�MN�xd�#�~'n{ᶨk�6,�=���D�s�=�{��~#���3&�X���h�#   �>%bN�wj Ԧ��m�^��c�     ��$(     ����l�9+��䙓S!,#z�H��|}��#+=k���q�/���4n�n�طp���`�qX��*��zN���m�7�zT&�z]9��   ��4�Ǩh��> j����      �NP     �N*//��?�j�>um\s�5q�sS�0UI�n;��X�vQ<�Γu��θ�Ҡ�S�=5.z��ؼ}s�n/�S�Ͼdݒ�Ǣ�  �ލ0. �����1�����fn      �A1      �`نeq����}o�SΘ]Zw�rlZ"-&�19��bH,߰�����9ƭ'������o��2��76�~��Z�V�g�0tB���3'G�'   �O���>��	��2~�xA1     @�     P��/����x���c�.�V9�C�q�)��I��Tg��q��xd�#��!_�P�8lb������ѶG�����4sR�i�' ��!7'7Zd���&;;;�����-ZT�|I�%vƙ����td�#�Sn�XU�*      ꃠ     �Z�|��8�7G��;�r܉{�G8:�~��:ۗdHKeA1�{����Ƣ��je;����<��X�n�� hBZ涌�9-�����	�aeeeE˖?_2ʜ�F����Ǩ��.e�e�)}O����M      �G�     ���-���{N�Yߙ���U���c��N�b�/��6,�m{|�?�H�9Cω���z���&�M���)�֒A5   P�N�{jd�e@]�oL���=QTZ  �������z4E�,   ���     �#�z'�x⊸��[�3l�aqH�C��_��}(+/�)3�ďF��Bm��	q��צ����;��0�-۷�C�
   �O���L ԇv9��=��'�>  ��R   ���      ԡ;^�#�uطb@�U��谋�,(&i��Iq�QWD"��\���1��Ș�`�.�?q��J��Ν�
� ����(���Ԕ~� V�'��>_�ˋj��=��N-:@}7`��     �^�     �C%e%q���c�S�s�>'EVzV���>,X� ^Z�R�=�B휡��RP����^�UZ�wƽ 4=ߙ��h�>��=������W�d`@}ڧ�>�w��c���     P��      Աg?�8�ѡe�J뭲[�}����{���a��I�Ŝ��q�����wj݉�&Vڿdݒxa�   �i@������%C��~Y�     P��      Ա�Ң�:gj\x؅U��꠯�iP̃s��N�-r3s?��2�e����q�kw�x����8���+��;��(//   �O����0�����[cݶu     PW�      ԃ��}j�A1��V��ߴmS<4��J�]�v�NŌ0:���V�?3e֔   ���:�u��� h�i�qJ�S��5��l      �%(     �<���(+/��DZ����%�ԕ{g�[iP��^ã_�~�p���7q��J��?�uK   �S2�!'=' �i�O�IoO����      ��b      ���m�RA,:�����}���k��><��x���3�����DL8pB\����^+�E~���I�֒�4   P���c��	��ԱE��}d<��      ��b      �ɜs��I�ߣN�b���b���q��*�&��>}mjLu�?`|�dT�K�����y   ԧû][v��6n�8A1     @�     ����c���e[����,Y�d���m���>L�9)�ue$������#�����Wk��C'V����ck��   ���f h����n�x{��     P��      ��2�e�i�'�m�h���������.���_��
�s��S����;��8��ڽ3�   �O}��; ����c�W�     ��&(     ���ڲj��V9��e?�a.�Ō<&.~��شm��O:����k�KK_
   �O���D" ��1=���޸-6m     ��$(     ����"�E���ԹS�'�2��>ן��c���^��ʹi��!_��6i�(//   �/��Zű����$;=;N�{rLz{R      �&A1      �d[ɶ�[d�OP̖�[��yǄ�*��v��b�:�ѥu�
�e�e1y��   ��tR�����4@M�06������4      j��     �zR��cG�Dԗ{f�SiP��^ã_�~�p��J�M:����/�{,۰,   ���%�bl���u��_���x��g ��]2�8�K�ES4�i��g   @�     �����W��U�l�s����c~�INF��ŅQ_����dݒ�ݮ����a5�='���U��m'�}B���;��   ��4�����- ���.( �ԠN�bT�Q�}��    ꎠ     �_��[�}�����ɏ�-(�Ef���3(���<&Ϝ�}M�����<uM���}���!gFVzV��m�G�=   MI��O���+�W���z���y�y�2�忾mض!��l��E[S�%�[����X�~il(�ԝq�@c6l�aѯm�X�aa      �A1      ��cˎ;�o)��i��Iq��#�H|�?y��~#c����8lb��<0�((.  ��UzZz�6$��9,��94�v{�Wd���)v+6����gƌ�3b�3��_SKz���qP 4vc������I      �A1      ��k��;���èOK�-�,�G���
�s��󹠘}:h�2�θ7   v7�:������/�-�k}][w��>1ՒJ�Jc����?o�O<��c����GyyyPs���|
�����c���hS      �*A1      ��G�;��wPLR2䥲��1���ŏ\����X�?��J翷��x���  `w�:�u�6��T8��#�=h$=-=�~`�]s�5�t������)����_Q=������ANzN�������     `W	�     �'���a}���Q���P�~�푗�������;xl���]���gpf��'͜���  И��72�q�7�}N��-���ծW\9��TK�p&�<�0�QP\T��>'F�̖��8}��q�{�GYyY      �
A1      � y!��N����5��mپ%�Ν�;�BmⰉ�����:.:�u�P/-+��3' мL̞m?y45+2Wă�<��sp��qI�%��?yܱ������_���Ѩ��=���О�����ߜ
���[⃍��H$b쀱�;��=�rX����  Hz��Gbɺ%�;��̉�:/z��   @�     PF�iU���bN���DCH^�XYP����c`ǁ����L[0�E� ��&r#�<7���O@������'L���D;+%�:/<����W���t��M��6���ߎ� �{㾸a��h���:�ˡѳU� �݌0NP �/O��T���i1f���q?   ���     �zp���wX����h(�/~>�]}���P���ߍ��Z��3   �Efzf���q�諢k뮵�fQiQ�ܼ2�oXo�8
�
��� ��l������r�`����h��:ڶh��tKԴ�i�K����N�z�5䬸뵻��g���VDs7��� �����պW,ݴ4  v���������ep    ���     �:��`p���w8�!�X^^�
}��1?�P��!߬tΆ��7�   -�Hę���Nӷ}ߝZ#�2gŜ��r^�]17�\�f����x�ǩ�L;#/;/�?�t�'uA]���m��ܪs��I��ǡ��N��_�=n��M��p}4G��ǡ]��Q��Wc���[f�  �]2 �Ư���V�y�6,�?��s    uGP     @�ڠ���(_����L��4y����k"-�V���~ �� @��27Z�����e˖4����hݺ��K�'��V�����w�zG��mk[ɶx��W�E�ų��W���K�Gmڲ}K*|&�����S�:�#��j#���Ny���^nfn�`�bⰉq�㗥?w6�fwu��ӫ���1:��	q��;ck��  h���0ɀ�dPLM�-X�<{K���m���   @�     P��w
�rԕ;�w��ѐ��[��@��~GVk|�D �yj٪e�g�GS�v�� VNNN��W�|�V�-b����䴉�z]|�oEFZ�N�K^�6�i1u���˛�M�6ECxg�;����
=9��qN�3���;�����`�{��vQ|��oŌ�3�9�Iω�{ ��܌�8��q��� �1I��^w�uq���R�7�kk�ָ����'��m   ��	�     �Cɓ)�q����ҝ��;��j�$/h|���  �!�e�Ż��{���ǖ�����=~������5xH�++/�Y�J�?��ԝ�'�_��h��z�s��94^��/ǩ�N����k4u��9>Zg������������w  @C�ަ{\5��8��ĚTTZ�:�x�S����+   �?�b      �H��;N�c�c������pz4�{8�8��h��j��&͜   %+=�Cb����s��/_�e�_9?v�P�ז��j���wㄽO�o���T�s��ң[�n���� h
z���qP���  h(�s�ǥ#/�o�v��lQ�yɰ���>?|⇱x��    ꟠     �:�<�����:�p��O]���1�Z�5u!e�UI������   ���uK��n�߾��(,.��ն�m��g�6���l�eq�^�E"�����E�����7`�� �A��j����ˣMN�͝�`Z|�ߋ��   ���     �e�,�?����|;����Sw�kL�q��b�~��X�ay   4&�>�?�������hJ^\�b���e߸�K�Έ���u�_2P�)�ux�h�#�m^  �!+=+&�?>��ѹU��}i�Kq���K^   ��5���      u�O�>���Ɓ��ḭE[�.���ť/F���UYO��  ��X�aY�0��������hʒa8�4!n�~c\w�u1v���ti�%Ft MI"��1���/��E  ԥ�DZ�<&n��M��5��z���cꜩ   4�b      jAvFv\��R��j�����⭏ߊƦ��<��  ��l]����ٛ��n��%ۣ9yg�;q�������[N�%����Ǧ.lhjN�sb�zޯ���0  �¨���g'�,��_�潻�ݸ�oWş��9u�   h\�      �Ny��ϊ�|�;ѽM�j���s?��3'   5�y���sc�ظmc4g/��r��cD�k�.�����8��I���j��:6^�p  Ԧ/��r�丟Ĉ�#j4���\w�vw���   �8	�     ����ط˾qD�#Rw�;��Q��V�C.�|�q��\   �����XڼCb>����ڂ��T%�d�	��j����ȢGR��  �j����գ������Ѽu���goN�,,.   �q     4+{�W\6�j�M$ѶE��#o���)�v�}���Q0̧�w����?��z��   �b��?= ��>m�ā���� ��ի]������#�i՞��hk����q��o��   �=�     ���]�����6��[��/~>   �/6�Ӑ�?  ��q�	� vJ�6����W�y�W�]��=3�k��&Vn^   ��EP     @),.����9~��OS�  ��I' 4�w;<���+�� ��h��.~0����ߎ�-�=���,��P\���h�    vO�b      jٚ�k����~��Í   P}[tL' 4i���L���� �i��2.�����#m[����i�ť�]�W�   `�&(     ���o=�y0��(,.   ����iNo��S�������V�-  �]fzf�;�ܸ��k�K�.5��ϥ��˟�<�_�|    M�#�      ;a������7S'W&O���|�p   �EY�Yqrߓ�9i��:��yt�u�_ �Si��3xL�x�ѯC��MǼ��bꜩ   4-�b     ��I�l޾���܏���~l-��L���j˪�^���_�5[����Ҳ�شmS�y�u�^�=�/������W���ߏwW�[�kX��]\�k8���ј�+X���wYy�N�����h��V   ���{�r�@s3~�xA1 ����?*n9�ؿ��5��t��������;}�   h��     @3����,߰<F�ft����G4�fNJ����Q'��k��}  @�;}���h; ��_�Y3' ���О��O���8���5������n�_��WQTZ   @�%(         j 737z���[u��Dz�m�6�D�n�7FIYI�ܼ2��_�A��08���K�\�0NP 4S{w�;�}M��ol��+X7?{s���_Faqa    M��         �B�6�cԀQ1�ې8������[�W{~��Ϗ�?x=^�����޴X�iEPQ2 �9;��Q��N��pU  �C���q�QW����i�՞�%���;n��M��pC    ͇�         ���z�;7N��ؿ����V��v1���TK*//�7V����h���������-:đ{ �Yz"=N�wj�zޯ h�:�u�����d�%���]�yť�qό{�ڧ���6}   @�#(         >�>_���8f�1��H��m$��mH�]=��x�'Rw����Fs6�ߘ�L���.�yx������( ����c���������⡹�O^�,   ��        @��o�}���n���j�n7=-=N��	���[��e�_o�v47iqrߓ������sT<�� �?��������Y���a�EeQP��%5��b.����nݛݮ[ei�kj7���e�e��i)nY�"*����"�o�����?�����03g����<f��s��sf�0G��: ��~mv\~����   �(        �6)]P�|)�q�7�0��YK�,愡'�7�f����7jjk��8��qQV\ ��s���( �w6��;.��D2��1}�Dk�f���ڿ   �4�         ���l�3~���Ƹ�㢥(�+����1q��8�3��-�F[��! ������w�?�Y @�ս�{|��Ek3c���r��    ���         ڔ�F����?�u�-ё�s�}n��ӓ��w^�\6��8����>����kk�      �HQ         m�=��>�Xt-�[�WTWĒw�ĊM+b�ƕ��jkl���5��.�]��dF�g��1���(�+l���:(����}$^Y�J�� �u\���{�~/֔�	     ���        ���:�E��n�kV�^@�*))�n���/�5�K�>ҥ-_�p�Jb�o\|��ؒ��eO��k^��ښ]>>?����C�O���)��=���ٗ̎�o9<�\�f��E���~� u$�����O^�I      l�(       �]��=*�h�����$~s�ov�����:�YtO�䩟��?���ݾ�t��＜w̿#�yq���Ӈ~:�qf����۱o���_Ǆ[&DEuE�3���� �~g>+��8-�o	     @��         r�-g�#z���ۤR���ٻ�~5�X�F�<��ښx�Շ3cp��q�Ǯ��F���ǌ�;&��/ߍ�ͿF��K�ř�� �\��nq��G�Co>      i�b         �i��{l\x��z����䙓��%�ƞ���%1i��8q؉1�iѽ��No{�a����'�x2rA���{q� ��}|���      �S       �.��[�����#׬]�6��h���덻��W�Vg�[�W�?��z�9oΉ3��+7�������A�=(f]8+��S�m�D���Ę��DMmM�v�� ��Q�F�����5/ �;��w�W=pU�ʚ�    ���        v�����&�f��W��5z��1�c���t��ן��o?96Wl��������[��?�`��?��ی�=*�}N���]њ������9�ǡ�b  �l�ښ    �(        ���H$�G|a�믮~5N�vZ���l�~��8�'ż/̋A]�{��'^3ΌT*�U�����o     �)�         '=���kd�k�5�q�gf�YZ��[����ώ���T�'���_��9b��
       �E1         䤳G��ӵ�~�ㅕ/DK�������9����w=�q)�      h{�         �s�yq��׻�nۺ���%����qE��u��qF�������       ��P        @��{t���ջv�[cSŦh��o[�ν5.;�:k�:�zϭx.       h;�         �s��Nצ/�������-�I���      �6FQ         9�~��;�x��xi�K����x���cX�au��E1S�N       �E1         �!eC�b�њ�i��-�ٷ۾   -M������w   h�b         �9�:��w�鷞���eO�E�.�3?���   ��b\�q�c�붭�)wO	   �i(�         ��F��=�]{m�kњ������+
�
���*   ��l/�9y�ə�3�   ��(�         ���+�D"Q�ڛ�ތ�dg�7�HFiai��  `O�{T� 欑g��98   ���         �SJ
Jv��ڊU֗���ZqAq(�  `OR   �KQ         9���h�k���њl�ܲӵ��   @c�kd|�د*�  �f�(        ��RUSU�|*���(���;	og'   41   в(�         ��W��;�>����$6Ul�֢��t�'�m��   �F�W{��   ha�         �S�o[�T���:wjUE1��[��Tmlض!   �]ú�c�=&�����^�{Ei��(�+�<�]�um���՘���x���c���Y��в�q�I��i���[1��   4E1         䔊�xw˻QVZVgm`��������ا�>�ί޼:*k*  ��R�WS�N�;��bd��;�]ג�1��8x������̥cnz��Ţ_d
T�G��������O6����}��o��/�   @�Q       �.;���(y�k6�o���]���?�UpT����.OV=��7׽YoQ̐�!���b�n��;ߚ�n   �5G�sdL�45��ݭ���=6�����	��)wO�7־�O�I��\v�eq�1WE�v�|�邘k�6~���\N   4��        v�ؼ��)�)r�[���@3�;�w�O��3_��ޭ���W>�9A��wH�䩟Dk1���z�[�\   �;��.7�zs��%[�<<����8�g�Ŝ7���v�:�����Lh�}<���񍇿��x    {��         rγo?qp������&;{���/
   r�g�6n9��F��^�=��q���WW�Zg�̑g�m�n��ŝ��.����k��/�>   �=OQ         9牥O�;?�lhf����h�u���w��7�   Z���?��M�ݩ�S���{������_v�eq�I7F"���y��ŵ_��@    �GQ        �,��4���"?&h��g���;��ɼ���{�q�C�DKwށ��;�f�X�|Q   к��O��i�'����z������鉛2�?s�g�['k��O?�����W��*R�T    �KQ        ��[�nѻ�w���� �Wǎ�_�~u��k�#�4</}�ڬų2'�}�'�d�$����h�
�
₃/�w��/�>jS�  @�v�aǐ�!>���<��v��_9�+���8F�?:�G�t̼e�2%���`    -��         r����ޢ������G<�\pg�T�x^��ԯ޵�?��   �u�K�ťG\�Oo�|��c�1������b��5QS[��ѣ}��0`B�8��8{�ٙ���t.���8=�x�#?�᧓������_�{ߛ)a   ZE1     9�}O�k&\�UƼ��?^������K�|)��G�=����0��џ��G_�U�C{(.���.;�8��Y�����Ƶ�v��?rc?���ro[t[�p�w���q?�	}&d�����;�z��f�4#F���*7��M��ѯO�u�4(���>�٘�|�s�?>;�w�*��.�E�,�a�)OE�d��rO��)�֦�޿����S�G����X�u���{��3�0�YeV�V����an����ݧܝU�-+��_���\��6����%��Y����ܱ���oO�vV�/�}9���9;�M:)�r�W�ʭo��������\V�.}0���U;�5�^v�KwǍOݸ��uG\':)��?����[w�����㨽��*���w���ɺ�����q��e�{�S��/^��s3O�û�*��=���2  �����k��>]����壿�x�QUS-M�ľ����޵�	��_�   �nG<���ۥ�`����q�7Ƕ�mu��s[��̸뙻�k�Z������X�y���7wZH���bs|��/Ǐ����}   -��    ��.�(�+�*�����(��oA� ���^m-=�mn}����7?Q77��mn���>�]~���L$��&!7�cn"��:3��ޥ�s��$߻d��.�n�N���"7����ސ�{|����^��ɺ���yS쑍��%��s�oHk�� ���M��-�%��/ߩ��_���s�?�9ᮥ��_��eC�]��_�"�m   h�3F��ӵ��I�'Ŭųv9/]��/?�����[��.���a%1O��dL�99�\�f    -��         r�O��4�|̗��^��]s�5����/��b@�q��W׻��bS�:��   ���8x�N׾�ǯ5�$f��ښ��o?#z��	&��1�������ʚ�    Z>E1         䬍��Go�o���:k�:�]��G�����t�-�Hƴ�O�E�]��7�   Z����=�׻�x����c����������3��?G"�����\83s�T*   @�(        ���ÿ�0.9��mp���םx]\��+��]����#�>R�����'n
   Z�a݇e�B���(jS�Y忴꥘���8n�q;���5K�S����   he�     ���c۶mYelܺ��ܦ�M�*w㶍��n�'wk��鏹Ir+��nښ��w[e��7o}����irKR%Y�VTUԙۺmk��e���յ�;\O��d����r�j��έ���3WQ]�un���A�c�߻[�~�n���$�M�Gn,o�=���M���s�5�^��i����#�_�:���#K�f/��K6���  �}���WH��G�}5�+&^[����9���/��'^���Kg]�y�  @�7�렝���_6�}ܳ�-��ʃ_�<_   ZE1     9&]^��+~���dM�����8��ߢo�=�1�Ϛ,7�ڥ���$�5�ho�ֵ7�#[~nS�e{r�l�� ��<���1�;��0����tqgsZ��1������\���    7t.�\���5Kc��Սr����Z�����   ��Q        @����磥zn�s  @�о]�z�_X�B��ǋ�^��&�:k�_����   �>�b             ��E�_�uM��Gumul(���;�Y[�|Q    ���            �=dgE1�76���߶�ޢ�e�   �:)�            �C
���W�T6���,��i   �=GQ         9���,���1}������c���   DTTW   �:)�         '�1<n8醸��k��W����o��mT�V       �6�b         �i������OΌ��ǌ3�'O�$���$       ��P        @�ѻC�b�����b�ܩ1s���\�9       �%S        @�4���[��So��_�?S�ȒG"�JM�6⡇��7�ѣG�5* rպu��駟���۔�      i�b         hӊ�cҨI����W���ϻ=��_4�DM"n��z�q��)�r��o��K���Dt      E1         ��в����~=�>��xtɣ1u�Ԙ�¬���       hN�b         �95�5QUSy�u|2��c�=63Vo^w>sg�>��xa�       �AQ         9g�ֵ��q�����1����D"�ح��Ҳ��_̌W���O����i����   ��r�����>6Z�ޝ��w��N�����K�)�~uv��؍   4E1         �u��eJ]�#}r�#Έ)c��A}����=��'��m�n��bƂ���DMmM   @6�w�Mmt��M��b�    ���         r�[�ߊ�=���ؿ��1i䤘<fr��u���k��.&���oox;�|�θm�m����       ���         ڔ�+g�7�F�0>S�r��s���l���t�WL�".;겘�朘>z���]��rK       @cQ        @�T���?���̸�����a'����pz�%���L$c	�q�I7�ϟ�y���że�       ��(       �]VZR�E��k���h^���QZZwɯ�3�VQ]��pof�����ѾGVy��;�%�]�/��rL{zZL�?-VmZ       �;�        �ˊ�����(rM��h^�����/��D�vú�N�!�;�x���b�ܩ�B����       �]�(         v������^�=�=���Zҵ���%���}�͌��V�����gO�,^~��   ��H?�����E�W.   ��(�        �]�h������ť�.���&�E�.�S85
�
�ճ}ϸ|�噱��bƂ��v��    ����͙   �P�b        �e�+VG�K�YW�.�浥zK�*_Ug���"Z��ښ�+��G��Nq���c��)1���H$��wLf�p�q���b�ܩ�ȒG"�J       l�(       �]v��k#'�@3{`��g����m�3�.�1���8g�9�Ҙ�]68�(�(&���o�+f.��ι5�X�F       ��         h/��r\��5񍇿����c&�y���J��w��㊉W�eG]�.y4f,��Z���Z�5       h��         @#�M�Ɵ��sf\:��8y��1e̔8q؉���kPV2��c�=63�w���E�dJc��       �-�b         ��l���\����ש_|b�'b��)1�lh��:w���]�Co��~5       h;�         ��l����#�̌1}�d
c�}n���58+��      ��EQ         �a�� 3.��8~��1y��8��S�0�0       �>�b         ��T�T�}/ޗ��;ǤQ�b��)1a��       ��(         Z�u���mO���~%�y�7c���       �)�        �f֯S�8��s�3�>��
       � E1         �:u�S85&���>&�D       ��(�        �=$�H�у��)c��#Έ�
�
   ږ�z�}:��3�z��X�|Q��M�-�yf��{��'.��%   4E1         ��F��� �;��աWVYsޜ붭   Z�/���������Z<+N��iYew*���.��rKT�TFcI�v.�\g���$   ���(    �����K�5����a�غukV��'�07�thֹ]���ݧd��s������+�un���ur��w�:w��}��vNv�:wX�:�%���sGu���G�5�Y��<6���G��TlMe�;���_�����I�d�{dّ�������_>��A��cKՖ����f�[����PV\�un�*Y'���Y禿�>�;�Ӡ�s�j���o?�I���%���M�<4�^ַ]�:�=
zd�;�dP��.�.Y����`n�DǬs�+�/�zW�0W\[�u�莣c��^;NVFl��r�rh�k�/�����1�ݹ @v�'�M5)���L�*k妕qϢ{�O�4�[�\   @}�~��3%.t���㗋~   @�(    ��]2�(L6�cذaCVǗ�w�ܐ�5zn߼�M��/�_����n��wȾ��{`�3��s�w�;��>���?�;�|/�2��Sz��P��Z"��3��Qgn��-�����_g.��m�'~�Ir��g"�ʃM�[�ޥ)rK߻4EnS�
4I����1|��F��~Lf4v��N�3��s��rDf젦i���m��e�/ۓ^���� ���.�]|t�Gc��q��EA^�ng����c�?S�N�{_�7�j�      ��KQ    �@�;���zC:�D��>QZXE�EQ�_�lK�.�T*m����cŊ ��o߾ѣG�hKF���?�b�rU�VEEMEl������77���xf�31����� `�ڿ���r��s����Ҳ��^Z�R�1���6Z�ڴ*        MQ    ��z��S���>4z��3   v� Y�����#�F��V^]ϯ~>�������Ǧ�M 4�>��Y#ϊ�0F��Uֆ��g3̈?���       �R    �h���b��S�̡gF���  -A"�Z����8����q���������/�y1 ����=e�Sbʘ)q°"?���W���9oΉ���]��[*�       쌢    h���q���a�D�v  �)��k�<>>:���7ϿYa d�ʣ��;ϻ3ڷk�U�k߈iOOˌe�       �
E1    ���OҼj�Uѽ�{   �	�D"�{x��3>�}�޸�cS妀ݑ|����5�D*j߻ �'���%��̧R-�����������q���b�ܩ�ȒG2       4��    �C����?r}���   h�D2�rF�����+c��9uI�%�)�)r�[�oŌ�.@�7!�(���|u�:�U��=�8ڷky��7��91��i��g�7       �.E1    ���>*n�xS�.�   ͭ��,�?5n{���3?�T* Ж�%�b⠉1e�8��ӣ�]iVy+7��{��ϻ=-_       ��    @;�����ߎ����:>}�fmm�����[  h
��7�����+�Hd�����d�3�'�_2���ip|��/EU��9 mϘ�c2�0�>'��v�*���&{���:wj��½�m      ��)�   �&4i褸z�Ց����WSS��r��1�.�| ��.�{����g{aL^^^fl/��g�plL�����ß���[ r�����Qg�'�|"u�u�K�^�;����O�U�V       4E1    �DNtJ\3�]:93]S]]�y  �;҅�ۋ'�ҥ1����Tsh�C�o��0*k*>L��K^��56l�yG�.u����.�"��>��Y#ϊI�&ń"[�7���.�ϟ�_�       �'(�   �&pD�#⿎��z2f����*sB'  ��RvH�W[[���[��.�)((�Я����L�N��#��9
���(���\SRR@�*,,�����/�廕��̏�0�?��8b�#"�Hf��jS���G�g�~�}ᷱ�j[       ���(    ـ��;G'
�;�MMMM�M'_  {B��2=҅1��w���G��|!n�s @k׹�sL�45뜿o�{���]1u��X�fi       @sQ    ��0�0�3�;�W�^����a�1�  �=-]�~>�.���˫�6���xz���� �V�W��}��f�/?5��{       �OQ    4�+�2�uV�Z���tI  @sJXVTTD~~~�0惒�d\����_��*7 �%�� Ss�;c��5       -��    h$�w�?&�T�Z� &]  �R������F�v�"�H�֭�[|��/�5�&  ׭ݺ6~�ܯ�G�Q,Z�(       ��R    � }R�5���d^��������	  ��&]S^^�)�I&�;��5��������W? �kjjk����s�ƽ/�U5U       -��    h'<!�����	��/  Z�T*�)��`YL2��K�^�z�S ���w^�iOO�i�ŪM�       ZE1    �>5��-��   ����b��#�F�s�� h�6�o�Y�g����c�k�       Z+E1    ��#�û�a���2jjj  ���^STT�D"3�~{Ѩ���? ��l���������ɼ       ���    �Ҥa�v�^]]�   ��?��lw��GD�α�|] @k��bs���]       �BQ    d���4�s���kkk���2   Z��󚪪�(((�\/H�)�O��/L         ���    ����������+�  rA�(&///��d��	OP        ���    @��������Q[[   � ]�YT��Ř�w�?��c[��         �y(�   �,�����T*UUU  �+�E��B����(H�!��'�z"         h�b    `7�ܫg�ثG���ɓ�  �\�.�LŤ�� E1     M�#�|$�_:?����z�o��q��+���20   �=OQ    �};�����  �\�.�L?�I������    �R��N1��&�ާ�>   �~�b    `7�<(�6}�d��I  �\��(��� �IQ~QL;%r�=�����       m��    �M}J�dަO�  �U����ѣ�G @kҾ�}�z֭���x�	E1       m��    �M{����	�@˔H$�C��QTT�ڵ�d2� 4���P555QYY[�n�M�6eF*�
��I��         �GQ    즒�ɒ@˓��={������� �<����� S�.�J����ձjժx�w��5�t����s����(�+�ʚ�         `�S    ��(��	��u��=z�� ���Ϗ>}�d���~;֬Y@ː~�J����DQ        @3Q    �)}�dMMM -C2�����G�.]�֭�� ����lٲ��]@�K��$޻     ��g�~&~�藑��-�   @�Q    ���VI�������FIII �;�u��ڵ�%K�d
*����    �qL�;53    JQ    ���� Z��*��Q�۷����z �KQ �M��y隥њ���;��       ��    �n���	�����ѡC�  wu��)z��+V���T*�A�/ hm�n]���M��Nq���c��)�O�}       �S    ��6U@�*))����  ���b֭[���4E1l�����&�Lм�D��K^"���J&�q��3�0g�<3J
J       >HQ    �&E1�����9��ܗ��������z �CQ�u��%:u�\Ӿ}� �Wqqqt�\w����\5���8g�9�Ƀ?�;�       �0�b    `79I�Wii�9ژ�;fN޶m[д��3
3 {��;�9����8��!����|cl��{1      @[�(    �V��W ���K:u�(���L �=�D2�|tL;%�yf��48#]�6��91}����pfl��       �-�b     h��E �=��Ŋ  ��в�q���c/�]�VƲ����w�ԹSc隥      @ۥ(    �V�]�vQXX �=%%%���555@����(�/�\�i٦ ��_��5��2��|Mm��ݯcQ�8��Sc��q��c"�H48cc�Ƙ�xVL�?=Y�H�R��%��T\u�U��v]�v�\֯_�]������     @Q     �O�(�����(�l� 4��6<9ic ���o�Sk���(�H���3�0�t~�U�W�3jS�1��9�r��g��͑��vX �u:tإ�p�s�      �b     hu


��+?��� �eR6$�;�`�1�ˀ��X�~Yܽ��:wj,]�4       `g�%     �N"� ڮd2  �\:u��8-&���>f��;���1k�>z<��H�R       ���         ��D2��)�9���c�½�Q���9o�ɔ��\836Wl       hE1         P�~��Ź�vq�2p�2��_w/�;�ΝK�,       �]�b         ��ס�C�v�i1y��8f�1�H$���|c�Z<+�ϟ�,y$R�T   �v�=>F��h��q���   �4�         Ц%�?`|��ϋ�v�ΨM�Ɯ7�d�af.��+6   ���N���8rь3�   @R        @���#��>�ۻu�w������,[�,       ��(�        �M�O6�O�6�o�Y�ge�aY�H�R��y<��c������M�4)�;��e�^{m���K>n�>}�m���=�P�����+c��ё�������n�qݻw�[o�5      ���?��ή�>����̝=�d&+� �����BYd���b�
J}���
�>�}����>�"}Ԣ��He�� �
��HX�0�d��r�9c	������~���5�s�����ef����        `zs�qϳ��q���N�v�c/������~���1ٵ���c����dr�����ٍ�����     `�	�         �nԵ����4��qC       �X�        �ݨ)�������o����uK       �X�        ��p�㊷^�=��~W�{u���i<       ����������Ҳӟ����۶m۱.7�}�         � ����I��������o�W�sU�y~M   �@}���c$�~�5�
�vY~�΍U�
   `Ϻ���zihh����?�^vD^����tww��c�        `J{���hlo�����gz�����q����?������       ��+c/����V�%	��r���b       �I&�	 �����^7��)�ZzV����8uɩQ�7����X:�p��'��$������� �{G�jq       ��Pc/MMM�����P         S^gwg�zhU:�V̍s��<⃱lβ�QTPgxF:^l~1V�vU|��_��^x(       ��W_�����Z��dYr?v&         ��B��;����V�����z^Ԕ�x�9s�c�~,��[�Z���v��Q�V       ͫc/����V𥡡!r�\0<�b        ��d�y1ټ�})~�w�΁�9E�첼��vC�1V��K2.��8s�q�����%�FA���Kb3ɸ�W��a����[���;       FK{{�N!�$����Kss�n�3>�        0`��GU�*&��0����軽Zwf|�T:�;b�C�ұO�>��C�<�q@�1PEEq��s��|��q������Z<��      0P]]]��2�R__�,߱mr?&6�       v��� ��K"/W���t���".8�x�!�iE�<G���Kұ���q��W�w�|7Z:[      ��v{�1�e��KB0�񚺄b         `���˅߿0.���8s�q����%�E~^���Hb3_}�W�K+�?z�G��ߊ[�%zz{      ��{ijj���2xB1        X~~~d3٘l

Fc-///�ى�����#V=�*�*��y��~�����x���8g�9�x����ߎ���?⩺��=����e˖�v���>uuu1-Y�$jkk�]��|�=������c��]�z��hoo���������~�566��?     L<�|���Oǫ�'�&����       v��d`w�Ϙs��d����ؚ6mZ̝�����ގ�'cBI"/W���t���".8�x�!�iE�<G���Kұ���q��W�w�|'Z;[��%a�O|��]�W��w�S�����8���]���!�.�:���?��ݮ���?<eC1]tQ������m����]     0~$���k���O?7nL�.���;E_��5��<C�㸭��$�{<�c�r�ܘ�k�یB1         0B��˅߿0.���8s�i4���O���Il���j|��/�MkoJ�1w<yǄ9P      F[������;����a�?y�o�ʕqꩧƼy󢰰0���<_CCC������*�3���ٙ��&��e�nݺ�ߺ��b�s뮾�?������O�����        �����Z��y���Cϋ��X\�x�s�dK���cɕKb��u      ����E|�k_�@L"��|�#����aT��\.wP��W�X�n��o�8��^��P         ��皞�+ve:V�[uA��!�E$     ��q����5�\3b�_z�q�I'E&�	a�r�܏���k{{�_�{�=�B�         #��[~�����2�8��4s��':�      ��k��뮻n���+���e+..������d29�         &����XX�0&�ј�5��}��/޾��Q�-	      ���׿�U�V������Eb3�L�7�|�}�~N(        �Igz��x�o�
      `r������\.7"�WTTĻ����������M7���                &��n�)���Fl�O~��f�XA.���b                ��~�ӟ���˖-'��               `�y��c�ƍ#6�������DV(               �	g���#:��0��                0���׏���f�
O�b                �p���Ft���Ҁ�D(        �I���>��☬66n      ��r�\�T"        ��������       LB1                 �P                �8'            0J>y�'����>"s�dK�]~��W�%'\#�Go��n�,   ��!            0JT-��V��>���oT��v��    F�P       ;�d2         �/B1     쵼��Q�_~~~ 0u���?w         ��@(    ����f'�� _��         �"�     ��h�@_P��m��l���         ��h    `�������JKK��k4d2�Q�9         ��     �Z6�MO�ooo�}0u���G~~~������M�yyy     0\x��X�Ъ��~���   ��     �Eee娄b�� @EEE444��~��\.     �ȸ�ޫ�   0XB1     ��3g��͛G���d? 0k֬����GMMM ���i�QY<��eee�����~�E=E       �     0L��l����֭[Gl���QRR ��̟�D���4b�H�dS�-�L& �S�-L��l���|O�P_�_z�{       �    `͞=;��룧�g��NNX�;wn ���O477G.�����g͚  L\3�gĖOo��jɕKb��u      ��!    ��),,�}��7�|��a�{��Q\\ �CIII̛7/6n�8��&q����/���         `��    `XUVV��ٳcӦM�6gmmm: ��fΜmmmQWW7ls&���� �k��Ɩ�-1�lh����ܱ9j|h���{�            ��g�}"???�����+	 ̟?? `w-Zyyy�u�ֽ�k��1cƌ `����WbR���}��/��2�~��   Lv���(*(�eyWoW�v�   �G.�K�H���M�x�<����0R_���w��<&�     F��ٳ#���ƍ���g��O�LH�3I( �$	����!�qZP.����      I�|�?ǅG_����1V~ce   0~l۶-�l�2��ihhH�5����eee#�����t�G�LfP��     0bjjj���2=i���^�����c޼yQXX 0P�f�J�$������'y�uƌ1w��Q{#         `(�b     Q�p�3gN���ESSSZ���r�&9I���$��$q���� ��H"c�/N���\a%���;�����K�:�De����         ��    ��HN�Ob1�HtuuEoooz�~6� NItl����H"1����ϝ���t$�2  ��/���x��a��c.�UvY�?O�Oܾ��!�[SVs��       $�b     �0 ��$
��  ���������a�����7s��wŕ?�r��.�Y,      ��    �M˟۷o��v������#���'  0��-;::����[�����~JJJ��wٓڢ�h��         �>�    ��Es���u�ە��G^^ވ>����hii	  Iq QDF^[[[���#���s�Fii��[Z�4ַ� �������û]___S�UW]�\sM��z{{^��[o���k��7o�Sե�^���f�~     �H�         &�$v8������!0PI( ���h*Gr     ��'                0�	�                 �sB1                 �P                �8'                0�	�                 �sB1                 �P                �8'                0�	�        0`5y5��M6�3ۣ�����Ly�Λ����\ol�m	       ��b        �w�+�rU1�l,���c������첼;����|       �T'            0��= .9ᒘ���Hܴ��    F�P         0!UVVƒ%K}���ژ�-Z�\n��+**
��9s�鿧����2�̐�.ӧO ��:pցq�[����[��%  ���������3`<�         &�+V��]}�#	��+W�����?��     `|������l�0��        0`�Օ1+;+&�m۶0����b֬]��t�vF<       ��?�������[���B(       �+,*����l
[Q\�����       �עE��Rl޼yD�_�zu�r��d2�@N(               �	��o~s\w�u#6����c�����/�b                �������-�����#2������W�0�z{{?%               ��TVV����\�;�O<1`}��ϾK(            `���ȍ��+  ��;��Scݺui�e$|�k_�ŋǢE���=���%��                0�}����������Gd�O}�Sq饗Ʋe�FK.��qIIɻO>�����B1         ��mY����,���       FG�������={v|�{ߋ�۷���\.���1�>��x����l6`��=����ҧ?����b         `/����?"���z�����u=��       v��d��|g{����~7��a��x�q��7ǻ���8�裣��2�o2`/u��{��}ϧo�y晻�a,        �����W�{u��n����O���{z       �3{�����������7��M<��3�aÆhmm��hii����]����;����t$���c�ܹC���#���9��5��[^^ްϛ��ҿ�+���D~~���+��)�<����e��|�3�'��}�[N?��=��-        �����~��       �����8���w�����јm۶��IF���uMMM;�\:::b����u�g�#               ����f���:�5��LCCC�r����               �A��L]]]�H`���9�����M(                F�P#3;3��d^+2��������'                ��P3��Ff����C(                &������ECCÀ3ɲ�~/�                �_C������y��LSSS�����                ��P3��Ff���7&+�                `���LCCC�r�τb                �Ia8"3uuui8f ��dYr��                 LyC�̴����I�1��477��I>&c��b         �t2�LTW�d���=�=      ��+))IGmm����ޞ9����         &�ڲ����-1Y-�rI�ۺ.       �:�b                 �9�            �Qr��wF&��e�C/<    �E(            `�|��o�   `��b        ��la�d��f[����~���       @(    ��~s}ln߼��jjj"//oDKkkk���K�6_rB΢E�  �'�|2z{������a�]w��ڢ��x��M�P9�2*�+b�)--`lEEŮ�_�z�       �   �!�޹=��n��v%%%#�ٶm[����|N� ��K~7�PLggg���HK"1]]]{ܮ��0         B1         L:�:�ť7_:b���������<�������m?�;�s���5   ���]�,:f��\����]_   `d�         0�u�ŕ?�r��?�u'���m�m��{�:l���i���   ��U�*.<��]���ȍ��+c"8r��q��svY���qW    #D(       ��������1�tn�`lݾ����C_�eyOoO    �����l�.�?���ƭ��   ��&       ��m���RG c�i{Slض!   ��[4}Q�����<   ��O(                `��                �b                 �9�                �qN(         )/�       0��b         `��
�       F�P         RUIU��K��ö�������w][W[       0��         � ž���w]eq���z��:�      ��E(         aٜe�����nִYö�Y���՛����       `j�aB+������ƥ�E���촾��+�z{�Ϸ�tD.�   ��R1�"�+���]UUUd^���p+//����a����K�  0T,����a����=��l��Y�fEII��{���  "ޱ��]�bފa��a��wyKgK� `�)��Gq~a�yq^6�y�;�ߞ�Ξ����ѝ�	    ��r��Br���ly�.��ŕQ�-�i%Q�-�����c���oYyAq��y_=�������m���������m�Ե-�ƦΆ��ј��   П���(�+��vI�%//oDKQQ��  �555�6W[[[l�>��Y���Fii�OS[ �TW^T�;�}�]�|��t���ֽ�����w���M ��K�c�]\3
+�����Ƿ��ǸO����q��?�}o�v�GK�h�j��Ǹ����dy�������;�?    S�3G5I}^IM,(�s��cVQU�J>W��g�F�队�{���{� ^���ѐ������x�����M�:        `����bNŜݮ/�/���޸Ɜ�j?ӊ��9���w݃�?  �䂧���ba٬�ST�K��ܫ�e�q�{s���z96Ss���q۶�Η/��٘뾩�1^쨏g�6�ǻ    ��P#"y�za��8�|n,(���>/��y٘h��e�x��y��K��϶o�'[_�g�m�g�^����+        ���������?���.>����o��ݝC��EtQ��Ϛ��  �SZP�׼|l{r�{ɌX\>'*
Jc�I�.�̎��f�.��<�Qڶ��q�m[�m/FsW[     �P{-�W�+�o�XK+���O�*SA�Y:mA:v����/�?��l�m���qCl�Te       ��,����Y��Lf��.��$>{�g��?�sT�?�:0.?��ݮ�� ����������ba8m~z�����
��L�IƉ3��a�����yC�m�k��M/���    �P�V�-}9��Da*���$���3yi�=g�92]V����l�G�6�ھ�Om����         Ʒ9s�+o�J�<h����o��h�l�����G.7�p��Y���-Q�-�w}GwGܷ�  ��e������x��I0��5�dz:N�up��־�+M�1-���gc]�󱽷+    ��M݃=����/��T-���+�Mc(\MQE���xS�A�[��������񩸯��4$        �y�>�;�sQUR���~��O�M��)
�wZ��d�ӧ|:�^xt|��O���V���ʋ��c�~,.9ᒨ(���v���-�;o 0��:=���鯏C�Ga���Q^P�O]:I$�����ǹ?��B     �WB�WE�4�Wp~������i��VP��.MGbC�ָ����E��5=ݹ�         F_xy����gO�l�~��_s۞ޞ��M���O�<�^zv�ۼ��o�S^wJ�����O��l~$��EGwGԔ����ih��'�f f���*  ����lX� ����5o��%���)����|q��}:9^�hH�1�X��d�uw    0��b����iql��xӌ���i�#�wct,(���s���mq�K��/_z8lz:zs�SYr@��N��^����MM/���x��xtˣ�ló���      �w�#*3�1�l�n���n��9����@�vY��w�f�7G|�I &��\v�eq�>��>����c��k�x��B1;�^>wy:�F�����  SEI~Q=���ڃbE����s
�h�S\sf��������և㾆u�ѳ=    ���U�)���4��y]W�4�> �3y��J�MN��"-�������Η��4<=�1LA�E�q�Q���[Z��ϟ�y�����G~۶o      `�f�͊�\UL6]}7`l���f��^�;�=�����������~������������؏�'�8q�fz���o��q �I�0/�V����Լ!����U�)�?���HF�Y��T�Y�H����h�   �Q%3���E�f�1�X�(��aƭi%q����h�j�_��H�d��x�����3���禣��9������?�K�^
       `�J1+����N�lP���w�|7������>����}�/*�+b$$�3���� 0%<=|�����㈾�Ey�`|J�1GN}:�b�3��u�?[������c    `d�L!�ύ�f'�X%�E��R�-�3���m[�[�oZ��m��@�KN�$>t����q���       0�$���������b��僺oGwG�͏�&����\.�ӺǶ<��?��C��y�=t]|��O �dS[X<sy�1爘YTL,�El���,u�[�-�-��M    ���I���(��]��9<�/�LJg���]xB�W�.}1�����|��������8f�c��/����       ^VXX%y%1��������()�����������G ��S.�7�y���ȦG�=�~O�����v���9�����_����5��Kw~)>���GOoO  L��8�z�8q��qL�"/�L|5����y��9�קǸ�S�Xt��    �I(f�گlv��{t�y�AQ��&��LAW�4ڶ�M/�:n߲&:z���>t䇢��"��Wo�7    ���l6��l��藗��.����ttww�����{+y.&'�'#�|���y��ӓ>';;;�?�TR9�2fΌɦ��9��UVV3g������#�i��&'�m��ⲓ/R ���9���+�w~1ڻ������q����_W�k�����u[��_����|  �AMQE�=��8e֡Q�-&�L�퐪��h�j��6=?|���    ����d�V,�s�GT�n��3�-(�-~k���'[�Ī�����;����Gkk7���v��Ҩ.�������GIv`W8|���Ƿ>��vY    �gIp���4=�o��=Ib۶m���6a-	�$�����a�3y�':::���5���  ?��ޱ�i fٜe��WOW\}���|&��n�}�x�8��;-N<�������б
I����o�kW_����va `RH.�zƜ#�Y��d�Ζǻ�)�9���ևc��g�m    `��:	d��������J'���҂�8{�Q��ه��b�sw�3m[&���^|g�wu����x��7���]�/9}�a�O���������    v/	qTWW{ f�d�iӦ���$ʑDc`O��󣲲2���FlI|&���Q `��-��U����8˪�V��]붮۫�p�w�#��,��<��اb��*��l~6��Ե�ņ����G����=� `2pTvH�y8q��t<Ҳ!Vm�3�kx<r�\ ;;pցq�[�ث9����sޡ�Ŋy+b�<��    F�P��AΜ}d�=�Ș^8-��v����3������U���� "=��'��$�/>>�s�wbNŜ�n��ɋ9�_�;.    �_iii�I0���"466Fo���ӿ�9�ċF������f�Q__  �ē��z�7�e�]k�_3�s�w�ǽ�ޛ ��,?�����y.�J��N[K</�o�������ߥ�F�e���pɈ�}�ҳ�   LlB1Pq~a�:kE�k�qQ]X�Z����> I}��g���W��S?�C��и���;����n�;v�c��Q����   �Β�hEb^���ӧ�Q�^���$���F}�;�{hjj
  `b�@ �T��[{`��b����=ٯlv|�u���q\�ܝ����    � �L ��8e�!��'���i����?��������3?��[� bS˦8��g�}�����n��C�+   Џ�����f�XL]]]zb$���X>/KKK���#:;;  �vb.���x�� ��K.jyd�����'��������ϊ�s��om���U�Z��    �k�� vbΛ|�U�C��!/N�1_{��xrۋS�Û����������6g-=+.��   ��UVV���c��(Hyyy���$'%TUU��R�� ��I  `x$�$p�Sb��9{kA��Ԓw�3�6Ƿ7�\0    vC(fK`~S����SbfQU�pKޜ��p�����ן�Il�l
������������Olڧr�XP� 64n    ^VRR�A�hkk����`j+--�������0�(yN ����'~��|i�~nu  04o�6?.��X2m^�p[T6+Ƭm�W��5o}>    ��5�G�ү����ŧ�AFR$:a�㘚7�/�����h��0mnٜvĂ#v�Ͳ9��:STP��;,�ZxTP{@,�^�Q\P�^����1��n��u�������;}l��}����{L,��4����&�K��u�����6<�my,�~��x����w���<�?>��c���d撨.�������F][]�w���קG  ��$�/f��/��ʢ��9�ڒh�x��b���  {�{�{�����  ����"Λ|�6{Ed�n0��X_Z~A��nm���?�-.�
    )��q�"[�-8>Μ}D�e�FKa^6Νw\�8cy|c�O�-��
�j�|����,�z���O���Xy��(/��*���<{O\���q�o������[7��5m�.˓��I_=i��N��������MM�>��{̛�9�p��]w��W�c8$A��x����k��}7�l���.���/�/=�)��&_�����s����wZ��NqƁg�ǎ�X��������ۻڅb   �$3��LqI�(/o���2��?{wUy�}���d��6�$a'움���REVAl�V�^�*Z�k-�����V�
EѪXq��\pc�!�=d��I^���Uf�/'3�o>�#�3s�0���<��    T}����֭Z��V   �c��%m�iz���E
h*�{Q�&��Pww�q`�^����*���1'<�8G�������    @`�b,�fӄԡ��a���x��c���~�&�����\����BIV^V��I1I�����֟&�I�:��}2���i��=p��ݲ��/���§�2b-�z��;�+����Z�}O�5A��Wy��)�����F9Ʈ�]�/#��ŏh��i����Km�ژa����lF~�|�N-8���%�K���3����7�����V���'���    �.�Ŧm6��v��^&�*��!+�$�   4;�=��O�����ۛ�V��L   ��a����x�D%h.�����H�m3X���(*��/����     �������'�]T��@c��N�S�h�^������BAvQv��?�pT%���&<f�B��f��ֱ�����u���5��iu��,۱L�Ϙ�wlt���
ŌN]�uN�>��@�(񖘫�ՕH������؇��`��!�hb��L-ٺDM��7��O���6��    ��	��f���!��P��0I   h~���c�ǘ��R����3_=�uY�  ���:ݺ��dH�,�*��^uT�z2�.�      j�5[6��آ4��(MJ=Ka��$z���rB�PO꥿�z_+�o���U�h�����~�	Z<{���z�Ð�C�򶕺l�e�l�g��}FfF�1#���O��~��m�������q�'W<Y�c$E'i@�~Ǿ��ˋ�߸�8-��@���D���ֻ?~W��}{����������m�w	    �6�(KDD���� tY��'Z   XK�3Q���ܶ٢�腕/�x�q  ��laᚘz�fw�(�C�J���\/��D���PEe���      ��PL3�w�h��s;�to�+�͉����w�]�/ X%�$W9^T^T�>��������:�U�c�*|����D#���K4��q����>�[��w�KR���.�z�y?��S[#����
�F@ǈ�x+j���n#���Y�c���xΖ�t��w^����C����K�0ߐ�k��&�=��:Gb�_     ��iX���ń4�=�>_�_c   �4z��֣�Ճ=�w6���ּ�%ۖ��r  �`�9&E��_���X�#<B?��#�ߪ���|[�=Y      B��&���v�H�[�Ҝ��g�;��=j�5���l:�;W9~�s��q#����Fb����v|�׿}]+���a�a+8��h�%�)=9]zOЌA3p?1��}��:�3�y<S��,s��PL�3A��k徕����kt=W�KC���{�n�cddf�z�C���j#1F��>0�����u �U�+Sld��ĵшN#4��xM�;��o �O~\�ٙ�׶���;O_�t���q�?���y��Ϲ��b���Jo�n�#�S��     �x�^EFF�*��	��2+=��k�V)   8]�=RSL5���,���e���ig�N  �
#�qE�9���y��Y+�T�kL�O����ᕚ��c���      3B1Mhd������ڣ�T����&iDro�i�[�.�&F$�*{s�V9~��;��KUV�_��޼Ik�9m���Hۏm7�����{�ޣ��>��ξ)`���,��HC�jFKj*cG��;�:�c���n�P̩�6d(&�$O�������2�/:��Ǎ�ʳ_=�?~�G�>���u
J�Y�i�z����fph�6p�����mzi�K��߽�XKC2"4��i������/�Vnqn��O�N2W�  @��<���j����,��q'Tz<=z����t:ճgO@u�/_��K��*�v��ӧ����L��r������7
@hZ�~}�ŢJKK�����v�����R"R @�j�j�9#����W{�҂��p�B�
   X��K�=��]T�����ɩ�48����Mm/�      ��4�h{�~��"�k3D@�0^Dv�-�s����F���c�h�#ั�uǻ%w���_�1^]��f�cv��.'�N��ެ�W�a#0�π�t��;��Ǐ��223̿�� �c��1W����I]���vy��DQ~"iF��6���!��ғ���}��S3�R���T?�����j����ٮ�j�_#(s��W��4�O
;}%��d�q�5��YjH���ϝi/M3�.5�]���w.   �\MN�4���P'�Vu?��}��p�\�zk�;yc���B�M���b\\� �����yC�[���	S�  v�{�#:�0�����z{��f4fY�2^7  A��r�a�i�ek�E/����L���N���T���**�u5      ���idFa}N�˕�lb�Q���T=�]O�|W�5_ Vu�{��vt����q�����d�]�kT�+��}33q�qzf�3~�.�_������y���>�����?��ic#:��3©�����Q�F������hJ�)rE��w��N����#}T�1#|S���z������٫�^���?O|���ʊ�������4C�-L�oRcX�c�&ϛ��v    �F�v[�����|!4����J   �y����|�0,�{�Չ�����3�m��͚�j�^^�r�ߛ  ��֑.��}���:	6��p]�a�'v�c�-ҡ�      ��PL#1^\��n�fuEaAot���A�mS[��	h�&���i�Uyc��@���K�]p<�x��.�Z�H�)�}��z���m���w܈���_h��sj�O#��/co��������^��w()&I��L����H3H����j~�n������15>��X^I�ƿ0�^��S����tn�s�I�?d�B��~���������]2�"1    �Fg�0l6�|>�����Xeeer8Bh�Z$�P   ��<�s��	���g�9[���������~��|�r�}�ś�k.   @S;7��n�6I�v��`�+����3=��=e]/       X�i�Q���c�zƥ	mN~�?��Z-؛�7�V���R@KqV���ʌW�hG ���j~����P��o{�6������>]1���������:����ψ��׹��w���4�b��6�ۨ�.77cr\J\�i��SǨi(�8F��a�am>�Y5�p�Q�@�Yz��\C�u����Xi����f�i��=��E7���@     4���p�\.�8qBVaC�������xd%�b    �ؗ�OO|���������!ר��S��g�iL�s;QtB�6,�_������S  `]N[�n�6Q�Z�*�푺��ru�ӻ�S��L      @KG(������9=.����d��ǝ~����z�7U�-`e��zέ�ݸ��a�z��n���;�]��\9�ʀ�]�u��5���|�z�5o�<��I�I�k�yk�ӝ��[�=�����?��O��>j���7ڠcǔ����v�9F�ֽr���&P5�����~Ƕ�n��֐r�s��W��Αw�6��{^�|��;޲�e�p��    ����nB1hv��n%�b    k21��>zH�;7��ꌫ�S��#����v���9�F/�y�܌�  �U�s&龞��1���P4&e�zƧ顭�j_�1      -������ѵ��(��ʆ&vדn�C�^՞�#��X�k@� ]��"�l�ϔ�J��6E�E��;��0L�b[��gՐ�����I����M&��X�P��ԣ��V���~hp�`%:�S�S�~F���,۱���#[t(��i��Ai��Is5� �����g�8f� W�+WC{�����b��cC�b^��    Д�P��X-���O(   @-TTVh���v�{w�����c�c���0�g7�G�?�w7�k.Rb,�Q��O����x�w�^����DG��{�`ll��?�|��aI=uG��c��Ҝ�zb���㎷���      -��m�ԯ�/��^�om�n=9�z�y�{���:����w�ڡ�V{�G�=i�j��ȸZ��ެ='��}L���ǵt�R5�o�^_���Ym�?�~C1FT炮�MoU��@��w|l�ט�fgƠ�Z���5��H����:�`L��)cB��.�;fL�id��vߡ����>��ic�:k����k��    �)������*�v����vb)   ��W�-ջ[�5���f�b���I9#�u�_�=ʌ�ۮ�]��z�毚o�g4�M�6i�ܹ��f��������b �1��]��|�h��(* �i��==�����w�9o      hi��S{g�~�k�:D���s�G�闪W\{�e���V�4��m��[cy裇��ZU9��YǌId�r5�EŤ��� NV^V���l�2�;�^�cF���P�=ܮ�>ɣ�W��w}��oDc~�1��mt��#Z�����;���Ј�#�Iy��ܷR�=��X���x�i�wo�݌���k�1cB     4���DY	���d��n��'^    -SNq����y�v�o���O]��衋�>���~����5/���H   �%���zNՠ���}���W����qi�ݶו[^���      @S"S�&�1#Q6� 6��3����(��$��
��x�=����^�_j��cF��1T�����k�1&�Т#N_���TgH�!���?���~���IƎ����1�V�3��XF���2�ݠ�coTc:�{�����-�ܝ����z��>�     ���햕�	=^�WEE�y�9!!A    �S��T���Z��x_xD�����G���W����6k���d��/�1TVV����v�$V�5����=C�#]XWg=1�=�u�v      �R�L]��l��e���j�@M�su���o6����Xٷ�Ս�n�7�����1���op|]�:5�E'�7g�:&v�;޽Uw-ݶ�F�2&��ؽBv�𴱞�{���]�љ@��e;�}�����ӎ�;���~�}m��^�s�>F��1��:U�}�ݦ�t��h��v��$�ر     �ILL4W_4N�B1����X���@(   ^W�|�
J4k�,M�?��,�It&��7�ۖ#[�`��[5������jݺ�fϞ-�1�߿_�/6����, �opB7��s����BQJT����:����V�l      ���%ce��u�	�C�vR�����顭�jc�V�z�j��?�����W��m����	]�e��MC1�ݯ�ؑ�7c0B0Ƥ�@E\�\��~�9u����>F��q�OFf�j#�cf���kuqϋ�?��"���V�����f����l    �ԌՂ���,h�'r���d%�b  ���r��l��6�$>>^ �����}���_�����B����ny�M�;Y3�4�;7"���;������>��C-X�@om|K�
�   j㢔A���D��lPsN�C��JٵD�Z)      ���Ԃ���=�����P7qv�~�g���c��� �9/<�U�W�]�i���vt[���:�u�1crX^I㝠r��D�����Z�kY沀c�d�@�g�Sgw:���=�����eF(�Ƴo�{�@��({�Ft�wlá:VpL���J8ַM_sk�c��K8    �<���,h)**Ryy�"""����xd%�b  ��f�)<<\��.� ��:����&k��l�	0�O7�	4���n�u�Ե��r���{���?�76���y^m  @U�C�h���0R ��XP��]'�}t��ٹT�'?       �"SCI�8=��ju�I�������S�Ι���-P/�|A+�U_�/�)�8O�%�����u`ğhGt�1#�RY�xoU���|��Y��N9�9Jt&�66:}t�۝��3��C���T���._����o���ƛ��/#�����Ֆ��9��OcƉ     �Jbb�v��-�0�5F���*��S��    �e_�>�~���mp�`]?�z]9�J�G��z_����[�ḿ5z�����W�y   �ɘ����KuA�~P�S�))"^�mSe�      ��PLt�n�G��RRd�ߴ���0V.pG���;ߣ��:�ؑ�Wֽ�lǏ�G�/iܓS�ڿ3�Y�}�*|�d�'��不��s�S��^�zd�ic����e;���<�([��V������$��)��������T%Pt����aV��Vx    @sp�ݲB1��j��˚�b    MÈ�ܰ�ݶ�6M�3Q���؞ce��t=#:������ɏ�-�јe��u�  �2�ڝz�����  ���Jt���-U�-      `5�b��-&U��{��#���K=S�Q��w����'���j�UxXx��.R���]��1�������+3p��8�C1���/��r}��3�V]&�   ���ƨC��'^���+<�qG(..n� Bc�_ ��j���U�C���o�á��m={�l�����:tH�-55UNg�!��7����J�HT�9|� 4�]����N���W����[�7ֿan�"-3�0�1}������c��jnۏm׼U����O���H   �$DĘsܻĴ���'��~�������+��P      ��p�t�Ƕ�#}g)�^�d8 uwAr?9�zd�k*��
hIJ��'��G�7�]Q�W%../�����K c����/���e��D���Þ��txS�ǹ�;���+���ˌ�㐴!~��j�*yJk�1/��w�Xy-�8G�a]�:  ��	����D����F�'���� ���B1yyyB����r� 5�=�6����،�]�*�0�σ�����
@3[��F��zF�(+/K�-�܌P���35{�l�ĥ�z_�[u��qs��Ʒ�ݱ�  BKbD�����Nѭ��t�i�?�����8_���      X�� ��:��3�E
@�;��C����.T��L@KQXx��XG����UQY�(ǎ����~���6sb����]����m�U�N��223�\%��]����H��ƞ��|����V��	恎a�*lS���"�E��{i�KZ�{�     @�Y-���>0��+?�:�    U�|x��z�.ݳ���:R���Ҕ�SQ}�  ��֑	z��l�uZ�5y X�w&����6�ס�      ��P�g���7=��! Mg@Bg���L�f��*�
h	{�;ڭ���حb[;��N�4"/ƪe?��L���Z�o��]6:}��}Tp)*/��{�6�0���Ґ�C̱�a'�n��C�CWd���L(    �:r8���Qaa���!//OF����@V���     �	c���w|ln�.�U��L2߳�m�9�   �?�9�5��5j������?������w�-<*      �����s��hN��e�	@����\���M���:#�b��h�V��~Z���Q�m�;����:�ӈ�����h���mT�}T{��e��b�c���Q(�Tl�.���������     Pwn��2���#��6^��
���4    �^nq��^`n=Z���3����wI�"  �N1)���%:b��qz��l3����      ��D(�?���I$�����h�k5g�<��ŕxK�'gO���$i�PLJ\��Ʒ8����:��X�,#�27c��g�ؽRz�v��w�!��1��.z��ct�G>~����w����c>���J����-G�hr��~���r�     @�������
����`��:!!A    �-Z  BK��$��{�#�� ��5���lݱ�E�+:&      ����_g$t�ݽ� XDט6z���������W&��6�03���F9��ϬrܸOu�����Ƕ�{���<B���ˋ�h�?F �&V�[)O�Gq�q߻|x�኎�VQy�Ƥ�	8�-#3Cue;��g�'�    ��3B1VQTT$��+���B�]~~��$11Q    P[	�]1�
�2K�;'  L�#]�ۏH`����s�~��*�      ��}R�����t9�x8 +��^���ڼ�B�UzX՗{�Ԥ>�����5^Q�(�xK���L8f�^���؋�P���0B.�x}C1�
�>���&����#�f���<Fm��ϊ�+���~z�as�iцE     �g�@Fee�<��v?�y���%    �	�}�]G�q���_n.�  pJRd�~���j�  �q�k�W^���\      M-��(=���H����9�z�H�_��B������>V�����\f�!�#1�]�����Fd�>223t�����@����
}��Z燡�S�0�����{���\}{�[Օ��|�纠�~�猜�77�i�L     j��v�J���ń���|Y���PLL�    �*}�����35{�l�ĥ  ��\1����F�7`E�#]����j��)/      ДB:�9&E��3SN[� Xװ�����T����`5k��jω=����w܈�4d(��C���؀�7-����g.7�����O�m�z��4W�ic�֙��
�1����������_E��Q�.��~�.�y��l]"     P;III���#?+�b\.�    ����T�4C��F}���׾�9
�W�ׁ�  �'��G��R��V`]�4��5�s�<�{�      4��Ŵu�5��l�ٝ`}�$��Ͻ�d�;�������3��㣺��e�.�?7����J�I�>p|�~3�R�E�����n�ic��kJ�)~o�lǲZg��M:�9r��h��iꀩoW���c<_��{����r�ǉԊ�+�_b���     h	�N���
�A���˓U$&��/   ��/���_���g꒾�(�Q�}�xK���w�Қ��dےz/�  �)���#}f�[L� X_��=��j��8O��      �BH�b���z���J����c\�!:R���|.�j����1�9l��Fx���;<�71�yşUQY��2b,�B1�p�~y�/ަ6�����~���]�u9�?�����O�[s���;޳uO-�j�&ϛ� �'     ��e�AS�x<����   ��ˬ!�4c�%E'�k_k�1�0/�y�\�  ���wv��qi�r�<�5{O�iz`�+�9     @��P�=̦{zNS�3Y Z����XY�2��`%�h��y�����wrw�;׾����،��Žc��5C�	8~���iF����;�/TS�-Պ�+�t��bÐ����}����g���a׫�����	�'��i/�7o��sV#�c�7��X]���     X��n<xPV`���#��   `���3��O���ғ�뵯E'�h�"��˿�ۃ�
  ���^��I�����]�u�H��Z*      ���T(&,,L�H�D:@�t��8�,_�sw���>�OSL99���Z4k��/������fmE挜���>\���z�.yJ�#�R�+����������ʋj}�e��jw���~UJ�%����ʸ1C�p���a�mh�KӴ���9n|T��x�~y�/սUw�?H�
    \eyyyBp+,,���U�   B�3�i.Bb,R2��hs^K]�*|Z�s����9-޴X�r ��1.�LMN& -ץm�����}�k      �)�B1�;�֨��e���tO�i����u��� �8ZpT��s��~��^g\�qZ{�Z��_��-�+W�WJ/=w�s:��9U^����U/�����_�.�������bω=ڙ�S]�������T�]�����o��6�u���wl�?��C�}�6�X��$:5��$]��r����i�     ���v�*��k�E�d����   ��f,�b��?s�L]u�U�������ݦ���k���:�9"  z�&v�ϻ����Ʈ�XY����*      ���L(梔A��V���X_�=Z�����?���BV�`�sB�ug]�:F��k�6'{-ڰH���ҡ�C��v�v��G�NӰ�կr ZxU�љ�Z�cY�C1�u�s���b2vd��=��#j�j�ξ!�u��v]=�js���wf`f��ڟ�_م�:QtB�p��	�ޢԳuO���s��͜,    @(�R(���@>�O6�MN�GV���(    ������>�J���J歚�o�}#  ��c���=�`~$�N~���rݹq��y�      h!����[�M�����{{]��6Η��'�*n���j�J������!�{��[�c-8���c���223��EV{=O�G�����q�v}��3-F�1��ϛ̉xw������h��ܪ�    ʬ�1ºFH$!!AN����
�á��h   nu��TTV諽_��,\�P�e,� @�Kr����3es@�p�G�^W�o�Qv����      A�q;�tw�����Z(���w�O;_�gv-`�rM{i����y�<�ю�y<S_��mG�5���U�
J[���g.���[���㤭���*��l�25��sޟ�=9{�ǉ���o     ����X3�QVV&+ ܬ���   �p�.�q�b1���9{5�|�_=_{N�  ����~w�+̹� �����^W�W^dAT      4���/����@л����YpH�V�U���4��YZ�o��h�M ;eцE����S���bo>�����W��>��q��s����Z��mVy��Ŝ��/��Ow~��N����r^��S���}      ���MLLԑ#Gdyyyj߾����U�   Z��i�5k�,M0M)q)��W��T�l~G/�yIK�-���C ����e��X"���3���?������      hHA��Y�q���@H���D�.<���C��/�һ[��#?�i��+������u���{[�SSX����PLC\2vdT�����';?QS�rd�������g��y�FtѠ��Vx���aN|k�[*,+     ���v[&���//#d�b  ������N~�[�v�� �|ڄ���3N��w�c�wC��WJ/3sՠ����^���9��|/��5/+�([   ��j�_S���7���zf�A}xd�      �����ѭh\���M����g��-�GAi�������ٙ���9{u�+W���5C���P��=k|���\36�p�B}��CUVV�����]�h�#�x��D[�n��q^��U�F�?�9�E'Ԕ�����h;�|�&����m�����F���|��8���t���o�돶�������    �)++��ÇUPP��"^?�!�ݮ��h%&&*99�ֿ����P�Ux<��=�f��P��
�h��s���D�>��a��IIIQ\\� �%i�����ٷ?|?���u曆m�v�7��`����m5u�Tsk��C��h�X�����_���o  P��1)�-}� ����;

      hA���F�u�$ �%%*A��~���*�t!4.c��ݠ`�+{����~sK�OհÔ�*]:(�� ��a^/�$���_��VmTEeE����w4��z�js���כ�=K�+ʥ!퇨{�����v+љh^��[�����)�0[��3�@���f,�!=��3   ��(..����a�3SQ�<�_�4N�S]�v�g��.]���+�b�������/� �o'N��ڵk�e��Ϩ��W�^�Ϟ֭[   �x�wr�ɚ����+{x����*|Z�s�����M��=a  �b�N��k�"�# t8���M�+�scA�r�      @�](&�����./�!�,w]�v�^;� +;�HomzKhY�̲��    ����i���Z�l���ʄ�1;�6m2���d]t�EJOOj.11QV��x��TTT��r뜌�r�ʌ~�����UVs����\}��W�fD�.��b�j�J   ���h-��@�{�W�=����rd�歚��׼�Þ�  �)#J���)5�:�u M�ud�~�~���
��     �ނ.��n�&�:�4�YGi}�.m�     @�����+���Ç9Y�!?~\.ԙg���c��f�	�s��3�=//ONV� Y)�����ݫ�^{͌���v�ڥg�}V&L���  �����є�S굏��|���m-X�@�2�qR'  ��	m�j��� �.�{��6g�C+      �GP�bF�ꯑ'7 ���9=.����UžR     ����\�����'�U�V)''GӧO'S.��|�|>_s��'���"�a,�p8���V(������[��=�x�^-^���<?�� V�n�VjD��MII� 4���8�k���K+J�=M{_�X��~N�.TaY�   �Ct+����뻌զ���SxD      @]M(�U�K?�:^ `H�r��c�x��     eeeZ�p!��F������_�&M�fDY�����wE��E||�\���d��{(:r��|�M"1�h�����W��,��Z�(��4SN�QH����������6�����ڗ�������;  P_�v��~�"�# �0���1U��{Fe�M�{      �OP��	;�qG��kw
 N�f�����g�7	      حX�Bǎ�ڵkկ_?u��Y����D(Ɛ��O(&Y)�����P�t�R3T��SYYi>����r:y/  �1�zK���w�Қ��d��*! ��sM����* 8�Stk��8Z���@      @]E(fz����Ť| ����Dm����R�,     ��������_M�/� SF(�*�P����W�˥P�w�^�ٳGh|���Z�f��9�  ��l9�EV/�+_����  hh�\�4%m� ����kr3�.w�      ��j���4�� b�N�"�Rݽ��檛      �h���*++��G�z���[�K��J���<B���J�������[�
M'33�P  @�)�����3_=�uY�  �X���wu�\a'? ������~�n\��<�b      �Ѣg����u[�I� ��	]tQ� ���     ���,�锗�����jӦ�Xbb�������J�+}�7~�4�C�	   uSQY���=��sz{��*��  ���))2^ H�#N?=���v,      P-:3��y��* ���۪��.�Ή      �ĉB�2sB1UKJJ�UX)(�����'�p�\
5��iZ���***Rtt�   Psy�yj�P;�  @S���[�! �����c�6w�      ��j���v�$]��<@M�آtc��ȶ�     lrrr���c^������������
�� TRR���2YEbb�B����4-#�C(  �v�|eDb  @�r�G迺M6_���+n;�=�uO��g��=      `m-2v����K�k�w@397���'�җ�[     L��Ѵx̫g���r������w�PL�x<�
��!�өPbĲ��
5�㞖�&      X׬�#��� �TJT�f��@/��P      @M������3�7�� ��~�u�6��Q��X      ����TEEEB�2N�G��n�%B1FTĈZ��k�R�'11Q��XV��q     ��.1mtI۳ �uY�����&�(8(      �:-.����c u�>�=��'��<��]     No<�5c�����SAA�����`�PLBB�B���2      벅����Kd�	 j����Ku˷��[�      P�����8�ڣ uuq�!���:m�     @K����#//ό��lL�����Ux<B1A�PL��gO��q     ����g)=�� ��:Ǥ��^2To�J �+�2\EEE    �������6-*�'���I�- ����03:u������R      -YNN���וrss���$f�P��iۖI����X���R��gO�      `Mqv���p� ��ft�e��+��`U��g    hP��嵾M�	ń�����83�  ��3.M#[�W���     hɘ��|�ǞPLլ�����������D�~�4��������p   Թ��zm�k�����Z�P��LԜQs���6�_5_  �y��4F��h@}�ڣ4��(=��=      ���P�ؔAJ�e�O �'�/����W&     ��*''Gh<��3B1F ������<�<��IHHP(�����c��III   �1�c���VkцE�k�]ڕ�K��as��7���7c1?���  �G��V�2X �PƵ������#      �i��-R�:� 4���x]��-ؗ!     ���ĉB�౯^DD�bcc-i!l\�	�4���\3��A(  ���8��S5��$�훿���A{s�*XEGD��C�;Gީ�	�  ��].�-,\ �P�O~O1��ܵq�       ZD(��(1"V ��.O���Ց�\     �4^�W�/��q�>��v�-�����Cyy����e�CN�S��HV���  �/������~6�gzsÛz����f���833g��Ƨ
  X��^��M ������c���*      ��,�i�tkr�a����Џ;^��߽.     ��&77W���B��d��1B1{�6�j�D��������D�"Y͋�  �j�a�:`������ۖ�ٯ�ՒmK��%�ۦ��v�f�9ی�   밇���N	 �u�/����l���      ��X>3��h�t h,�%�ћY� K      -	���e��o�z����P�x<�� a�PLBB�B?{��?  ��UTVT�;���k���;�W���yA�r���#�u��+�@��Ϯ�m�>�  @��f�� * 4��(����C+      �'K�b:ƴ����
 �1ihF�t���     hI�P	����UAA���Xѻ*������***RLL�в�i^�J�?�  �-�8WC���/}ZC;��i�4�����mˑ-zc�ze�+�~l����Ԙ�1�:`�.�{��"k�Z��8<����j�  @�q��ue�� ������#�TVQ.      �K�bfu�0��'��w���zƵ�6�~     �������PLլ�1�B1-���E��y�������f�	   ԭ޿Zß�ϾQ�}X������[�_x���9�Fn�P�d~�/�|�²B5��p�K�]Gjt�h��>FQ��߾��B�W��]K�ұ�c  MkBۡJv� ����m�譃_	      8Ų��N1)��K �Tfv�{6-     @K������t��Q,))IVaFRSS������*\.�BIee�*A󩨨0��Y)�  М|>=���zc�f,��3�U�-�F��6���u��}��f�7���Fm8�A[�lQ���A�g'w'�O�on������*9&�N�2�6�|��}  M/����v� �ʕ��ӿ��Q��L      �����k;�Q�� h*������6��     @K`DJмx�%�ө����+f\-_^^��"�b*+c"zs3Bq��b   ��h�Qݰ���?���Դ��^��q�s:�cn�x+��}b���?w��߃��xL~I�|�>��(��H{��"�d��M\��o�v�vj��ތĸ���\��N���^-ٺD  ��LJ=K��X@SqE�hB�P�q`�       �%C1=��t����S|��.�/�-+�xʋ�T�(��=�e�U�T�|�^Q^�<|�6�p��",9�����w�m��0{�3��6&���e�Nt;b������fv�;7�     ��UVV*77Wh^�������VVVVs�y<���󘐐�PB���K�.  ��vߡ�^�G3�Cc���k��OF�%=9�ܚӖ#[����o�� ��m���i#���2��DyA��[�]�-�*��.�,?R��ey}���u��+�l��
��>[xxDEX;��v���=,�m����fK��;��G8���1��8���5��9z��*�J      X23��(!ty+}�_t�s�8w��[���[���2����.m��^g=>��#��8��c�N��������f;���������T�ӧ��V�@A���c�i�o��>�Ev�&����V� 	K��"�Yd�d�$��m�~�3��*$�����s������dH8w���;��~�:'�k^6+�>���b���wJt���//&w
     ���PB�\��h��X%�L&��*����K('!�e�{   �mk�V��΋eA���W�eg^&a_X�Ov�D���^{�@  �igI��X�)0ujc���P�/?�k��y1].��(���\�q�˻��h�'����,��ϛJ\�9R�(2�����ϒ���"      ��b��dE��sTkUٓ;��;z�C�콅b��w}a��S!���G��ݨ��ޟ�xከ���3�h~S炸�yr�BC��s�      �c��5M���Tʐ94�T*2::*V���i��X�  ���1�C����7��\����U����\��L!#��t�\��k�  `~��i���凋�3/,��KW�w�sw�Z��W>�
�7�}�����	�n�G~wns�i��_�jt����X-	      ��r��O�8[`�jY�H���=���R��w]��M��o����؍�Jww�����O��cW��2���D@`k�Gȼ�Nٕ      �b��5�r��5
	��P�J:��Z�&V���i��X����a	��8`8 `6�����c��������z���3W�%g\"�:�S�n���l=��i������?�v=  �����$�k؛:��st �+3��p9}��k7>!r���������W�̵矓D�0�����M����fX���mц��      �f�PL�?"�/ؓ:p�=�;�c���C��?�]9��������w߾�e߸��]��_,��Y�5���r���ϖ����     ���$n��Äb��*��d2)hlVZ�NŨ�̧������ `��p�4�7A2
 s��~ijz���[��an/��P�~��/��.���a�Ȓ����l�%[��#o>"m{Hx�ٟl�aT  8��o||�{��[*��޿q�8�w�y�a*w\�ȓc7�*���+;��>1:�C�վ>1��䡾�&ֈ�     ��
�\<�,�<{�Tr���=��d��Wm�(~��!��l�����]�Y�<�����r^��r��Gd���    �51Y�:Ժ�>}��Ȭ�)�˒���4�t:-V���i��YC�T�l6+���  ��˕rr�+�կ�Ү�r���e嬕��¶�S������<��9yrד���'�P.  hg�.���6���ky9�{מу�v��7H�{;p�1���7�����/.�̞�s[j��ӌP���X,Om      8�e���<����}($K���@-uŷ��x@l����G�n�R]/���f���uyl��~�O��T��c�Δ;vo      +b��u�.�M�^��X,�}W$�L�i`j�YE4')
���AE��   L�W�_�_���|�r���'ssen|��k�'a_X"���Ai4K�R�L!#�B�ٟ�/��vׯ��v�+�����  ���8[`�J��5�{�|���W��[�<x��͍���4-�z����s[�aΊj��y6�      ��L(��]+��4���p��#;n}i ���ݛ�� ��ݨj"�}���6/�q���R_o|�Z)�����@H      �FM�5��D"!���f�I�R���%hL�tZ�"�������>f͚% `�Z�& �SM�ow���lޱ�~  ε�y�,��4�ty��BrǏe����?: p�U��:vsޟ�ta�O���&���6�Ė��-�#      p&K�,<.�\<�,Ac;TL�6��]��k�w�g�iaMp�6�8vsڟ]��Ýw�[�D=�јT������O     ���r9���k �3>V	�X)4��S���F��$�b����lW�x��Ć��� �}��{�wO��;�oF(  @�Č��-_-�~:���ʡ?������߷��x`�����M��������<�b�j��O۾+      p&K�bV�IG &hL�JI�~}˛����_�0�R�ܹv�c7']zÇ.Z�<��%��킆��i�����x     �R�n-���Q�+�Rhg��$
��Ų� ���Omm��4�}�֪  `q��ݶDИ�{���v����{w�ѭ������৯�`���+�OusRԆ�[�K���"�EN�      �D��\ԵBИ^J���Fn�ŷ_����p���4vӱ�Ə��{ZO��V�#h(3B��,2G~��-      V��pkI��R.����!wˊ��b)B1�*��*�g��bY�     �xt,�����h���Co~���=�m�;�u��7�nN��u������	w4	����ǶQ��yB      �<��Zo�Gde|���3է���u���K�1]����ޒ������j=�,���Ý+�      KX�:#�������,�H�$�IAcR��L&#V�F�i�X�8      c�\.�P���R����m�葋�w?\�
��]��i�;�i[�����4u��{z~,��      ���Ṗ:O��兑�o�����ݫ�/��\�����{���#W�Vb�u큨�?��9�K�Ɲ$S�	     �09�z��UB1�TJИ��T�U��x<.NC(�Z�٬
	     ��wJt���
ǎl�š7w�U���ms���f�?�>���؂�4M�´`\N�͓Gv
      ���P�K(�7��J����+7���?\+���Vo�9}K凋}���/\"�<��+�8U~���      X����url�HD�^���eS����e�u���I��V�z`-*R���%      �z�:C�*��<;��������4*����n|bG�y�+��󾎥��uy�wQ�
B1      dj(��	�p�@�F�+۟~6���Z��s�����?�7vs��7~�t�rE��Xۇ;W�     ��&��ZX'��r�$����M��bQ����AAc�R(&������H�VX�      cD�a9;�� �p1]�r��+o^��:�q�ܽ��Y�������e7��-�b,Nm�"���J4�      ���P������m��[�~��`J]���Wf����e?����5��SNl�)��=     `�R�$���fhhHpl�D��P���#�bO2��P�#'agM�      c��y��ܦ��8���%�=�ƹw�ѭ�)��;����hY����̄��Զ��������      8�iG�[�!Y�X$��r�"��z�]��s�՛6Ԯ�,:%�����3Z����     f�Z�&�&돏U�*8���!h,�tZ�"����}���     `�v�&��g��غ��s�ݟߜ��ᾳ2cdh��3�NX�      �1-sv�I�uy֔�j��^���>��	w����|�����p��U��K��޶�r��R�U     �,L
�&Q��%8�D�'��Rp�J��
����B!qbX�488(      �Z3Cm���K`M곘������������!�S�������;�����X���m��p��=(      p�B1�-X�`1Uy��/>q�ڇ(������ϺO>򾶓?(����IN�Γ���      �0Yߚ��r=b�FG���
���Xe��b1q"e��z     �z�3�ݪ�ղ<r��_�ƕ���V�z��>^�����;���6m

�✶���      �`�Q��/,�F�	��P1U~��/.�c�ÏL��?_~�����<�]�ه�F} H(     ��P�u�uC(��Z[[�
R�bR�P�i��XS2���ʼ^&f      L������B�$���7�~�_�P��������-���;� w�y�)�b      ĔQ��V�q���[*lz��o�����T�v���vK-w~�i�q�Z���[����r�"      fX�Z7��I?��x<R��{|-�NK�V�L&#V���I�c?22"��nT,�*.     �F7;�.s�:�2Z��xi�-k�Q`���n���F)^�qڍaO�X���
�շ_{�      �gJ(�Һ��GJO��r�7���E�%����}i�)_ر��.�8�UD�a9-6_�~S      �044$�&�ͱ��n�F��?VD/��訔�e��H$"N�J�,���T��P     ��x_��k)TJ������e�"1q��7�n�/�8���;� w9�m�|+��      ����b�f99:G`��Teˁ��������_�ߗ�oqG/�8�����     f��j�L&�4D(f\���U:�4+m��s�I�ضY�     `꼷u��:�Ւ<|��knZ�����|�Cw�nt�?�q�MA�_`�S��=�b      �@{(�춓��r�a���>z��q�#O
,��.������$��v�K�����=R�U     @����T�?&�r���sϭ����p8,�@@<�1��T�V��ǡP(H.��r�|Կ��+�����_L��D"!;v�0�>��y)���3x�QX)����IԾG�U�V��+G�^����|��~H��Q���P�������۷~����      �on�Cf���P�Uec�����5�.���Vo��{�g�E]+����K�j�yM��+;       �7�U�EkP��͇�^qǚ�X�W�|�����X�X�L`�foH�Df�/��     @']����y���577������k	�0Y|Z[[�
�ɤ��3�Q�R)�
��btF�N8���ZZZ���THFG(�H     ��X�X,�������<�-���V��w���s/�\~��V��     p ����+'G�
�W�lx�_o^��:ACغ��"�ٻwitv��tg�O      ��5|��F��7:
�f����$8�x<.V�N�	�4��� ֯N�k����,��]�B1      Sce|���:��3���{�@�����i�m��Ӻd��tg�m˾��c     ��iŜ�+!�}x6�'��������a��^_����B��D@`�3���ݏ     �N�b&GW(F&s�DB� �L
��ȈXA,�a�39�PH�r�~�V����      LN��%�Y��;�����
ʖ�������'������li�%[�      �Kk(��u+x%��?��E"���?/�/xm��=c�!O��&��V��q[     �j2�v��Ũ��̙3G���A60S*�4�t��b�Ѩ8��}��B1����r����D" :}:�i���j��^�g��<gzϔ�>����.7n   #,�.��#0סb��ux�{7wo.�Zg�����oy�#�	L�q���|���      �����1[~��rvߪ;�o�
�mWo��1|�G�����4j"ˊ�	�q��     �����`���:]A�F��z�����P�U�#��E�>*t�$�\N�y=g�[������b�h��Ծ�P �®��k�����. ����ma�������  �8��|�jI6���w]��MAC���6�
]���G�����c&�M#     `o�B1����
�	�S�U噑mWܹf�>AC���^�yG��|2e"�"     t�!�[(&�7��P��$	��)��G0>VY_�hT�DW�L�[(FQ?��P�ZOs��      LΊ�	sm9��wo[��{��v��~�>vk��>�~��L�2��~R�Z�&      �'m����Es���+o��;����w��B��@�/0���q��&`���Γ����7~&����j�v�eChÄ��2�2Y=g�<��3R(&�o�=��%�eB���������'^zBj2��z�=��O&�o>�����"����w��y>�����%�K��)�ܶ�&��W}��/��    8�L&�e��b�P����߯���
��޽����L&�!��I�T+����$:�Wv��(*��1$R     0ys��pV �j^K�;��w��|_��½������ޓZfw
L��ȜP��=       �'m��Ӣ��ّ�K����Ʒ��x t�w���W�s�����!9�y����`�x�.�GZ�.��m��W_^��bub��Ү��l��E-/Z�N�LCՉ��X-���I�:���2��\���Z^�    8]�������v�	��ZB1###�c�Bl#�J	���U,'��1�ɲc(&
iY��� ����qG�n����h��D"�ܾ�.�  �)wZl��<�R��ud����^�Ym����z��?+��R�/� w�,۶�     �/m���"��(U���?^߽Q�醡ͭk7�6m]�����x��K#�	�      -tMW�<�؍��#��d�A��/8�D"a�]�\.'�RI|>���ŘGg�D��FWl�P 34�4I�o~�o�
 s��w���y��  0��8P��'ï�t�U��*��ۯ��r�-�uu��\`��ƶm?�}Z      `OZB1ӂ	I�[�xj�M���x���ި�~hAaZoG �l��2[�/O	     ��tMoi���P(�e9�ZM������Spd���b*@b���#K&�bj;�&�:�ڞ��v�m���3�     ���Z8�Y^K�;���p��������n�����|hf�e�9      ���9)�t�����/��w.�|(~C�?���U��F9�     �C�d���f�#�?��c{��Û�PLcH��b�hT�FW����I\.�؍�PL>��\.�-�     `����"�
��l��w�{%����4m����Pu���eZ0.}y=�1     @/-���j�f��������Q��ݸ恿_�ͮ5K"��Zq     �s���<�k]5�@ P�e�YS�
�������8ҥT*I&�Ѳ,��{t�b��1c�      `��n�g�_�r������k7>1��O�i]z�@�%�ٌq     �)=�����^I��a���,p���{�paˌG�.�@���9D     ��s�����u�\��U�K$��b�ɤ�����F��$j[V�մ,���Y�Hg(F�/B1      �4�w3ӕ}��%p�����g���#r�Lm�;�      �~�4{�2��]�W�V�W��>-p���nzt��/��X|�@���g�#/
     �Q
���������А�����۷����N��g�PL,'���k�,���J�b����      Lܒ�Y�~:���ߺr��#|��͇�����F�'|    `�2���w�}�T�V'|V?�C1� �k��^ٹ��5�H�(;������R���sRt�      I�d}B1�O��jd�D��`� 	��*�Iō�DgxĮ���U���R��     ��&OP�;z�凋�
���R*V�G��3�����Q?�s��     0>�`�T�M�c|(fa��^�ZEve�.8�ݟt���;���ĉ+��	�K��|�(      F`������x��mdd���<�B1�dR`m�bQ
��XA4'ѹ�k�L��ѹ�      �`A�4q���^J�顫��A_hs��:�����/�vƕm�	�ն]      {1<Ci]��w���M[��w��%+����@u}v�]���      #������tM֯V��J�$���
��+�|b��8���e�=����     `�:z��
/���$p���:5>|�`ܾFZмp�      2<3��K�O�V���_8�]_ڸm��/�L,Z&�F}`H(     E��簾&�3]�E�3B1Gg�P��訔�e�z���d��O(�`0(N�+R�r�l����Q��g      �7/L(F��S��ks����Ժ_qK�ӂ�?hC�zOxJv�v���z�]q   0�*��Zt����v�ev|�,�X$'v�(Mc��y\	{��$�	H����C��7�'�������y�UsՎ�Wj���;�����]�v�ԕ���D���#�n�L�?��I^������8������6����At     ` ]�������t��:�?���T<A�7���i�A��S��%�5xw�dR� ����׆��^m<�ؕ�}�Zg*R���.      86�	z%K�ա�N��p���ڑR�S1_��5�� S+UNI*�X{   !�wqc��/k]V�.m]*K�K$�3�e�JE2�L�$e�T�~��h-*��q��|�o�YEc^u�\?�}�T*=��/~�_p���m�BzmO������]�i��o��[�3M�     #���:���A�It��it*����k�}Pp��.�x<.N�"1�C`��	�BږE(     `|\c�9��z1�s�]_�<"p����Ԝ[[��۾��-ԶNm�jR     `>�91~�,I,��m[����V�U��r����@�A'z��j/�\��Ǿ~�T*=�v��A��343/L8A���H���ʯ�<(������E���@���.q��]��2+2������ߜ�A�5�:v�T+R�U�������x���z����7�SV������]B���y��ӟ����k��c���>3��(d׮]������ۂ���^^8�/o2�#�ˬڬ	����&ٳgϤ&��:YN��0��%��'�3��t���k'����/;]���>Y&��J�U#�L̔�`�/�<���ͫ���73���c������������b���   �Jj�����Css�ؙ����O�S��C1�^_���bb��8��ؕ�C1:����|�     0�C		z�=*��(}I�1���k*m՟{8!�j[7=���y�    �[{��ׂ0��0j^����0L6���aԭ��T�Us�[�=�=����^���Δn��hL����&B1:��ڻ�k��ㅃ���_}O"�������s�%�K��"CŴ8էN���w�{�ԛ�N����M�m�������\���7bp��~�2�;w���m۶I$1t����`P�n~��q�ݻ��M(   eddd����C1�	{N���B#kmm5�.X&D�w�N[�+���}�3�h�d)     Ƹ��Zz_��W>�s����M/�r����Zf�B�d^s'�     ���� ��&�	×[.���_UF�N���j�*Keq��z�'?v-��`�]�7����Ѐ��0��t)�*ҟJ�� o�ܽ�|���'�۶�<��ƶyN�؉zd�]�`o�b����!    Ǧs�~SS�ؙ�P�����r	�,��},"���JȇP�q���Q�Ǆ��     �c��ڙ�E�_�3;p�I-��J����=)�
     8~j,،��(�H�׃0*ctF�?+
��QW5�t*�VG�1�����0c��B�kS�?CC13B�	�)�����K�	�+��#�0vs�@�i��������L&#�թ7�R��e��$    s�����,v�3�~_�f��L��B1V	���%�I���b����-���I��-�`�����t�7     �F6�1�ڤK��h8�/����s�m�+-�0g\Ѐm     ���k�b'ԯ�b�~�u�k�xd5�9����9�(���?W��)]N���݅ݲ;��U�a�ˌAk��b�.���[z���o~�k~���Z4:;ܮo��u�5Q      �kҷ��m۶�K��@@�R�ԃ���S���]3���J$�=��xX%D�wR[��D�Qq�����^��/v����b1:��Q��Ծ      G�`��.�e�m��3��q��qk���sn���"q�"��:�    �Qy�^��2KD����zF�No��e�j|�:9��
�Lu�X+����zfW~W�:X4.�B1큨�]z=:]�Z�d9�O�����ͳ���3`�ُ    ��蚬�&�X�R*�Ď�^��A��rZ���ݬY�G���R��̒J�֤֍���фB����ItE������]�=jߪl�|��(��_�b�   ��СC��A
ٲe� FPg3Qg����n�]��X!'|M`�.Ƹ    P��0���zf^d�,��u;?:_='�T��TF�'S���T��+T�S�=�=�[蕾b_=S���aX(��>۳}��\�q� ��@~�ڱB1t��!     0�����'�؝�P�N�!T�������!��+%�:��qZtC�&tśT�����'TG��!F(   p<���|����x[�n �[�.�$���e*�����x�P��l%��&O�%0T��\���    p�X &3�g����̼�zF}���7^M}F�Q��TGaF+����O����0{�{�@�������X��b&�t�	����6m<��?�����rz ���"     `j�j5B1SL�ϩk�5�D"aj(F����4aR�ڬ w�g^:#W�{��Z���      ���`L\B�B���}���R����g��K��{rt���ԉԶ�'wH     ���?"3�g�um�!b~�i���0���d2R.Om�5W�Io����Ga
{���Gơ�tP��H9}� G�{t`[G v��PoX�ހ���D��v     SK�+��C�#q�d�P(�mY:c�L�b̖J��X��ZA4'��
��:N"e    �ŋ˶m��_��a�?� Fs�14.��P����F���0���2�O��$    h�GZC��l����׷��w�C0ӛ����7�>
�z�pF�N�x��Ҡ�/엞BO=���{�aƅb��:��Y����n�$�Q�'8vC(F��@\v��ŉ:��l2�����R���\w�u�3Z������I�l�rܯ��˗;�L�   �/����~�>0�Ig����c���T(�c��ⴈ��ȕS"e:C1D�    (+W��_ ��w}��7p��z���@�q    ��.�w�|��OJ���? ~�u�3�y�*���������멜��A�z���˯s՜ Gc`(�Y�f�ғ�+�1d�;k��_�\.��:1ٙuf(&�
ϱ����)��T��zA�x81,   �b����9Y_�~�����v�Z[[;B(ƚR�bL�3r��:v��l�b��e�     8:5��;P)���M/
pw�y��󿻼��6�o�"�    ��E�E�k3�>�j��x��Q��a���U�����_����/���`}��Dv@-�k�P!�� �p��y�w���qm�x�m�x�8�����d   �[�L=��#>�OJ�����BWW������wA���zŘ�}�1B���P���     @#J������P1N�F���#s�����    ��*�1\�|�����j�:%�PA�����[蕾b��ߺU��jmj�(��b"���x�������Ю��ĉCE�l� �x�P   ���k������%N�~���Q�P��E��z��R��vFFF�c�P�z�:	�c��Yՙm��l��      ��Z|7�a��~F�q,��se��PQ�}     )���qT�"0�+�K�x=s�*����A�C�C2P��aTf�̉���!���#a�sv��X-Ir���a��ya�P��"^�a*�xh�b   �_7<���'M�W���tZ˲t���b14�>�z>`�T8(�͚}7$
9�x�:[���]��^��ia9:�Gj�C(��\��$    {!��G�4�#�!]�o���Cq2T    �ݨ��v8��VA����M�BFb�ظ���ZI��d=�W쫇`TF�y�4$ձ`&CF_F|aG�}�,}������E�![��x��SC�1��9��b   �_�+�>ٹs�̚5K�:�,�+?ذa��r9m�Ե]<75�J�֢�=V8.���N�3n�֯��,Y�D�-[��   �cIDAT&v���'O>���J%m�T�q�̙ FjK�I[�M������\*x�����K�Z�.   �-B(�p�ZU�J��è��`MjDi�6	     �BE`�x+}Q����χC0���B-�0�JRR唌�G޺�����åa�V�?�p4Ƅb�kq(��/�8e���j���D��ř&�^�H�(�b   ���b&��&�?8Y�t�L�>]�R���Ȉ��:�����U�o7oƟ����n����F��$:�V�5���H$l���x<ڣaD�      �,�	�_)���a> ��|�ʍ��βRg0��H    �����=���H���d>)�BF*�ʔ/g��v9X>(��Q���PL��H�G�	0N�y��}��)�V�!�{��� B1   ��0c��݃j�~KK�� ���'���|�d2�D�`�P���M�̈[�b1�33�CD�  @#R���3�+  �Q�.�4y�d��|� p���ƺ�i��3���&w�u     ����s�+��1$%��E�VxM�	.f2��{��6ۿ���� �G(   �L�7��u(��d}���K��h���w����X�UB1vh�&3�Vv����~	�B���-�P  hD.�K|>�̛7OJ���޽��  `ʵxC���X�rn� 0����!c �;�����     ��g���P��J�%& Y=8vc��>&ja�7��8K � �k   0g��SB1{��ն<���
����
��
���I���'l����:�@�
�Ř�����s�D��ۆ�
 s555����eƂr�����#)UJR�  �xE�!����n& S.��Y.0T�&     `��b���x�j�& [����,&��o�U�U�n��~��B�    ��鞬����vgF�AM�'stj��M����� c�p8,>�O�.�K���e2)���l `��<.�tH XDG�C.=�R9�����O|]ny�  8^!o@`�|�� P�^����P!�@      �0$�s�ů(VK��m�%�䫥}Cy\nq�]�5�& 0Y�`�P    �'�B!GL(�D"ڗiF���x��z�hddĴ��J��a���NQ�T$�Lj]�SB<fE�:;;  ��͉ϑ����5�F�}˿׃1�r^   &�'��JR$�	)Vʯ�u�     �cB1n -]�U������Sы�b���g�`��=)	   �"�q����9�d}["�05���b��ᔀ�a����x�SB1fD��   ���]�|�/�W�����M�'   ��0�]�bMv0�jy��p��     �CB1����-�LP�Z�'0�O�b�$���G�b    �+�˒�d�.�)����9uG�
��ܹӴ�R)�5�c������)����V9e�c�s�}  ��r�,�lc,  ��ː������M&�]�����<      � Ӡ��b^�	*��{��{��� `��    "����'<E"q�h4*.�K���d��1;�A(�:��T�U��F}{�$jߣ�Sc3�8f�O   #���ox���_�l1+   ��u��*V˲����`r���ؽg��M��H<�      �aȑ��P��ʵjI�	rWj�t��#|�8�8�<�b    s�"fLb7��땦�&�d2ږy8��582�C1*N�z��D{�~N�fFX�)�3�8D�  ����)��s�lޱY `���yٲe���}���ŋ k#�`�R�ĠOLJ�V���ˇ4��      �aL(�H��V�e&�䩎
��SˌP��������իWp�-Zd��53�-�b    s&�;)���:C1�r�!�D"�#kmm5u��j���hii�K�^��������8�1�B�P(h[��%   ��/���u����(�������޽{��bV�ZE(h �q7^�Z%�I)�*���qBh      �0�f�%�`����$�<�]osDo|*�a��3�8C��e�	��b    &�M�bzzz�.SM؏�9*u<F�1#|X*�"cj=X��Z���=v
��h[��ȈT*�x��  4�]C���{.�Ƿ?.   S���N�U�B(�R���1'C     �C�����0XM8�	�U�%���.�`�91�9�    oEEtsR(ƌ�U�̙#82��/MMM�ɘw��d2)3f���*�'EL�qX���P($�@@�B�{t�b��j����  h|�ZU�����_�l1+   S�%�q׀A����0`�hn��      �aH(�R���r�H�c�j~W��p�jY0u�`v ΢&��n^�   p4�IM�W�����F�H$LŤ�i���觞���c�N
�)f<���	B1  ��l?�].��Ryb�  `�r�1�Fs��&���p�N���     ؆!��R�H��<�2d���<.O��p%bYS��� �
�2::*   ��߇GFF�.�I1Ō8���O�R���{���|�J��
��p8\��:��(��{�
�,X�@   ��Z��uO^'_��-�!  0��y]B1���Ȑ�8*     �}�!�`8��C(��H��p|� ǏP   �,�LJ������3��q��$3>*c&�������1־L3��f2c_k�z  ����;������   �1��x>�L��Ȑ��     `��F8�d���`���.0����Π��T(   p*3�"N"�1Y�P����I��s�c�VXN�.����D"�$D�   ~]�V�o<���%�%N @��U�NV�Z ���w��~�'�?�_߽�(�8}��w��O`,bY      �aH(����y̞Ƅ��;K`8bYS�P�\�b   �d���ڗ� ���P($�\N�2��|}yj�82�C1�dR`���Q)�͏q;m�Ⱦ�xfD��X�   �sp�\zϥ�y�f �>�O�%�\2����}M�z�)И�D���چ�}�� �T��O���6     �>	�p �x;�!���u{fGm}����P   �lhhH�2͘�n�x<�5��u;c����PL:���b0�yR��X��"&f�{��755�CeŢ�)���6  X�zo���ur�}�H��   �8����!�	py\�+���     `j!�`�&O�����	��}�� ��z��R��*R ��!   '־L�M�W����۫u�j��9:��`(��9�R����h=� s�1�=T�����ږW*�$��Jss�   �m��N��=��-;�  �YJU"	:�|�yL�W<s���      �aL(�Ұ�\c�Z"�r�KFO`��� ���*���c	8�   8��А�e:u��nf�Q"��������d2I(�D�b������L~���r����QԾ�P  0���ݳ�����l1+   f*��" ޥL@���9�A�y>      �aH(&]���.�b0���4��Res�tlW�b �"   '���z���ï@�jD�x��PL:���*���B1���ڗs`�L1#R��=�f�   3��!��s�l���&  `i�xj�
0aw`��p��     �CB1�2�t�'01_�3G^k�� ��"8�   8U6��b��u�jҺ���1#R0<<,8���VS��L&����Y~�_�m�SC1D� ��*�*i��Mқ���] �Y���=(7>x���ny������,�]~\��   �$c<�h�(cB�� ��     ؇!�j�z4yK����"̺7X�P֔"8�����+�rY    '1c2w<'R�ݘ�?>f?'���<Vx��11c�d�6�
����3<gH�f�}�>�>B1�qR�/��^ٽ{�,��{j��e�  p��ՒƮ�O`�x��K�	�{�Ck���      �`H(&Y�
��7/`�Nh�?�q�P͒��>�� �
���y   p3&s;-�p�?��G1UG�H$L]~*��'�L�}�]dߣ�2  `g����^6l� �bQ   �J��l83d�KW0���v�]��z�L���b�;     ��2=U�	����;Z%�^ 0ѧ��ق� �   8���#��8���C]����e�c*����.82�C1V�8����qq3�=1"eژ  Σ�S�{ｲ{�n  �:B1�k�]=O����a_�S��9�%0T�1�      �bH(&W)H�Z����)�o�|���u��78�_p��p�2�, �*j�&   �4fL�v�d}%�j�(j����knn��o��S����\δ���Զ�I���8�1>Lm߼^���em��f�R($ L%����7�ˎ?`$D}���eÆR*�x ���*K�!$��B1�����pi�}      �bX�%U�I��E`�fo�Sc7�Cg0�L`8j�SK*�\�b   �D*"�[<�R������4c7�D"!����,[�b�q)&8�g�H��Z*X�N��/ש��]Q����A��U1���.�����&����n���z��e����iӦ��|5/�]   �[�X�Q_��n�F�cHZ> 0\�ȶ     �N�ŔF	�h�7_(�bp����v�-!0\��LB1���  ��Q֝ʌ����cS	�B1*����$�2#X�n�1Q�$��a�^��__f�b��B1  `����۶m���~��� ���w'pr������VU]���{ $��5��uT�GQpA�g��ܙ�;�2	$( ��@e�fS�%l!���tWU�յ��4����T��T�߷?��,Os��9�O��w T�47t�غľF`L�y�Pq"Y      5�b��̓ݚ�8F��1u	&F�S�����"����S ��   x��s}o���@ �hԻ�o�1�j�L��^��i�q^*��U/�lī������+�2�=  �\���G}T�7o  @���:OGLn�|�¹M�/h���YpzlR}kL��M��     @�X(��$gLihm>�y�o��\���c'8b� w�.��b�}�   �kl,��b�^��H$�F���xm�̈́bƎ+8+������بp8,��q�Jq���{  ��*
Z�l��.]�|>/  �j���<���T��JO	؎x��Ű�bKZ�.�X�     PK*�a"�!P�B�����.`;&4�+T\��Wg��B�Za.4�m�b   �56q{}��	�8���{8���@�H���X߄b�T���|�񸼄s��l��� ��a>3>��ڼ�{X ���5��i�4�]��v�
����"Y      ��b�&��3���"��8�y��5�����#6v�X� �G$^8iP   ^`c7�����7w^71�o��I&�V�'cG&c?ĝH$�%�������㟍��   �~��.˖-�ҥK��  ��+q���ч؁�u�	���     P[*�a"�1�������/=
�J\��������.�e��C 0��p8���A   ^`c����n���8�sG6�ut\j&�C�XL�`P�\����b�p�v��{�s��l�c&Pf���
  0�sb{{�:::  Pk�C}���>*kR����/�7�'�?�T�_9��yGN�o�*�?�>�     �vT�j@�	�i�ă����Y��?�W&ֵ|Fp��Y�D(�Q__O(   �a�!Nk&V2,pz�y��O�.l�����s˖-V�O�����K3k"N���Ǆ������cc��Z���  `G
���-[��K�:�y  �i�S��0Z�,3�?�����O�+�#�6�*o� k{      jM�B1=�~��� ��qu��E(��+�6��0Ep�&B1eE(�QW�gI   x��P����c#c�̎�K&��B16�^��f500`���T����\��q�=�1�Ѩ����0ߜ{�  �1����� ���k��{���~���P�̍	�8cZc�)�azØ�Gp3T     ��S�P����K3��	�73:�ж�6�Q��H��R��8�$: ��   x��K��0����D��1mD���͠A&���N��6�	�؈V��H�י�ӡ�=  `{
���-[��K��O @�{��� �m� s%N��86��E����zJ�_|��y'L�om��k�     jNEC1��6�qHK8|���o��^!�/�5�����U����)� B1   �
�X�韅}>�b���.�;>��8C5���f����W}}����bll�1�s��:�6�=  `[�g���vutt  �KV����)f>�5����ӓ��غ�0W��q     �=A��W�����$8grc�E"�����ysf5M#8"W�km�P>�b �b   �6oG�Qy����6��(�LZ߄K�8�����F��ay��s��c�q�  �
-[�LK�.U>�  �׼��5�N: 6�s�=7t�W�<oιsB��&+8�c     pHQmbq�C��M��Կ|%J��/:y��>y��>�\����~�_pƚ�-ñ�� �   x����,�����f���;���%	��g2�C��)n�x�h����;ہP  x��\�裏���C   ^��o���/_���G��������?�;�q�4*�n1�c���,      �n	���V(�Bs�+��8)�jB�ea�驂�������cS�
�y�w�P^�b �b   �]]]���L(f��h�y�	��	�����;�ېJ���q�2{lls�1��>��  �*�ղe˴t�R���  x[>��]W��1�a��D(%3��/�q��t�     ���pPPeU�k�;�J�)j�qpb�Ig_9���o�w��4�?�%Li�I+{	c�� �   x���ijjR0T.�st\�O�8Q�>�1!!%#���!��n���̹g���`�s���  ����裏���C   x���P�sfE'�~���>������Y�.���}�&��5�     �1>B1N
*W����`&�j�&8#j��'~Pz���fŧ|Fpԛ}L��� F(R ஆ   �y6B1,�����tvv::��׼%	k��T*%8�P��z{{500����x��������<�9�r� �[
���-[�%K�?  �;��ݨcZf�0�a��\VzJ(�æԏ���p�J�q     N)*+8&X�2ϛ��b�v@|�g�l;��m�y3y��}��'׏��$: TN$Q__�   �Ze��a� �B(ƽZZZ��oX��/�d2��O�bl����wĄ��Ѩ��s�2e�  �7�s{{��l�" �N:Ip�c�7N �7tށ��3��蔣~t�CO	����wP|��Qo�r�     ��h��TAY*7�=g��K�'�y����sOikk�w~[pTz�O��,)'��
�����	�   ���8B.�s|\��ƶ�i�66�F�b�c��n���K�E�*s��X,&���oNg8�  ��BA˖-Ӓ%K���W������o�r���B���ԍ���t_�sf���8���l�:     ��'RV�&����y�&�>�̅s������3:G?w�Q�5�z��\���nuuu   j���`���^�ZZZ���J�g�X�����F0$�*`��̹g��Վ�ɹ ����٩�����  ��m�R�P��C��si�>��N=���|T��/^}��ǧ�en��~�ya     �����c����� k��(��S,H��I�±��`�G��+x��7έ;�n�E��^I;{!7 x�   �:��
���؈C���*��*ۗH$��m^���AE"��2����jD=�~��.��e��C( ��U(�l�2-Y�d�9   v�ī�Q�N���4#:���i�g�l�xC����rz��y'     pLQ=�c�j�Vedf|�`x=�FG&��ut�>������ߛ���kB�k����IV,X�bj�P^�R���  @�c��}�����3Fؾd2)��gm�(�N���U��T*e�[��q�s�}6��  j�9Ƿ��k˖-  ��y)��P�ŧM������Y$Լ���cS'�{���     '��!8&�6�t��K�+v[NS"&㼦@�ojc�/JOj��/;i�-{}\p�P!��z��E(���  @�3���X����M��Y�G(fǂ�����p��B1ΰ����׎��{쳱=��߯��z ��W(�l�2-Y�d�9   v��"
6�@����ߟ�6������P�J�q���W����     ��M���v�����([sXr�Ͻ�g^���5k�Q��A�`E�e������ x7B1   �u&�4뿗	���yGǵj�F&�c3���d2��O����������XLx��}�|�0a�  @u3����vm��uv   {��(��00�
Κ���0g\���焚5gl��)��q3T     `���{�۳�檁�*5�����
����6�����3������Y��w��i�1K���*��� x7B1   �u6b!�x\x������tww;:��HP5J&�Z���<�g�a;{)c�=6�`M�	�0�bs�q��0�;�  P�:;;u�]w�P(   {Ƅ����~�ɂ�m���[�����,j��W�z�1�f��`�9��c     �c|�N'z;�Y�A��!��Y�Y�I��L�{ڸ��KO?&Ԕ�,8=vĨ����a�K��B���n�b   P�������^
"���&�b�ɄblI�qD*���-x*bb#Pfp�y�`0���F���8:.�  �_GG�  �2z9��P�%�:��Uz:Q�9�'&����V��5�     �y�b�v(�����*B1�2����?�c7~��_	5c�����G���b����@(����~��ae�Y   ���܆x<.������XC���qC��2���o�S�E���s�ys�q:ù     �^H��3''�q@|�o\�����+��P��X��E�ǧ��1�6      Gd��x�z+�+m�
��_ڵ�It�"���5�����ы/hw��ST�W�>��j��P��W3��ʏP���D�   �&�Z�m#��v6�Iww�������}6C1n�ԺB��x(c[�1�q�ihhP0�˜{֮]��6BA jSSC���Tk����](RSS��v&���$  ��e�75T�)���-'��w~z~��7|��'�����'s|�~�	֘c��c     ���b��֌vA���@/�W�??��@D�crCk��񏔞!T��/�7����k��	{�t�& �3̅�,�  @-��X�|�61F���H���R)�!�j`s���i�������э��
����N��H$���)��P{���UWW�Z���^&6Z�￝��F  T�@>�ҫth����@�oN�޿ɴ%Z�-�nbU�����uoc����0�v��     pؐ�	�y+�ӛ�(W��O��::9K����>�_��#�_p��/T��ms����x"���ZҵB��C ��/v  �7�X�m#�Rl,�7L,�P̎���	y���:>v���,�+�1�EL8�����b�L�\N� w�     x��q ��f4��m���X��QB՚\�،Ʊ1�*n�
     ,ȩYkǼu`Q+�@�y����X���tҘ/X�m���#T�&�}|Vt�(��L�_�{�U
� �P   j������(ngk�����	y��&����"T�B1^:.
+ۼ�s�6��.f�ݜ{Z[[     ����¹�>(�utb֑-��\p����s�5�/sS[�:B1     ���jSNp�[���V*P���e����ߑ�f�1p�Ќ�����*��k>z��-�)��Ү* 8�P   j�֭[�����ņC�Nlm��ȄZ֮�s��T*E(���8���[�|��q���~��=s�!`Ouv�_��5]YB�p��|�6l��  P)��:�y�[�#ޙ+t����=�}Wg�х��J��.���F���.s,3�4      ��)8�P��[�REg�ߞt������M�o����B��������w��g����/f��t��$�dp?B1   �E�\N�L��q�	�lS P4u<ZA(fd�����2�enؾ^��tu�Y�ιg�l�{�{ �ÿ���I�jU��-O����   �k���tƸ���QOn=������7]���}���r�b��	�qsg     `EQ+G�������J���5B1.�w��D*ۻt����j_^p�}�Mu��`���,�Z!TF�P �5B1   �Ef���Xj,�̈́��V؊6T��A'/qC(����4[�B1����Р��>G���     �~&�@(��h�����5�i�|��͂k�s��GG�z�%
�`�W      �qػ'�ސ��';_�'&#��aɽg�ˏ����~���W���|౭�?5�Wx�g���=Be�X ���   ��Z�� ®2!�իW;:��� ���,�H2��6v*�*���x<.��!�}f�8���     �͞�~]�����;Lm��_Ⱦ4�p���sѮ��pn�A�I/Onhm\��̱     �q>�)8�ݡG*=/gVk�`J�#޹���k������{��ˋO\��<n�q�f?=�.\㱎 p����Y4IL
   ���"m�o��X��Аzzz�F���qCȤ��޾f��K�E�����l�9��_���1m�      �l�0���^��Q�0;:iT�PX�x���tN����/8=rX��WfE'�\��̱     �qEgZ%x�;��^��n���';_�ߌ?Zp�G������;>)��YW͛v\r�����(�����P9D  l�Y�UWW���~   ���"m�P�,�ǶيE�}�P̎566�\80��u�iB1c�M(ɦ���B�i��8�؈pU��������s     �;̍	Ÿ���)�r��W�l;s��m���u��"<'���A�iW�f�     ���Bb���	��̩A���9e�A�_x�{���$��s����-��L�Ū�y!��:��r� �B1   �5[�nu|L�P��&O�,�X"�І�PL�HL>���=���Kl�b���w��s�yߥR)k�=      �Z��5�����qp���!ߪU����Ӌ�e�ޢ3�m:�)�ʁ��Db\�??�%]+     `�*]���wB1�,��ո�J�瞵�<��������?����w���+�^x��'$|b\]",��c[��-&   ���Y�c����}�%�I+����>�r9�A��2�Qn/M�'�u���͜{v�湇�     ིŜ��zU'�(��~�)c�>ߊ�N���[�;7����<::��}��F�󇭯*[     �/�{��+կok���]�A�Ţ�xQ��x��>Ǎ������s��Z�u�umw�	�9wѼ���r��p�.T(�d��Be�s l�   ���oww��� |���|>���[�r=�H�P�-�t����*��	/mkb���}��c���M�&      ��c[^$�R�c�[��UMN>�Ƌ�^}���f1z����S�K=��z,     `�����(jY��f�P�{�i�kf��s�;��X#T���|�Ni=�@�Op��S+Օ�*�P��!  �Zb��|��q�	��P0Tcc�zz��"32�bj�ٮ�5���D"!l������%      �ߒ���'ׯ�`��>��65����������o������>pBr����%+���\��     ��'
����M(�;1�k�뵾���sa�[���l
�/\�����*��?��sG����/ �W;�u ��P   j�����87��� �N6C-&���d2��Om�A����P$��pt\�=      ۖ+��d�+:m̡�;���C���sOdQ���	s��������3l�F�.�d��*�     `E�P��ŘZOљ��Ţ�ߴT�L=Up�	�-uw���"W,8�����+�6όO~���^{	�֟��-/	�W( �B(   ����l���Fk׮ut�����@ ?��X"��6��&�(�N����WN#R�^�ܳq�FG�$     �}�oz�P�˙pɇ�����>�غ�Ƿ��S�(���6��ė�9!���~�_p��6.     �%�Z�������998����?�)')��U��N{ط��t�+NY|A���ӭQ�.���#�g�fb<��oyA��A��LH ���   �%]]]V�%�s��f�7n��}�hT�`P����z�!hR�R����}>��"&6�=�pX������P     �{��^�U��5�q��^f���Q��iZ;���ܛ�����=v���f�F�m?*z���̱��     X�+/8�+�NkU��'���3[�똖ق�O�'g9�tG|A�g~t�}w
���{�=���[��l$�ý�� `{�   ���X�m���ي�}�P̎�y�D"����Ƕ4�U�L����
yg��ƹ�@����N�lV���|6      ؎�6-�W��.�߾��c&ԍz)�(�ݫο�߄�v�5����~/n�N�U��ұ
     ���+������C�����"�[�>2��;��5�r�z��^ܶ8+���r\sb�/���"T������g�  v�E���   �[WW��c�����v�V���>Q��ɤ�P��I-2��t:m�{�R�dppP}}}���L(fDl�{�      l�C���s����/(�_<��?c�a��zC�+7�v�W���]�kN��wx�}�%�ޟ�'V�l1�G6?/      �~/X���뢞�O�q�XڵB��5:��"�փ>����;q�i_��k��Lء�ms���K�xܨ}?S�0{^e�ݸDp�Y  �SWW���   ��V(;gk��֭[��ki���N�RBy�h����"&�bT̈́bF��9ڜ{&N�(      �_&ׯ�oyEs[��	���g���V7/j������{a��_��;69�_Z�Q�HU���9�#�      �??�[�?��דrp�~��u���t֔���2���~|}��o�x���O���GV	���E��!�闚�%T�laH�t,�A$���  @-��������Xdl-ַq�6�D�ʸoGM�A��.�L&c�[��q�V��H����9�      ��o7.!S��&�����F���՟��>,�����}�&�t�ؔqBU�o�R     X������￢�I/*#skLǮܼ�s���s�����t��Y�f��������;#]_���A_��q��'�v`l*�b�b�oyY=�~��b �	�    ���b�fB1#����0q�����$�I+�y+.�}T>�t��� B1���{fDlE�8�      ���7���S�[��|��Y��M�ѨgVv~��X#蜅�&M�kY|x��G���պ�N=�^)      ���y��^�
�����>��7�%���/i�(���*���:�O�^�3G]��}Ն��-�ʃ�^x�����^H��L�W����^  �   �Z�b}�3���P��f�r9��)P��J�x��B1�c�L�����ʸ�gF���~8T��:��5B1      ;f"�w���.��a�:��e��WM�>��������`�Y��=���aɽ>5p��*��uOq�N     `�OO�l���B�E�9�1�\�{B15`T8<e�!�]�z��k?�����_��#��SO��8f�!��$S��zC+z7�� v�P   j����^
"�)��֯_��f^���[�F���D'������cg2�|��I$�
"e�g�=��i�3	���/}�|>՚���B�p3_�+��k��ͼ? �n��>7�$łB���G|ǌ���t���1��Z7�:=�Rp�U�M��xhb�)���@L(��zp�     `UQO
�l�f��C��N~#�{��ԛ: >U�~�뒑��ܮl�3�k��`��Z�L?�ӿ0�~l���)��>��k�k9?9�P��	�B   �����ֶ2���3���������ةTJ(ۡ�/y)�e�����♑2�"�C1===�f�
���]u^�yj.���k�ktK�p���;���kr��.�L   N,�7�է'�(T?J��z���B���~ܺl���o�p���S����N�T7j������õW{�0sL�g     `�]�?�l;Ӥg���ҳ�N~3w�{�PL�I������1TȽq�O&�}�o�U�7vy[[[U��眅�&��7�i�''7��5���jI�
�Y�b ��   Ԃ��.������F����
���7�Q2����6�5��gSS�g�r����mB<&ȃ��.2�1c�      ����O��U�j�	����#4�9��H�����U�}__������L�\8�i���;�G��t�Dn�Z{�
9�z��     ��^��m�V�����`��g��f�޺\k��hR=wL�5!PƦN,=.ݜ������o�l��ݷXU����5���	u���':q|��/{jٝ�$Zb���   �n�V�/��bñ���P��}�%	+�f2�|l�bl��mH�RV�^m�W���H�     ����#�����j���5�ql���l&����n�����wt4,Xܶ8�*pfۙ��־���'�0+:aV4�@���=��yu�     �*����Q��T|�K_w���.��B�i�G��}���fW�m|�c ��w��ڛ���-�ҢS�jD/I��WӸ�u��P��f3�]���� ؙ`�P   �[6�U__�����qa�lm/�X;g+>ab(ۡ/mE���)"e      �v����1����Q�L`��^������־K���o�v�f����[���J��YW͛��]4:���^M�f�C�1��u��X     `ِ��`��W�f���*��9:i������)'�9�(Ծ1��p�a��s�C�r�>���^L�ޛ
�n��+�op����է�4�m2?n|Cr��H2"xί�?��BN  �	�B   ��Y�m#��b�]�b}wkii�2��I-g�d+8d��cK,F�H�j�E�$Uk��D"%����ۙl�K�^E  �^��:�L�r��G�}&�2'1c���o��os��=���o�y8����o<����������|�%=eL8�ϔ��&��6��<]:�c     �eO�*qQ�e��\�]�%�gG�A��}B_�v��-�@H�4Mh)=N,���b�y��7�y ��=��zfh६�����OO�t��mmm����+�6��c���a����x�ဖpt⸺D�!PG���ҹ>ݽ�i�� T�@     ���Z�O(f����?L��I�����#܍t�l>zzz����ٴ����q�V��s�.!R���5�)���444p;sc�h���;3Pp�gt  �m�ٚG	�x�	�Lk�TzZ�S���3~qXa�`wWg6�F&���`n���г���37�Ӿ[^Ͼqn]�7|D�:<6�5MiN$�MTa<���g��     ��
�w�W}���l(Ƹg�3��c�{���,�i��Kjǿ�׆F�t���!ߛ�/d��������|������B�;P�������Hc0j
Գ���?k�T_nP��P��	�   ������f7ntt�\.�L&�X,&l�	Ř�c���x&�ǅ=�J�l�zm�@lE��Ucc��ܗ98�P     �Ƚ�Y��������x^s��_z������o���bA���Bo~`�??8П��T��|���3O�l��}�|��@��>�k�GB�P���L��t�س�g�      �+�q���b~���M,��k�Wg�!`[B��ᦀy������jc��P�����`� ;c��X   �����q���l3�C1��G�����l#��t:���Lp�6/ELlE�x��3�e�Ygg���ci>�W       v�U���L��}+�~~�_�P�����<�(�3�K޲�     ��J]��v������z��lo9췛��S�Uk��Q θ}�c����FF��?L��Ĉ�������[��/�o�}i�   T�������®����>2u�Taǒɤ�P�������rx��x�ƹ�DG�Ѩ�k̹��PL�P~O��*      v���Mzr�+:nԾ '<���^�u�      ��s����;�;|�E��g9l���mk�E3>" ���ٌ~��YyY����ޏ[�̢۲٬�l�R���ܙ���C7�|��ϟ/`g��'��Y�a5�)��ټy�6��̙3]���,4ړṖz?���m����ڵ<�\   @�lݺ��1���XL�5�B16��jd�+W�t|\B1��d�����4����s�����N9殼&�HX�Ą�      ��-kѱ�f�'�� TV����5�     p�p(.��`���|(�x`�s:s�qWg�H �qۚ�4X��� ��	��!����"����Wye!   j���ڈLx)�PN�b��VL!�J	{��v������1�K۸�l���~2c�     `dV�n֣/jn��Jj�xA+{7	     �������
;_p�^��z��l_9,W�׏/��o ��y�[�mZ*��H��D4n�8=����� �����>��n����#'N�ׄB!   �Ȅ
����X��\���kii�2n&��������]]]V��ܳ{lm7[�	     @5�e�#:~�~
��{�/ ��/t���	     �|���#��lQ�(�pm��M�G����	�J��h���6��'�M��O���[KN   ��� ����H$���b�������ia��ގ��8�T[�&�2     �]���S�lxF� ������     ��b�dd���n/�pm��X����{u�_d�>��{%�F�myI�ϫ� �.�GX   �ml-�nnnv]CC��ᰲ٬�����_�����%����8=��J��=c�Sf��K�=��־I�     `�ܲ�w�@끊� �ԓ��OW�     �%��+ł|�*��������ӡ����j=������ �\L���K��%x �T(   P�X�_}̂�����5�ʄ	��3���F���8:n&���"l���6�-�H�+l@��)�h4�@ �|>���ñ     `י�í���g|H PN?Y��ҹ>     �BQ�
�2�P��ӏK��1�[y��H�T���` ����?jy�: �K08�   ���X���Ȏ�P��W�윉}8�1!:��b��I�R��O�l�{��)'j1�m��rCCC���USS�      �k�����{��6� �����tl     p����Ip����ꧥ��ҳFY�1�ҝ�~�OO:Q �����ɪ��0�l `$�]�  �j����y)�Pn����}�ڴ��h͚5���N�	����lz;��������m�F��c#c���     �]W(�Õ���� �õ�cJ�tl     p���J�\e䡘K����E��9���5����kt�����JǓ�ٌ��b �T(   Pm�Ͻ���V��J�lm;B1#�H$����0��'lo?�G��jf�6�H���g3R6i�$     `����=��U��G �'�����v�     �ku��:�v%���"�bC�����}>% �]�:u��?�B(�Hye1   jKOO�������Q�pX�=��ۊ;T�d2ie�T*%�t:mu|[�klE����+�f(      ��7��!�
���	���s����     �"k�F�
��k3ї��Xϗ�$K~ױL'���(��&FrՊ�5T�	�B(�HqGj   T#[�����X��n�B1�C'�.M(�1��S�DB�}���D�      �����m��秜, �?]ծ����     ��Z���:��,��^̢�ˢE�ߣ���T�N� v�}��ӟ��܇P��
�B   ����ׄb������ӣ��!~��	B1�����R��Vt*�	���>J�     `��b��:�e_�h' �+{7�uO
     �E
2��Ү�b��EC�^�Y�,�<��ͫ�W��. ����x��;�0R���   l����KA�Jhjj�$��9:��'���Vkk��}���Ï��~G�M��#����"&�"e�����)#     ���ł������/��� F�X�ZP:v�ܜ     �ʽ�B�W��U���K��&�~��)?j?��, ���ߣ����F  �   T[��m-6�>�oxvvv:>��g�윉!��&����g�{�R@�ֹ�P̞11#�߯B����900���:     `�-�Y7|��'&# �;��^�d�     �U|�\p�]�>]������|W�_�[W|��>ر����'��,���S6 �D(   PmX�_�l�b�s�dR�ׯwt�L&3<�eBB�5oo;��r\4Q��mh�ܳGL$��b���ی9v�X     `��d��:�e���y'\`�l�֭�'      �Y���.���^.�J}[w��3eћ���x���� �ӛЂ�ܭH(���Z�   �n���2���`�$v.�&32&�|>���^555	�&�JY��}�r\4�s�^�ƕdb;6B1��C(     `��t������N �=f�k�V>+      W)������*۷^\��㧫�5'��f6M l����ά�;�bd�� ��@@   @5P����Bs�[��V\����&xB(f�e2v�i�k� ���Tcc����9[�"e      峴{�~��Y}h���m1�s�      p�7�������W�Y}K�˧�eQ�������U���?$ x�Ƿ��G6?/ @�`�   ���EבHDuuu��bV�e����
���T�t:mu|/ųlŦ�	���2     ��p�����4M�% x��}�~��     p��T�r����*[��P�n(�x{��� ��c0��+~-�_�X ����S P>�   PX�_����q���U(���������T+�����b�������     ��`aH���X�:WA_@ `r�t��#      \�K}�Ap�=�4�ne�R��~�����tT�,@�����w�'�/��Y� �"
�  @�`�~u���|��j�:�X4U8V6�ut�4��ݒ�d������"e^�ƕdk;��o      j��=��U�S�	 ��J�sl      p���"���g��6tq��b��V�R?�^�d8* �v��G�,�R ��p�   TB1�̈́H�� 6b�f��uܹD"�M�69:&���c{�y��Ĺ���ڎ�TJ�\N����
      ��?k�Ԝ�tp�t�Ro��u�     �u+�+����W�]�;t��Xzv�,K���w���%��' ޴<�N?[�P=�Ţ `W�X   դ���ʸ�x\�sf���b����־SmZZZŘ�v��P��
y��o�q�28���َ����ܹ���q v��k1����������M>��7 ��Q,}}��;u�!�+l o�����w      \���u��x�J�c�����W�t�\`i�
ݱ�I}j�q�=f��^��rE�����G(��
�B   ��֭[�����,���K؈.��w����G&�v����ݼ11��|���Wb<�f~755YyϘH� #��'����㾉Dn�D<��k�0(  �j�9��^���m֧�!*�A����w�c��      Wڢ�U����G�ҳ��7����5�՜��;�����ІbeՆP�]�Ż$  �:�r9ka��`k[���عd2����tzxN���G�m����+�E���8瞲1�7�!��     T�S���kӧ'�( ��5��魯
     ����T���(V��b���r�B��K��?����4����^q���٭� �}�`9?�   �cB��f�9��ֶd���$	��4���>566
#�JٽCf4��|���T}}���P&��f���%R��&M����ڭ��hI������<E�8����   x�ͫ�^M�uxbo���_�OW�     ��6*�EBU)��W�A]��J�N��s}��MW�%��!�m��nJ�N6�$�:�B|�  @u����|fnhh��f(�̛�|>a��ɤ�q3���]�N���o�^a+2E���lD����N��555iΜ9������?J�F��N:d�>��	   ��ͭy_}놨����p���n]����!     ��O��6�	U�ܷN�V��L���޳A?|�^]��G�vm�������� �*   �6�)[��l6���>b$;a^�`0�\.�踩TJcǎFƄul�ݰ�V��PLy�ڞ�� ���ת!D���V����e�e�����5�B^   ��'ׯ�x�6]yЗᆨ@��s����J��
     ���ԵB�)o(�
-�ź����r��n\��M����w�' �-��,�c ��,    ���k�������1E2����NG�M������^��O6؊�yi;!�Y�|v1qw�s v��`���z��i  ���ѻQ�_���a�O	@m�z��z�g�      \˧o�*
U��+ls�N���7�gv�^܆E��F�Z�ol� �s���ݥ���f^K ��w�  @u`�~m�F���m�a���&Mv�����PL&�F�v(�K-"e��V�,���l�j      �䑎e�'6Qw� Ԗ���Al��      \�a]����T�P�|m�ź���?��bNm/�LW�eM�k��pӪ��hǋB�+
�]��c,   P	�B1,�/�@ 0�����U�d2����TJ9���Vt�i����ss�=�e���H�      g���{��똖�P��Z��W�/      ˩�o
U�2+l��\�]z��\"��ӿ�x����/+j��v����� �Mf�&   �vfa��0����lS��X;g#bc�f�L���^9.ڌK5s�)+Jnhh��8��GS�L      *�X������e��Y�IP�^�Y����*��&     p���J� T�ʄbڔ���?�gw�E6l��{�v]����W�?@�-�Z�+~-�wCP�B��    �3��\.ge�x<.��	��^���qmF�I2�t|LB1#g� m�b|>�b�����1�sO�����P���ޝ��Q�����t�}�!	9!܇ x���/tWD��*�?wQ�x�G�@ �,����E.E��k�oP��}O��L�Ꞟ����WOc4H��1]OU��W�t�g议ꩩ�SD�      ܕ)du������U��d��;���ܠt>#      P�~ �Z�j)�u�.�έ��!K7h�������*��_6o�OV�Ny*��P��a��   x��I�L��"�bv�o3��|>om�����K���F����Ɨ	�l޼��q��      �o ;��,�^��5Vs��ܨ�����k     �ӊ�H?Q��k�=+6�s�+έy�c��hJ]�>3�T���LR�]z��ri�r��7��    ��5�ڼ_6Q�/3Y��UMM��s��1qx7�5e�Y�R)��!�HX����[��X,&�?[�.�      ;:Fzt��蒣>�HU0��@%������j�p�      <�5�����O�^�u���\󛍏*m�'�U �/�K��%�i��	  o�D"   �n``�ʸ---�`Ɨ��Y�&M�$�	$�u?��:��� ��ݐL&������}Ɵ�ǕP     �=/'�k����7=SU�*�B���+o��5     𸌳|^sT|����Z����s�y����T[�D�}k �3��E�\Ge�B�y�g ����+�   ��lM�nmmƟ��Y�Ō����J(f�ĉ®��ɦ EL��T[�k:�V*�"�     `�#=/+
��C�Y!qq ���9�?[�G=��      |�ǚ��BE(��[��l}NE=�܋�Ć�+W�AuUQ�<��L!��/�Q+�6��P��a�   x����A
"��<��P�ʱ���al&�v�ZW�L$��l�b�1�d2�2v+��������1S�L      �닪��˳�/ ���������     �,WF�	���c���wn}KS(4o�m�G�����;rż~��f��X/T.B1 �FUUUi)
   �*�[����Q]]����>6���cB1nK&���l?NA�.�����D����k�=�b      �s˳j���gf�* �r�t��'     �U��R�B�p'c�g��s�Py��Q�h�o��#�֛c��}&�tي����+��F(��2�4͕�   /V:��26����Lط�1���F(fppP["��:~�B1��)+�h4���:�R)��&R     �����j�}l�?�7ܶ�)�v�c     ���~���x[a��,TJ�l�����ǘX̏�߬�)�<C �1���+o��K��G(�ފD"�b   �Y6'W�b1�<LaӦM��K(f��X�mP��fP'
���YA`s�C(�|�ck#þ     �;�{��G���o ����^w�      |!�ejҷ���^(Ƙ�E�@?pn�P��gt�+��{G~\'�, �3Ѧ�V��HL������    ��9����E([!#����4����R���M�dR��PLSS�����u�-��=�񭯯���{�l����6�C      x��Zs���i�=�d��MO�W�     �O���Oh�F������M�DI���)��BV�_r�.<��:��pO���OVܢ���	 ��e�   ����j�0Q����	���q���;�D����j��D|�k�TJ�\����O6�������P��=6�w      ر�:R����f�[ ���M��W��      _�H�P�ܟ];G}C�V^/9���A�b^?^~��?�u���
@����`�o�||�,n^�@e1    ��5����Y�pX(��	�N��y���d2��i���
;f;�����=A���`��5�Ry"�     �-&V��g���G�p�9�������O	     �G�W�
�Ι}�k�.��[�ȣ�ł���R4���@�������t�CB1 ��_  �eL֯L6߁�al&
�~�zW�41B1;788hu���A�P��X��)/[��9vo�=&L      ��[�U��׹����� �Rt����;uO�"     �Ȁ���� T,{�����k��sV�Oˣ
ł~��e
Y�1��0��a]��:��"� {��  ��lE=��_^6���C~cB1nK$�v��tl��N���K������o7��o      �tw�s-du�!���P� �/s��y+o��=�     �3��m*��ٵ_v���hy�	�皻�9կ/����8ڒ�w�\�M�^�>S�OT% ~�D����T�*���q�    �*��jxx���6C&A�FU__����Ƕ򛶶6�ǴB���A��e�h3&��-D�      �3n}I�̰.:�c������g���ӟV
     �g�;n*��P�<����
��s�ӗ����i�e����T4d������F�Yz��Y;���zy���7���e��=�wL� �V8ޫﶆ۔�f   ��L���3ok���V���0Y���$ėw�v(&(�E�1�V�=eUWW���Z��i��H     ��-���/�R?8�P�p6PN}�������"      _)�I��B �/���*��O)�;�{U��{��wtPs�<[-��;O�.��+oU����P( �Vu����   ���z0Y��ZZZ������f��	�B!a����]�v��l�t��żf���'(��M�1��!R     �놻����.�bf5N����y-}o��:�E     ��lQAg�j1y? �1�v���������<nYr����5��Q�Ҕ:�O8��-��5�8/w;W� T�H$"   ��L��&뗟�O.�S2�Tss��s555�����Ȉkc��;g��ijjR8V�
z���<�(/�����v}\��i      �g�2I�~��ׅ�}Ton;T ����5����j$7*      �1q����"�7B1F��hH'����㶤�u�K��{G~\G7�����|����?	��\ �Vu�w��   ۳5Y?
�q��P�a�-B1ckkks5�HpU�]����b1��}��������=�����     �C*�ќe7�˳ޯ�Oz� ����ו���\1/      ����	!P�3�v�
:O�R�LEb�<n07�o��k��A��{&�  ;7�ѥ+n)�ց���/�rEp   �����]`3300��3g
�fB1�6mrm���Aa���2�����2�YM�Æe�������ؓ�}      �L�X(/�m)c�C�c�y��zÃ�ݦ�     �S����Jo�X�~]�8��t�6y\���OWߡW���Yg(Z��Z=�E?\�u�휤o#`_D"��  �7���L�v��(���ߘP����P�Ѩ�Z�d����XLA044�l6kel�=�)�y     🻻�ӆ�]t�G�m����$���7k�`�      |�1e��@�V(Ƙ�����I��ܫ�<����u�G|\k9Q����/��w*S�s�: ��UW{�,   P(488hel&q��fx�V��o���u��~�	�ek{�MP��6#R6�YAbs]���Ӂ(      �ϒ�:�ūt��ӑ���U����S�n�     `,WD���ɛ�k��q���(��8�B���[t�KW�ۇ��7��d�BN?_s���^$`W�Ţ `o��a   ^�Ǖ�筌�d}w��Ԩ��V�t���m� ��ḞP̎��e�h3"�J��6�e"e      �֗I��/�J��q�>:�$Aww�s���sE;��     �*�]*N�
0o�b��Y��P����`vD�Yr��eƻu�
��q���t\?Z�[��0B1 �E$   �5L��Xwuu�>.��wO[[��c��x���%(�E��V�=�hhhP4U&�q}l"e      ��/�����#գsg���*λB��]��=��      |,��>��Z-�wC1��P� �֗��@�/�ߧE�՚}��m��.����P.%  ʭ���oe  L6'S����0���PL*�*-uuu�Ι�BMM�FGG]3�H��L&��mb�A�.�	�>����>.�2     ���@��Z1�I�<�,�0Y@P�Ln�e+�ͩ>     �X�Y>�yzZ<�ϮM�+j���{�#/����/�\��!���p�l$7Z
$�����=Q( {����4�X,
   �
���c����a3a�P�����͘����z6:MMM
��
[!s\�<�p��P���6      S��ꋿ�ǧ�K��~�B��R�s��zV׬�O�b^      ��W5O�	�B1W+��t��t�s�d�H";�9�n�i�ӿ�Ն�*͊�Ra�3ŉ��s� ���je�Y   ^as2��@w��p�®�����I&����贵�)(l�{���[��L&���a544      �!_,膎����z}��3�_�Y@��M�����z     �^Hj�~&�/��1*������׹�N���/j��&}밳4�q��J`~It��'u݆�(�c����"��   x��x�PWW�h�P�[l�b������b1WǳD�2��KP�Y�tZ�T���n�΂�v��P     @�y)�N_\�3�{�:y�1*��Ku��;���9~     0�j�~"`;���4�o���!�t�|fc�W_[|�>1�d}d�;T�
���[�p�Z��(  l�����Y   T>D���Vƶ9y<�l(lň����������Z&�j+`be����om�V�=���x��l�ԩ     @�Χu�[�h`��������N�_fGt�ڻ�P�b     T���|�/���kf�eJ�\�GQ=��;R>�-�t��H��:���&N����yݶ�)]��pi}���< �*&�   �R&��26���e{�>��v(�QL%���:~P��6�Q6�YAD�      �t����U:��������7��.����Q��      *įդ���b�+գ��ңνY������K�轓N(L�Gx����t���0� L�  ��0Y?8����F������{��&����.��P�;lƣZ����H      �-��ܕ��.�z�3�������?�ޥ���	     ��ܬ}^�� `��1j���w:���ν��CE���]�����{�:��`^4Z��ƎG���O�Pd_ ��j��  @eb�~��8OO��Q�d2�\.��Cchjj*=F�r���2�M��bʮ�}��]߮mC(      X�ܿR���C��~�>2��
U	�3㞮E�f�}J�G     P1��I���nQ^�N��L���l����9���Ou�t�+�鴉��s3ޭ�h� �x�w�~���f�^���X,
 �U8   ���f����cn#c���um	�΅B!�b1W�#�a�I$��6�ss��������^�Ǽ�����m�g      ��\h�W��׳}+��?�Y�x�ʡ���5wiEr�      *JH�P���9*���b�yڪ���u�s����_��KK���N;Iѐ���ۚ�.]��n��X/�\� �HD   �W���[�P��l>�bvO[[����x<.���p���%.kk߳-Zw�
�)��(�
      ��$١�t��c����X�Q�-���n�xX�v?�B��R     ����<}���l���5��*��z������;M>��gJ.��~^��q�N��Xn̍覎Gu�g9x��#`<TW���,   *��P���g�1�����	Ÿ�fŋ����c��� ��Y[�8.c��H�ĉ     ��):��(�Ǧ��H��\1�����_oxP#�Q     T��.�}K�n��#��4���A�u��"x�|�g4��+o-c�x�{5�a��r�v����i8��B1 �CP�   ��F�����e{�>��v(fppP��ᜠĳ���6��Af�q7�s�      ۶��>���eƻu�~G	(�g�W誵wkK�ߏ    ��d:ͳ����������!��y1|Q`qb��}�*�{����'k�N���2{�G{_�����t� 7�0�r5   �bttT�T���Lַ��d}�-��:���J$���v�涠�}�D�      ���~�x��zc�,}fƩ:�i���t�C�nx�4�     �BeT��@7�C�5�v�r��/�-�I�H!�\�X�}�����/�'�Q��v��k���k�����5C[���PL6���͛����:Ngg�.\��}�s���1Ƈy�<��#��{���}��cmذAӧOWs�w�{D"   ^�d��!�}mmm��G(�o̱���k�e�h3��1M;l>��{      ��̹�f1���q�m�"`_���M��K     P�҇5_�����f�����t^�9�jUrż��zN���B)��駨-�$`O�_�����2�Y ^���W�6m*{$�0���zH��u�9��SN012��+V�2���V�ZU�Xg�1�pX^S]]�og  �?�b������3I.�s}�D"Q:�
���^V�a~�u�X�a�(f}�gU)�LZEe�Ⱦ'x��     ����|a�?jV�d{j��V����[�ًQ     ��u������	�K�{��ݢ�Y!����Ob[0桞�:c�[��)�PK�A�X�W��kyr� /��/q:;;�e���5�f,X��K��_�"��S˗/��C+W'7�@���4k�,����K��  @0X���Ep����Ǿ�����M���b5�ZUUU�9r+n`�w�c=�XLAg�O�������������� ��l�o      ������?�w�>9�M���S�QF��ꆍb     @`�I9}PW�[�>��������PXw9�TI�3�e�����k���蔓4�~����?�_��l|T˓�x�W~�c�����[���ޫ��}�;�QSS���=��S�7o��٬��!��hŊ:��=5(�   ��?W�2Y�����f�>������\}}�@J�PL)�c��8�������ǎm�w<w}l�}3���      �s��/��Wt\�A��ަ��&��-Iv���O�ɾe*     �xE����I�ш�}T١�Z���&U�&���0�BNt���_�[�Շx���:K�T>�����n�������0�;�������f�ҥ�袋t�%����Q��j�*-X��j$f�B���kזb1^��V]]�og  �&�a����؛���3�	Ÿ�f �K��������9�j����v�}��P�96h�9���      �'�y!����0Y�<�D�<��CUBp��"��iyr�      ��\ͺPsD1�"3k� ޫ����"�Ĺ]qG����������5��][���;��P.% ���۫��.yɺu�t���?�����`���)�����
3	ɬ�f�Uss��oG\�   ^���gmlB1��|�mƉ����p����%`bb<�\����e4창�!     �=�zx�殼U�u<��Oz��?��j�
�a.��p�bݺ�ImN���*     ��
�Ӛ�;��`�b^U�<]���y1]�ܯ���L?}��u����^c"7��D��ֽ݋�L�
�y~`b6e�YmڴI^�|�r]y���7�!���s+W�y��]�VGq�jjj�~/�HD   �mf���(Buu����;l4������b1WǳH�����s[ln��{��P�Y�f͚%      `ot��������M���L8V�t�j�$T�5C[tO�"=�u���i     �K*��Z���Y�B1�Z�?��z��͹w�*�9�~]�C���a�z��7�Mz{������$���uw�s�Js�`�K�P��-h�ƍ��Vz���u�����O���'��s�='�2��9���
��}�p�4���   ��m�'mii���<�l��잶�6W��>6#n��{��<�^e����\�      P9�riݹ���rH�:m�q:u±j���o$7�Gz_փ[_Ғ�     �դ��(���b��Z�/���/�٪pE���5��=ڤ�x|i�\��&_,�O+uϖ��\|�
E����̕��pB��W_�c�9Fp�,�\N��կ�u###���Ԕ)S�~����f�   l��`��]6�&���q30�H$���7���477����)     �x[5�YZ�]���5��g�	:�i��?K;to�"=ֻD�|F      �RQh��K@3c�\C��O�|ݮ�~��D5�/��o6>ZZf4쯓ڏҩ�G4��L�gir��Y�G{_�@fH��ٺ��6����L&�k��V^x�,O?���n�*?0��	&(�Z��   �6��B1v555)+�ϻ>���h)�Y__/����<On�KL�8�̱��!{Ǳ��]d�\D�      P�R����ZTZ��iՉ�G�	G騦�wu����W�p�bmN�	      ��(��5_��YpC1�,�-�@RQ�;/�� ����:�!�贉���G�=�$���8L����Ae��1��l^�xO�`�ҥKu�G
�q�w�/�빳�S3gδ�=�I   �M�����f��]�PH����&Λu�P�����];d)&dBAeb9�B����X0��6�=Ay����w����qv�ޙq��      @�l���ΧKˤژ��vx�<��&�m�Øs�7�z      ����Q����p�j��ڠ�t�fh��2���f�Pgi�j�=:�e�Nl?\o��)u�;2��'��O�+�d�R�e��,*��P̶��䦛nҏ~�#!Lte�����<y�jjj��O(   �ي�---�]&�ck0�N�:U�5�X�n�+c��N&�䈓�H��W45#�Ͼ'�L�ʬ�6^k�lV���jll      �����_�13���;�;Jo��C��($��n(Z1�YX�'z��B1      ���
�s�����Y��ܢ���2��c*�z��,P���8���\�{J��[g��rB�����3�RmI�������j��P^�DB~�x�buuuiҤIB�[�h���L�����P   l3�m	r��+l>6�=?ikksu<B1�B1&`b"�.�J)�N[�P�}fc�f�=�b      `����Z߱U7t<���z�z`������h0"�nId�K@5�?ݷ\�!     �u���>�+EY�cV�ߛ��u��QH�w���W*���]0����+-��j�<C'��1-35�a�¡*a�ų�Z:ء��k�h`U)��Jؐ��522"�1��C=���>[�|�?�������32W�v�   �d~f�����o%c��`�� �w�ۡ*�6m���f�9(���>kc��Ԩ��N�+�������&3}�t      6�F�x��r��t��;Doh�����6v_*����F��X���Wi�H��s}     |�\��ۚ��X¬�Y����[��~��~��>AP��+N�b�TEtp�:�yzi9�Y��99x{&c�0K7hI�C#=4d/344�����O>I(& �-[&?�d2�SCC��c�  �M�����rV���jj�ꈶٌ�،E��ۡ�]�d2iml���(e����lml"e      ��gersi�ɹ_�Ҵ��tT�9�}��v�����^&�UC�ZR:ϽC+���+�     �1�t�F�o�R=,bV��Ջ���)�X�;��3�=l��}5��,����l�_G4O׬�I�퉚Y��µ�t�]���ֺ�n�Jn���FfG�;���j�ƍ��Mcc�P���x����Wf��1�c   [��x[L$&
	v���X������P��P���%bbs��J(�l>6�? �M5Mj��w~�{�յj�oS��e   `G
ł6o--ww=W�ڤ�X風��K�D�"��٬/����9�]Z3�U
�l�      {d��|I�t�  3�92��B��U�j�.a�L,�Jq�����Kᘃ&iz݄����pT~S,՟��T�֏lպ��Rf�s;����)
V�M�R�+��Y�b�N8��r� ��ي�D"   ��u�b1�>�σ	vf2E��;��&�����[?�&	��PNP"&6�=6�X���"e �����Շ�������>���^����   `�����!��ׯ�DJ�X�8�H�\צ��:�����t���w��0k��4��§      ���&�TH��<ٙ@	� ��ݵ@+��'k��PQW8�vKw:^Z��_񚯷F4�6�I���X�|�i-��߹�\]��H���t��ȣ�l� y&���x��{�}���Z���}c�'6��S~�f�B1n�֭�;�P���--   ���w�n&�{CSS�B����f��ĉ�]kkks-388� ��	J(��'(����|`s�      �S";��kJ��µ��N�i-]uR]�纛���R
������s������o��ʏ
      ��a��5��bì�=5O�yz@a}EE]�|�I�+��piY�ܴӿ�\]��H]�sK�ܮ/���T[QuU��i��-��HUu��E��P.]��90n0�H~T�bQ�|��I�K�KK.��_���5q*��w�)���Vhe��z������   ؞�t��d}o0?��X��8���cB17nte� �b�q���!k�e�hs�C����`+Rf�a��i���
      �D����w����ה�mo�4�.����hU�_���{U��ҹ��a�g�*8��_�.�����|�s2��y�۟�n�}     �k֨�ok�n�Q�b��B�����<ݠ*�Ĺ�Ig		�n�t�{D��' �W�BA~�L&����PL>�/MN1�T�T]�[Z   ����oml&�{G,�����	Ÿ��1ǡ���4�؆���y����U�٬�����>s<�����1c5�4i�      ��J�GKKW�^�      �nX!�S�.��x�j��Bmv>~Z��ҋ^z�  c�q�S�P�nttT~gb1n�["��    [�����*x�y.6l�`el�렟��1ǾL�#ђ��H$��m� �y�k���U�H�w����1c)#            �B�+�]�*}Ws�%�Ō�z��x�f�4u�s�� ��I~�(RSS#T�Jx�C���c��   �I�RJ����	�x��p������b1W�d(�f�8(�D�q(s���^���oڴ����{             T��B����-�J>¬��4O8(c
���0/ �g��a�Y'Mcc���Dbl�����  ����Yۼ���D�������vW�3�� J$��J(�f��<�6"��1�=             �W��r���;������rx5�&���ď��o ��X,Z��1���&���=c�*mC$   `��I��g�0�Dϰ9Y?�+�ϳ>�������R)W�j(&�LZ�PL��b1�;ZZZ��ms=            �}����M���|�PL�5O�ݥ!�߹�-�k'
 �f(�����d�}5y�d��M�6M~VSSce\[�   ��$i����z6��B�P��p�y�ŔW"��6vPB16#e��͂w�\�m��             ���
�v�5O�'�Y��6G��J�:���Ug9�Y��+�@2��l�����v�aBe�9s�"���٬�����ʸ�0o�   `��I�A	"��	ńB!k�\-"3���6uvv�}�.� �3�<��������v�f���}���|>L*��p            �eI�ߊh�.S��
��{n��E��O��Xy}Ź����j �HCC���|�S�N*��Xab1�V��ي1����L   ����DA���\b��d���f]�5k��kn�n��|��ӣ�!S^f�2�[Z	�x���ٲm]loo             xL�B���u�.��+�eD(Ɔ�Z�|���ՏT�Ϫ�/8� �͐C]]�jjj4::*�y�ޠ��*���-o�e(ƄZ������KW1   �40`����͂��	��B16�E?ikksm�L&���Z���q�q� l��81�U4-��GFF��o"e�b             xD�YRHרQ�k�2*���������r�Np>������� T(���\9���K~s�i�	�p�I'��o�ߘ	�����Z�  �۲٬������d}�1�ɦM���m&�cln�bL�!���T*ee\�	Bd�v�����}��P             X֥�~����\��b�b�9����m��)��9�r�  ��L�[(Ɯ�����0e�r�!Z�j����Ճ#��FGG   ��LַC%�=6����p3c+�b����M:l�9L����I�����26�             ���^g����G�W�G���2g�^QZ��Q
�,�q����
`s�QWWW:y>�H�/�������]v��y智��K�555֯(�k   n�9Y?
Y�׳�����s1�v���Q�hT�L��c5f��c�#A�g����m��I��>   {+����gv�5���������~�5����g����Ƈ9�k_��&�;mڴ�ޯ��Rmm���^CC��f�����g.hd�5       \SPQO+�[T��5W]��^�PK��f��]4���� >e;cL�4�7�3�C��,'�x�f̘�6�8� ���   �m6'G��חNB��؜���fK�L;g~v5�Swww��"㮠ĳ�e2Ծ
J��ol��6�G   �Oے6E�_T�ºx��;���TJ������9�dG�
��~�6s,"Dts����>��r�Y��X���8�W�l�%;{��}d�0��}m�cG��R���秿������h,��#      �R�t��t�.W� �T�o�oј�5[oSQtn��Y�u~��7��{3i�Ll������	�s��g?�Y]|���:�~ڜ�M5�   ���������b�IB1ckkks%�N�4�x��cA��،�����$�����<�^  �;���z�^��W���ÿo�
��a�Kl�RB=n����}���՞0gA�v��V	       *HZE=�*ݣ�n�e���aF��5OO;���m���*�]
������Lm ���ӧ+�L*��˫=�P�~��B0��Mo�)����~X^eN2�%/�,D(   n�9Y��F��툂Y'�M�&�[�3��f8��Wj�v�f�,(1�����r��1���f            �>X�,���T�{u���K̨��y��|����q�ϤNTH�9�w:_{��4 <�愑�+O��S�ׯ��+��[�"~p�s�/^���>yє)S������V   �6���mI�c�hT����2��x������6ֶXLPd�Ykca�8<<��+I���}�'����C�b             �-��Bz\ݫZ) {���d�r�����Hg)��:\Uz�s�*�]�s� ��]A���]�TJ���򒪪*�w�y�0a�lMMM��w�[���iy���2q�Dy�   �������mO
�Ι��V(�f��O�Ř�GMM���g��KB��v*�	�c�1���֎��rƌ            �]X+���P���PK��ޚp�3j+�-�;��e�����t�Bz�����g�c��@@@M�2E�������3��+_����0f͚���?_�^zii2���Wt���P   �d"1�|���---�7�禳���ض#~�f(&����SP<��V�5�)�1�Jg�5ξǻL�������D�             l'�,��������T�E���`\1�6hj���,���k�T�r:FEg	�h�pLH3��& S+ 'Ţ��P��X�v��X��^���/��SO��������7��y��&�����T�ט��K�   �M�'E�	��X,fm�~B1���.�ϐn�|m�0?G��1�`�u�&��qs(H�ߘ횭P�             �̉C��z�F&
Sp�a-���
@�1��eJ8����Z_�dU��1:���)�W�sn��|n/�~�s� `^��b1����=��������[��V;�w�C��K�J��|���O��H�A(   n�=)�L�7�|nFFF�N�U[K�{W�ϴ�y��+��)���$���V�J<�f����Y�pX�&"e             �I�Y�	�=
�>���|~5c�u�8�_m ���ص�j���,O���}Y��S��SAag�o֭m��lp�u>W9_gP�"U���O��;^�f�Ќ3���X
�
�ƞ6m�.��BM�:U��w�q��+4w�\�Z�ʵq��ì�&L�W�I(&V�jr4�  �8��c�,��csRt]]!�����4i��kmmm��bL�'Hl�m�ϲ��iH�ǯl>?�b��ЦC�|�_ ��������AC��������W�OG
 0�jj�H�Z*       ؑ�rz5 c�J������R
;�S�ӕ _ ���s�K��e� R���+T�#�����Рe˖�=�Dt�Yg�#�H�6�;&O���/�\�^z�+�+FO�>]555�=	ż�o/\��  0�n��!plN�J��l�̺I(fl&� �b�q4[��րDL��;����;[��t)eBv���������W��w��"�}T�M�-��TX}�� @Y���zO����        �P �5�&��)se�P(T�1L�Ƅ>L��S&�b�-�6u�TM�8Q~�'�   `_1Y;��P��V(&�˕*UUU�t�l��ح�d2[�5 1���bV�7��              �f� \�P��������z��b   �&��ۓ��k555� m:��2��u�O�|�XL4U�K�R���v�v�P���z Rv�              ���  ��P.�b   ����!e2k�2Y���s���eel�1	�hoowm,
B(�lm��jnnV���b��muuu�팭�'D�              p3j �!�\�   �-�'C!��w---�B1L��-&z
�\9V�J���2�yl�sY�lG��v�f�k[�n�2v?�2              \ŌZ �k� (sq   ��'C����6��Q"�P.�#�9�3�	_���e*'NT����2nP��6#P&�C(��l�b��             �.� ��P�r���*M����   ʉP�b�92�^L,���]ص��6WB1A	(��X�HP��6�=���ħ|�f���{#              ��3;  P̤%B1   (7�чh4���z��lN�7̄}B1c��b��344� ���I(��loӰ{l��ɤr�A!              \�{  ט�Z@���a   ��d}��v���:�'mmm��322� �d2V�m@(�Dq����[��;�ϓ9�oBz&L              (?B1  ��PN�HD   @�ٌp0Y�b�����d}�ͭP���*�	����V<�z\�}�?�~-��G�b              p�   T��j��  ��FGG522bm|&��C]]��Ѩ2����mƌ�ĭPL:�V��f��ƶfr���SK b<���k�}              �a6- �6�z �   �ܘ���e����+c�^O�bB�PُY��~.���Ym��ᰚ��U�l8���C}}�"���p�              �S�g& <�P�r�&  �2c�>vW,��1�aL;g�
���J&�ektt��fu�1��	�zξ�üL��������b              pO垙 �B� ?���Q>�/�����/J�YW˥��J~RM(   e�d}�.3Yߖ\.W
w��v���͕����`�g�J���ieܠlm8lnϰg�k�V(��{$              ��ٴ  ��GQ����G-`_�y��k�  @�1Y��v��L�'36�ٰaC��I$�<y�*U<�2nk@B16uuu�F��?�|�`��bQ�PH              ���M p�9I ʉP   ���d}�~���Q��Q5�9s��k&���aU2[�AŘc�6#e�XL����|>_�b�$�             �M̦ ��P�r#  �r�9Y���Y�PH���mF��ĭ��Ȉ*�9�g��/�d2�\.gm�V��b�5a�=�3              ��i  P� ��k��c��Ď���?���ۄ@s1�k'ΏK���t(��DT�?Z�R�*jz��q�����J�;��rIU��Q@>(��,���@�c��C�������L�;���@�=3��x���3�̰_�3�<3�|�@#�A�K�.���������fԨ�4+����:U�ĔJ�T��f��ӥ}ꆟq'ɵ@�lǎ         h,Ӵ 4E��� �$ @#�HL��m뷗����g�JC�q�v111єuC�J��[�ZiG��{�Kڏ׬H         4�iZ �B(h4�  )��F7:I�$Ձ��/����P̆���������u�bꯧ�'����N��k9������X��Q,SYƹ         ��4- M!4�P  �4cX���>i�bVVV��A��&&&¹s�����z�҉�[RY7��b�����Φ�~�9�>�D��zϒ��         �E��W�  t����   �277��������v�'��\[|���;2�����ʺ�.	��)�
Ŵ�)K�y���         ��P MQ*�@#���  h��/��~�������[�l	\]�Ph�:��YXXHe�n9&��SZĦ�P�Ǚ����ndd$          �#@S��� �H���� �8i�g2�ԣ#\��Ci>g�I�B1�����F�I+���P���JX^^Nm�\N���Z��#         �e� ��  @���i�э����K���333�kkV(��Q_�|>t��"<W�b�R��=[�n         @㘦���@@����$I  ����|X__Om�l6h?i�7j'�
�P_�p\L�5��iK9�         �xB1 4�P�,}}}  �mff&��s������X���	�b1���~޶�������VWW�#�χN��k8+R֖�~�f�{         ��b h8��Yz{�� ��fggS]_(�=%I���S{���χ��5A�(
�����L1���{���dB�TJe}�         h<��  t�8,  ���гa����b1�;776m��:�����f�!�N��Í�������4��         @�	� �pq0	����  �[�C�1�@{J;���B1�C1��\�LҊL]��Ӿ�c�V(fqq1�������          4�P '4Ko���  �_����E�Di��~|>h�pL\__����2<<hO�5r�̙�֏瞷���         h�� 4�P�,B1  4B���$I���x�=�����	\[�P��\�b�y'�ߩ�xR<�Оr-p��        ��1I@�	� �" @�-//W/i�>���=��f䨝Ŵ�l6:]ڑ�\�x:Yι         :�	 N(h�  ԛa}nFڏ_���v1>>^�<���h}�|>t��_����di?~3�=         �P&ih8��Y�b  �����T���okccc!I��~7277W];�xs���#�����/����=9����)        ��f� ��! @��=�3���zzz���x�t�R*����ڞG�V(�b�@|M� S�s��f��\����CG         ��L��pW��� �!��2�L���ۯ�' @���f��0�PL�ÞGז����J �ӥڈ?g�ו�ҫ������Ce��         ԟIZ �j�������� j�� �P  ������G����3gR[?�bv����B�h}�pL��KM3.�{�^����)�J���*         4�IZ  :�P  �#i��޴��ôcG�"��Z_7Lb`c}}=��c�wtt4���k��ٳ���=B1         �&ih��Wp�!�bs  ��8������!+���[�;j�֗�PL�q�x�I�$��r-p�ٹsg          �O(��*�J�Yb(fmm-  @=�a�4C���á��?����O;:�.�������b�u� �vܩ~�� ��         K(��Js��>}}}B1  ԍa}�!�ͦ�~���v��d����Wk���ӥ�H��E}d�{         �c	�  �1�_ �z���Ku�B�hqX?~V)������������P���kNܠ�e� b���gbb"���~�~        @'��=��S�7��\.�f���� ��I�3�;��@���S�m�N�>�ڿ!�b�b�-��ZW.����N��C=��Y.�K-ز��         ��0I�M۳g�?�l��v�F�a�h�84�$I  �zMm����p��:�{����B1�3���@��&&&�+��v�g�4�=�6m
[�l	t�;�3|�{�Ke��>         h� n�׾��-I����|�4���t3=���[\  �c�Ν�a�Xl����sO	t�ݻw��{.�?��ko޼9�-��ZW.��`׮]�?�a*k:t(�v�{�7<���aaa��k�z�         hS� ܔ���?-��qJ��o��Z��8���� j��P�P  �244�����6u��۷���?�9�g��}�c�_�B���6f˖-�ֵm۶�b(&F6N�>��u����w�+�9�O<���/������#{         @c����MMM}�\.�j��V(&���7� �U<���ᥗ^
�Νk�z1�я~�:dMg��r��ѣ��_�rx��W������>��066
�B���	��P��w"G�	_����ڳgO��>�<1�Ce�<�LXYYiʚ�
         hS� ܐo}�[ٕ��?������7�  ꩿ�?|���X���['�T�����{O��n����O�cǎ�S�N5l��طo_�Ї>�>1���|'�Z�򖷄�[��n#���'�W��p��ņ�300P=��߿?йv��>��O��~����ٳ['F�z�p���          4�� n�����l�\��ҥK�I���������������˕����os�L& j$IR�p���?�������R�~�̙Ϯ���/^�_^ݼy���]�o�PX
  p����ѣG���?������ٺ}��y������j��7::�x���/�g�}6�>}���ݷ��m��Î;�/3�㲼�h>�`5��M6m�>��O��~��azz����x^۽{w�����$:_�}�?����s�=Ν;W��_��s�С�y��          4�P �mjj������~�ӟ>�裏n8� �(�c�L͗�sss~�ǎ  �	qz�޽aϞ=���E��/~��_����I����^����Q��[��]�vU��>�|�;��������<���K��ŋaqq1Fx7�=2�L��4>>����W�ߖ-[7.�F�9�y智|�q1�/�(��b�)��N�:U=�\�p!,,,�˗/o�{V��1s�-��m۶��;wV�7�%����;��W^y%���1�\���2=����T�=�\.l߾=�v�mհ         ��+P ���O?��>_���'|���@��.��ͽ�u�$��رc��c�  p��u����C�P���^h�y�{�=��~������G���n����z��!�����         @{����ʦv���f{{{K��600�7�/_~}z*I�?y������_   p������·���@:b���ѣ��?           ��P 655���������~��d~�T*�@����|���r��ym�����?�l�e   ����B.����7���b�yv��y��          x� 6��ɓ�Q��we_�$����w��� �*��b��t{���?������ϧ���9r���   �w�qGرcG��X��O~�����y������]�v          �7	� �!�������[��P(�MeS�0��R hI��b�jtt�,--�T�O��n�T.�yzzz����>   6dxx8<��ᡇ��b^x�p��Yј:)
��[ow�ygu          �9� ��رc�(�˟���������=5_�@�����
�\�/^|����y���ue��   ����P8p�@�R,���\�+W/���������/          ��� pU�r99~���U�������+۞��	� -!I��CR�}}}}����n���3���;|���   pzzz���D�          �,B1 \����'�$9T�ott��L&so�R�$��r�\�g�{&&&VΟ?�Q�k�*�����z��ş|             �-� �����R*��}�$IGGGw��_���9 ��r��*Ǫ��ձ�u���###�-..�]s�{��}���|              �6 ��*�J��l�����t�$��e������T h�c҉���{+W�*��q����������qm��t�ĉ�<�ȹ               -N(�����㏖��߫����{f``��׾\���O����� �b&''�zzz�@�$_���Uvm�f�5;;�`��Ƌ���+��              Z�P ��ĉW�	����+������J�҇����� Т&''���ɓ�;>>��r������}}}����n��ۣSSS�w�ȑ�              ��	� ����U6[k���L&��r��+�#���g@�;x��J�\~bzz��$I�o����W^y��7��sǏ���Çg              �(� ������͓���$Y�f�o�\����{�� �D�V�l��я~�ROO��^YY����-�r����              �(� ^w�ĉ�R����r9S�?��=[�wjaa�<xp= ��}��}qzz�T6�����qm����?~��_>|��              Z�P �+����yO�L&s~pppjrr�@��˾����}vii��ܔ���?��7��;��              �� j�8I��߰����C�ݻ��'O�|�r��/o�muu5W��     ��rE          B1 ��ȑ#_ ]�������y&  �$�  @�)�J�        �T�    �J�D(  �6�         @*�b    ��+            4�P    ܸb            �&�   �T.��b            h
�    �q�            �@(    nP�"            @�                 �8�                �'                ��b                 Z�P                @��                hqB1                 -N(                ��	�                 �8�                �'                ��b                 Z�P                @��                hqB1                 -N(                ��	�                 �8�                �'                �����3��>    IEND�B`�PK
     �k�[����  �  /   images/7de8bea6-aec6-4ad5-83ac-8e47725efc1f.png�PNG

   IHDR   d   B   �s   	pHYs  �  ���R/   �eXIfII*            (           V       ^   1 
   f   i�    p       �     �     ezgif.com  �       �    �  �    �      �w��  �iTXtXML:com.adobe.xmp     <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="XMP Core 6.0.0">
   <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#">
      <rdf:Description rdf:about=""
            xmlns:tiff="http://ns.adobe.com/tiff/1.0/"
            xmlns:xmp="http://ns.adobe.com/xap/1.0/">
         <tiff:Orientation>1</tiff:Orientation>
         <xmp:CreatorTool>ezgif.com</xmp:CreatorTool>
      </rdf:Description>
   </rdf:RDF>
</x:xmpmeta>
�[n  IDATx��]	�U���{�����F7�Ѐ���*h���$I�$��8T��c�ʤ�d�d��JU&��*Sٜ$f☩%JD�
���4Mw����}_�s޻�nO׭��������g������oy1|����߹���hT�.>����v#iK"�f���!�#���8/�`�9-���UaK�q�aN�aIZv�`��)m�rP�U�9��:a��\v�'�w]!74CQge!�,b�\A7���]w#mM!mNɻI{Yc�0��<�c�,
��a��G��u
�!OIsRڲ�|!.�,D:���}��n����:~�_T�w}�i�O�<�8U�<�ن��۾��˞W��.2���p j`�ۋ�� #����]7�F�9]���n����b��jőA?�m8T3z����`6�7@���5�1���L#�a4�*O�0��|w%B���8Z<��"�OQ�##a$�,�{�	�r�c�8�8*���p�ì��-�� +�#Tv[	G�	wc�~|�u6�_	�ǰ��J�W����{g�)Mt����CX2�6�9��g��4$T���;��;��� Ӯ��Q�U�$1N&��O�c*,�
��13�f��b�F=�^,;M�py��[�٤��r�
M����R�Rw�`	Y`�6"�5��J���E�6��z����
Q]�".��Q�����8�`6�-�h�z�l��v� pu��Ը�%#��eWT]6���I�P/��c�~=�fŘ�h�<�������ճd3�""߫A��|�z�ë��|/���@$q���ɀl.W*'R�w�IR��S��NJ9N"L@��?ǸO���XL�0R���ap+UU!�	�7�~�7�A��zy�လ����C5��C>�O�K%\�^q�g�d�R�W�p��n0L�HB�*XC�e�i�o�1�Buh9g��~�%�V��f�����Nt��겫a%��)�'��z\FQ����K��\����h����x�?B>���Յ�����\�%�b��PSmCo_v���V��rZ�v�I5E����C1TU؉��p��s����%�PW�T:�?������}Ǎ@(�h4��f��cH&�C#Qd2�z00��
8���=S��XE8�u�݌r�E�q�Y�v�1NH�BX]��-��:y
�Ch�)��:�FR��[#U�D�jcƸm�?v����l3�usF�e��q2����ߡ{0ؠ��`����Tfc�7h�2�,HO���20i�h���<�0��dΩȐc@���S�@=�ޑr� >��
_W���yאe)��1#x1��n�Mǋ��sT��u�ڐ#��B��[��b\����qS����+II��\��?�&�A�{��%�ep!E�nfB�:��ݻ�p:�t:�*s��r��U�2g�B�U8]�}��`~��26�|�T��>�0C����W�n��f;�C>�ZB����,�K#�����hA����p=q�����Hw'�,���e�%cApI ���<y\!t��eDx^���q�#�at�w4�&^V7yS9GqG]�e5��G{Y��l��� -I�1K8���0F�H�~�?���,����Ŗ<A����`NY� /�6���g��`C^nQL�aZĳI<��"z�c33��s�Y+�=fv��arYT�V����"���G���Ov���H�6m��l6��3��'؀_�]$���`���ǉ��F��R9RF���cu�jx^8MN$������*W.&&g0�2�2��~��w��RC�D�r��X�gj�>������K�c�X�]f"���.��o�\��
eG�T��x���k�rw����%�"�3b��n�%k9��Ʉ��r��ԉ�iR�Ia���COOrd�X���4!~04����Kh�^����X�X2&��,0j�N�+�_9_Ž�S�~
���Y�U�a$8�zo=�c�r�����D$U�O|��1�yꤧ��qy��Bv&�B8���D:��g]��^x�^�3q�n��>dHO���kE�������
�'�b:�:��WͿ
ۻ�#j�N�m4100�w�yG~3�-�v;���p饗J�����:U���3��1���R��'��	p�-�-XZ���c�zہ�Hf����BrG��i`È���R1D�Q!�4�t���ف֊Va �J�D���jTQ�G�5���ar�33wU�@�܁XJ�i�{�|��֭�33�I�^�3�TJ�Sq�	��$(�F�.fÖ�[P��Қ��ӻ/xQ\B�نFw#C��uբ?�/�r#���t��v!~�X.��@�"���W,C�x�0��l"3l42�D&1{f�"���N� aJL��gF��b��o>g�gg"��L�h�֒�%����o�i�&<��9|��Ϣ�]���0�8ʬeⷳ$������p�/���1 z(2��+�a溭n!<�5�������%fp;=6V6�D�x���ܹ���.�"�UY�0�9T�bC���Ð ���PSV�M+6�C�����U"ꨨ�G"#bK����?/b��a�j��K	��C���Рq(<$��sl_�^���ƌ�;�U�'f��-�S�t̛7O���>L�b��0����rfB�94~[۷bm�Z,�Z�n_7�D �ԃ�!z�R�����Xd���L��}gO"�}��>�c�R�I�W{,[�L~��bO��ߝ;wb׮]%�rf&"�;�ueuBtڏ���;�{3�������v4�[G�B.�C�*0�6����q�ݻW<)6�2`$�����Du��3��`,<�߼�X�A������g X��� {�6�#xy\�R�6���IT��mVLf��I�`,h	�������R))��a��!��F�>:���Ư{-���uk�e5���m�iarAB����r���<�~�h����&T<�^L�*Y��w6�z]<
_C�,{~0����Dg�S��>�]�pGBGND���=��@����#抦+Ļa���o7"�Ȝ�����h�9P�^M6&�ug'w���N�������-�>�.2�rX�m,2�*op7`�W�A5.]��˰�gϩ�TH x"���@ޜǜ��Z9âAS�*�}֓w@jN�*�tm��L�afn��������!f��?e�(����h<#���9�4s��+�H�ϐ!��C����x�`l�����	����L����g�!�\R���Ig�8��y΂N�+��M[]��B/�p��ڊ�����6�s�=������|��1���G��f��b�N��#���;wZEBlZjZ��(vD���с�a�@veY�2ll�(㐅��b�;�0��i�x�8ĻԶ�WO���*O"-kZ��6���\��Z�@RQg��u��	Cd��hjIXp��p!�[����f����`����3��C��,�c���D��0K`� ��MN�ӅK�"֚)�����NHp������_�fM�f�)�9=�u���XGi?�� +"�7�t��ȒADZ�S�}�7��o�4.?s�aWT�(��?���ق9x��XV�~��er������)��DB�B��õk�ʴ.K͉��u��ˬ��CNX*l^T9�$z�JN�a�p���S]]��(�!֒������p|�9�Ygsn�#�T�1�a줃Y��9[w܎��v�,�gY
jjj���(L���uR����O�����(�/�Bm�[�H[�3~~jJQ��k[����#5y��
�d>]�GWUU�1�L�ϛ�k��Μ�T�-K�T"��uM�pB�Ф{Lt�ۡ'��Y���hmm�ē�rY�X���.�gƪ�;�;�t[WY����Kj�8'<p��믿�����^��h4����YԴ���?� �R�P���s��(��wvj�	ӑ�6g/������԰*[�`�̭�'�N��5 &d�3�~|�RE�z�8׃��4*�k��Zθ�:��A_{?���%#��y�p�9�t8eĞL'U�'��X:x�'�8�w���H�R8-Pp���Z�p��b�M�J��^/L�Vf���"����'��P�j֭�;h�r��N�ө�/r�礄���9�� R�3����+�wC���ց������؍�7�x���,G�B�i�HR�$��A93q������l-\4fd��:^�x���Dw_7~�����M��G� ��b@�H{�s���%R�ϕܯ�:Cv8uHd��6��k���j�*(�nչШ�����<r�#b@9��#���,��TA���»6�qo�^��z����X�-�[���H����.}���bD��"!��Hޱ,E��s�I�K�R��O6�;�d���i���u�oP"7����r�L�����|�|!cD��w��f���5�U_2�}�1����G�rT�����C烺bpU�*D�D��=����6����Z�x5�*���g��[֣�V~J���TX+িH*b�a��k�5]�����b�W�^H��o��-����?�_<���h�"49��q����4�{ٽXQ����i(�,W���<<F�Kz��<�%'|�po������� >������ JK�Kp�^�VX����tUK��dCq1a"p��N!��n\8�BNF���T�j�"R~��'�2�����U�i�|�����<�s�rO]7��9 �3��]����W�%���G^�;cߚ+�%��K��b�yr���~�_�Jl+���a���*yy�Ǯ��u���tY3�����W�BK�emQ,����?������/�><2��e�Y_��ax��>Z�L���X����zdÁ���.�x�+�U�?b�v�`��y�fܵ�.ɗҁ����?~����6�͞f�}�m�84Œ�3�8��u�2A]{��
�>��o��
&V���$1�d �d�(S&o��j5Ye�ˣ�+�D"�8&���~\U�l<0�ph���sj�\	���l�d��pV�]-�B��;���ϣ��(�����P�W��xu�[�o���W%?�cU=���i(�D�tV�s��1Z=�2�Y���ό���ے�󹔜O�r��b8{�Q��������/���0GGFq��<nϴ��^�Ep˂[D��e������薱��,&����Z=/��\���0#&��d͹�)�+��}4^�ۡ:$$#s���S[W{�tV����sެI1�''��h����9� 
�<L���x�^�=n t��$��:C �:��*���cccbG�˺�(C���;�~o�	����e"���eG�˨��*�P��L-����o�k�����$� ���H�Ux�&�͜-ȹP|��esΑ��d���ק�=�;����"!����Aڢ(���*�K�`U�j�����x��^B������!��Hޯ����!�I#K�n�)={O�'*.�g�C�E���{�K�o�'��oO��x.[��7��M�j(�*fo�ĉk%���\[�+����zo��6sc�*��,�ņp[XR��=�N�S�b�z��|�����w���I6���j,�\ ��m���]�n�t`�{#��Ll�!�SbXd9��$�����K/���.�Hz4�N&c�r�G;�ʸr6���
K���_Jrf����K���>�h#6Ԯ,П~�~�O~	�ӻC$���⭡�^IXдi��ɀ�"	��9Yz�^�rO��t-74�f��	�b����WV���α�׿�W��`Z�f]w����6���ͺ�l�";�0��ڄ9zV�+�-��ό�t�[o�����a��h(���t9��#
��"�ب�wE�aZj�u���ɺ��=N�5���j5u��4�z˻�C�s�}��v��Ų��Y\K����/�Iy��'I]}O���<��z���}7|?��?�QB�zŤ�Q����]xz�ӳ
��HL|���\r�H�T2#$%��[�װ(oܸ���B@q7'���4^��F���֪�}��f��7�w����.�t<dP��Jb����-w]�nA7ｨ�FD?n�1�F{A�f)$,�U�*xN$	�����`j8�f��<�ؼ �y �Oe����n��이��L��S��0�����%K�H*%�f��J��ҥKe�H�'��80Umlߵ�=�%Ǟ�sv��ŋe�Fuu��É�ŬVr����r�U�wl�HG��	�ۻ���y�������3��[�T��2�l�� 1���÷͍\:���x�����)�Q�l���Ɲ����{>�0^3�q&���EOJf�74xN�YGʦ���=���'�.�=9��Ib��c˳�:�߇��~�÷IK�3*L���@:
V����K��C�O=�����'����Zn4�������Dy��c�s��l�}~��L XJFͳ���S�,�ng��b�0�a�>�TUWU�*J�ܭ�[Q���϶���Y��E_Cw���bX]�M�cB'��s��� ~ֳ��s���}&*��:�\���j�Z�y�oO�+6��e��y,�l�::�EԈ1������R���l*��țb&�/�f�y�����%�����6�U��R�4f3���[3�&��6ILVF�Zs}�eq��F�G�F�#��t\ֈiYʹ�/��-�VQ�:	�A�o�!b��!��W���~�wdW���ށ��L1���G�xQ��&)r���/�~Q�\��<'�D�t�u���:����uAk����Be�Z����_'�r�K���x�՗�!�����B�1�y��;v�J����3��y��+����}�髷������W��?F�w��]A�y��f����󹛖�/?���8>�i}���x�!���K���Z�8�;��솽���
^d+U8O9mq�"�󖓷/�!���r8�	�\�M~�;o�5�k�;�;�#w/KPt��:�����r.�+΄O��Ϸ��<�R�223x�A�~\q�B >n��Fa@}}=�7�:c�����o>���#��$��ƫ�'�~q������\�kw�1{��4J]���{����mYӂ�5=	���ţgeϖN�U 52��    IEND�B`�PK
     �k�[�I��t� t� /   images/89718c7b-e32a-4492-aa2b-d7960b76d502.png�PNG

   IHDR  �  �   q�y   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  ��IDATx���	�\U�7���[�tX�6	k l��tWw�� ���PqQq�?g�gtt\`@��m�QD�t�"#��2���������DGgT���n���<��J�t���=����n�}�"           `=�           �w           ڂ�;           mA�          �� �          @[p          �-�          ��          h�           �w           ڂ�;           mA�          �� �          @[p          �-�          ��          h�           �w           ڂ�;           mA�          �� �          @[p          �-�          ��          h�           �w           ڂ�;           mA�          �� �          @[p          �-�          ��          h�           �w           ڂ�;           mA� `�x<RE�,�D{���gYY�85u����9h#Ͳ�T�����S ��'�jT�:�<f�>F�ZZ��gWy� ��G ��� ��-�����4���#�N�0�ǗG�?��F��6?�cʃE�����~����q�A���e�����w߼�{8&@�X�H����=�֌�k� h'�z��D{k��?��� Ƃ���{           �w           ڂ�;           mA�          �� �          @[p          �-�          ��          h�           �w           ڂ�;           mA�          �� �          @[p          �-�          ��          h�           �w           ڂ�;           mA�          �� �          @[p          �-�          ��          h�           �w           ڂ�;           mA�          �� �          @[p          �-�          ��a%�7Z>�]~jV|l6ذ����_�li����x��HEEk�z         ���G�����	+^�5�ٌX�����d	���opg우A�-���b�ȶ�&b�I�6����+��"�V��,[��#�|���<<ZEk|����o�fY����          ֱ�i����Z9��<��6�d4W8f_]���#�9�bt|d�k޿<O�"[�ǀ<�1�t�,����H��i��#=��o����]�׶�F���������(Z!���t߯����G�#~yO�(         ��h⦣y¬��n�ȶ~ZĖ[G�l�Sk�����6�4�U��?�8��E+��������{5�),Z��_�;�9�N%�N�}���S#�{d+�1y��WA+�ߺ�u��{ǟm�?4�15[���˺��<         𗥭��4u��v��<S����W�FGj�λ�����Q�������;o����(�ס�S]li���v�+�ݧE*+�f_U�;���yY��C�,7�⧷F���"���        ���j2�����;�i�}"M�2:RW�򟱬?6�m6F�6o��h����GQ<���*p�:ƍ�p����鉴�v1�M�4���e�>�dٲ��E�Q��/         :U�n����G����=Gs�cV+�󮑷����ї�{�-�b�P4o��h��@������&��gF�{��f�FtO��rc���)�ʟs��ﭰ���Q���({4         ���wG��Gd=������kH��p�j&�
�/[��?��o.�(��Y@�p���Q5뀲�����jjux�s�h��H4TnJ�͡�",         �ݥ7��;+�V�p����j7n��pުX������
�_�"�������:�r�xz��v	ְZ-��}�UGѺk���AĒ�         �Ƹ���h���3��+X�F�����j�G������;�o�?ny+�~ࡑ�8%X7Z}��YY1<<�ѽ��E���f         �:�e��=3��G,Ϸ	��3i�"���O<-�����|=��;��X�Y��λFvȑ��9d�.+֣� �u�hŃD�ܐ�߸.�~         ���M7��C";�H[m�_i�)Q{�Q<�Q,��o]ŭ�#�"`]pg��h��:|�Ϊ���A�|R�Ǟ���G���,7����        �����>�7�V�}�z�΃����"̉������o}5���]�Y�Y�ZwSeG���G��*��P�zg�Vq߽���u�(7�X�4         `u���g�1'E�n��Z����^ټ3����h|�s��wX[�Y+�λF~�q��>x�N+�)m�m�g��q�D�?�ͯ��(z0         `e���Dv�a�sӦ��4z�CF���Ń�������'k��;kNJ��D�̓#�u��s�..�cO���c���oF�K����	         ����:�g���Ftu"�"��?Z��{+�޼yA��"�����7j�</Ҕ�A7>�C��l��hut���x��         �?�|R�ǜ�!G�v��s�����E�Fq�����碹h~�S%��S�v��ygF�c�`�k�����E�߈�5���        ��+M�$�g������>Ƥ]v�څo���E�_?�����Y-��=#?�y��c]mE�}�����u����Q<�h         0v�7��y�vLĸ����ʗf��2��.���?1��V��;�$m�E�<7��疋0j|w�Ǟ�!GF��ό�ݣ�         :X���	�g�i�M� �6#����ߏ�g>���	XYq�#?��Ȟuj��	цE~�9�=�1��D�x(         �<� s~�ّv�9�/J)��9����׾�/~.�'�<w�T�3��/����+#m�]t]��h޼ ��H��:         �����������2��V��cO�|��1r�'�y÷"�"�p�݄^������:�����=3_�l4��&�1         TP���'Gv�)���V�擢v�Q̙#�@����;�[�G~�1��;3b|w�SR^ȴ��l�c�����        ��H;�����J{ό��}0��K4�|mD����3i���oBS��Ii����wE�;_��|<�'�         ml���OxN�G��ek̸q������;({4�#���z\Hv���&t�hwX+�����"ߧg��{���        @�iuٮ��呶�:`mI;N��e��u�D���D���i��Q{ɫ£CXg���k���׿���c��        ����sumg�k�wJd��b�o���c���X�R�s�����G#�T��;♑����w         �O�n��sw�����v��+����S4��oE�M�cT�d��_���z֧4y��z�{lH         닆������8<'Ҍ�h|��Q<�`0���A����Ͻ`4�m�R�����أ        �:��Ĩ����f��E+뚽��1���Ƿc���XҺ��#������lf�{����{��]w         kO�i��:��"��:��l�Yt���h|�����"��`lp+�'D��WFַ@[��Et��1���w�         �yٜC����G�ж�,�O�����л�x�Ѡ�	��i��v��"M�>����v�y��e�h|�C##        �S���"{�Y��̀��z"���1�+���σ�&��ᲁ9��s~��	U�rTd��#�}s=         ����Q;�H��P5i���u��b�C�����%����#�����>��*M�3jW�'F�yy?�+         Xui��v��&mPY�Fo�h\��Ѣ3	�w�,��s_١Gt��]�]ox{��-Q,
         V^�{ft��ڈ6���"?�ћ5F���##Agp�0�{B�/Md��:Jylw]ti�������        �'�tX�^�\d�Β|x�&m#�{KĒǃ��l�A�f��vѥ�v�%�#��NP^h5��!��HDQ         A������t�*ۧ'�.}G��҈�:��{��frt]��I[t���gF7>F���f         �'�,j��O�ti����7�]��T��{H����k���lR�X��="j�b��h�         �,��E�G6琀�"m�Ut]��n��yOPm��v�%�^󦈍'�5�~F��;F�����         �j����5���s&n�׿-F���(�=�.�
KS�.�o�Q�X�����o�ƻ��K        `L7>j�.�}zƪ��F����_���$�^Q�^ӣvѥ�ƺ��!.�,�L�        {�'D�U�E���c�F�5W��;/���#�^A��=#�����'�=��^_nH�E,[         c¸q�uѥ����R�����y������"�^1ٔ�Q+?p���X+e�*�tOQ?/������\�����gY�l��/.�li9<^���e�r���eu�_7���L*�����cY;��y��e�fD����\12         �,uuE���E�s�`�y��V����+�����r>\�)k�X&�y>�Ÿ���cy^w��k�,�-Z��Vư��P�w.��e���5n|��!�7_�=w�!�^!i�����+F��S���n-7����G�F��F�qw��e�^^��|ppp��{�Tn\����e�blmT)Xmپ������?om]        @G���_��Ȧ�OYQ��e���E��,�n�g֬Y��o>88�U~���������4���)�i�\G� m�Qt��M1|ū���_� �^�i���+#6�8X-?-��pC��?���~��y��5��_�^��:�/^QW���n�a����z9ݿܘf�������*�����9���G�+�        t�,��K.���_�Z*�Ƣ(n,��/]�thΜ9����̊Ƽw��o������*�u�]wo6�����e��݂U��Ĩ]re����Q�wo��ܫ`��u�["&�9��_��WSJ�gY������F�� ������E��]���ud��P�<.xR�O�|ɒh|�        �I��4��
V�Ҕ�����������������OV��Z�-^�x������La�l�6��J�n�<�~���x����	���	D׫.��|R�n.7�m4_���[\΋���W�;o��֍�񧗯S�O(k���/ߦ~��	        �N�wJ�<�ʺ6���Z���3f<��9~S�oUQihhhf9U��'����Ui���vѥ1�Ƌ#�X�/�v��Q;ﵑ��)��~R���.������4:ܴi�-��۪�����)S���/srY�.k���O}~>��         U��: �����Z��r�����kӦM[lE#�E+�ʛo�y�F�q\,���/i�)������;/�h6��$���jg�4�}z����}�?������V<z�V�q�?��C'�����ܲR�\JQ;����}Ѽ�         ��l�i��{�h&�?�L)}�?�����N��-3gμ��ת�e������6	�(���s_#��A{poS�3�E6����|�(��_={�lφ�S�N]Z�m���Ю���
�?�����q�"���Q\va��:         *e��Q{��#���?���,��c�z��������R/|U9�\�O/J)���=:����/_��64��yg�Z]ʯ)O�����[<���ޟ��k���o_6q��3����z����M����c���x��         ��7���/��h�`�me���G��ܹs���z��x9|�UCCC������_Vc\~���ͯ���Ơ�����ݎQ;�|��h�P?�h4�;00pw��Vl�iݝ�hѢ����r='ư��ɑ���y��f         ��,���.����b�+��)�����~��`����M�p��dY���=}A��cU��u�1|�/���_�C���tO��y�D��1lYy��D������<e�F�Jr�U���s�����c��f�G��S�q�g        ���'�����nJ)��^�)X#����*��/^��������ye���j����������x���=����] /}U�m��1j�܀���h\����6�����o(������)���|f�A��ώ�ۣy�`         ���wV�Ϝc�PQo����J�V̘1�7��E�}��l���?/�b�x��Q;�y�[Z�
ֿ�w��V�6���(�������z���`�������<44tR�|WY��X�e���UQ���(��u         ��V���Z���M)]����rlk]�^���^�p�;����)<:Ƙ�o�ȏ=)�vu��	���4�7�g�c�EqA�^�>X��M�u���7�p�W���/)�,k|�iÍ"?���e�        ���	Q��ulc̒�һk��[f̘�X��������:�(�w���b�O>3�w�ŏo	�/��m�͢v�ǐ%��r#zOy2֫9s�<R�l�����wsh�َS�v�c��!         �A~�9�&�cIQ_m6�/�;X�z{{�t뭷~�'����ݼ�|�;Ƃ,���\ïyi�>X�ק��v�y�&nc���:����?��R���,��O.�V�{��C���x(�E�        `}���Ev��1��.�����ޏ�c��iӦ-+�7~�(������X��q��;.m�y���Qv�1���1�u+�E�&�q�P{���W�t�M߭�j�/��b���1�ڗ�G��        `}H�o1�4w�H)}��W����6h[��EQ���S���^�41:\���ӟ�o~9X?�ד��Q{�Y1F�T��+:�S�fͺ�N)7�-���Yt��ɦQ{�1�7��
        X�Rm�mc��EQ��^�*����?�hѢ�6������p��ώ���/�	�=�� uuE��WE�n�܄����7o^#��V7�rCZ�h4��ܠ�������F�k�         �R~��]�;]Q?(������
*�����W]u��)S�\T.�(�+:UWW�ν �/� bd$X��׃��3"�qJt�{ʍ�rZTڊ�rCzC�|]YYt���gE�G����W        �.��v�lޙ��ZMr/���ߢan�����m���˲�s�|��Pi�]"?�h|����%ྎ����Q�E��NWW�)3f��M�VlH�.\��ҿ��͢���p��1�Ƌ#��         X��,j/xy���m�]z �tZoo�ׂ�������`O9�LY�E�ʏ91��o��;�uG�}]����l���e������;wXu������iߢ(�)/8�с��{F6��h��W        `m�;&�n{E���h�000pw�q����W]u�QS�L��\^\V�N��Q;��~��M��u�c���(?�h=��C-)�⌾��k��VnH�<��~�����N}^߼ ��        ��!M�2�ygF�J)}n�ҥg͞={IбV4D~�����EQ|��wG�I;N�����k�uC�}I�L����D�z��g�����	�z��r#:epp�'�Eȥ�i6�0�^#�,         ֆ�y/����===�L)5�1����󃃃���+k��0�ɧGs�Q���`�p_R��_1n\t��l4��������(�ᲅ��� :�|���l`N4�o        X����F�3h�(����}<s���������c���r��$��G���[_Q���Q��v��>8Ҟ�D�I)����u�����Y�ȇUN�.��n'�O?;��F,}"         ֈ�	Q;�сO)�P�׿�Y���?�?��<�[!����#���ƹ7}/X��׶q�"?��i�M�?�,Yrly"z$���//Z���f���r91:D�|�ȏ=)���         Xj�?;b�͢�<�R:����[��700���ŋ�>22�Ţ(�R{�c٢˖k���Z�?s^�I[F')7��.]z�9s�������E�=��l~�\N��}b4��Q���         x*�V�D:��aJ)���{S�
3f�x�;�8����(��9�'m��'D������lo�c;Iy��v	�.7�e�COO��+/V��ro=�������yk         <�s^��+:�oSJ�����0��:u��[o���%K�\U.���{��ƹ���kQ��Fñ��n��s��p;U__��,84˲֣f:�9:٬"��uѼ��        �:���G�7;:��Wtnn篚6mڲ[o�uޒ%K�-�GG'��)ύ����kI�m��Pl�ֲe˞պ�&�I����288�z��W��0:@~�9�|���f         ��,���s��<�e�Q===CO�r���O?~��EQ �n4�q]?�i��	��%�S��Rt��&L�p\�^_�����E��l6�+��Qqi�]"��?�7}/         VE>��H;���%|fOO�V��ٳ�,^������V��9Qu)E>�1��K�5O�}-H{ό����!�sܸqϘ6mڣ���������3����ʢ�j'����l        �JɲȞujt�fJ����o��3f<6��g�y��r�{T\6mFd{M��O~�Y�kA~���!�/7�c�O�����T�ׯ�RN�U����f��         +#;�鑞69:AJ�����/�����.\���Xj=`���|ޙѼ�`�p_ò����Gt�%Y��!򳀧�^��mppp�r�������D�ߍh�        �ߔ�"���EQ|�^��7�)���k���dY��r�ATX��gd�{��á`�p_�R������^�C�===?XCy��6�x�]���Qai�Ev�!����        �o�><�V�D���w�]��������CCCgE��r����ψ��ҷ��!�e��"�KT]y�xK__�5k�ܹsG�ϟ��<���NQa��ώ�ߊ��        ��RWW�:�{���<?}޼y��5����󃃃�rzQTX�25����\4?X3�נ����ꊢ�����k�����-zV�ټ1*�X���V��wP4���        �9�Dl>)*nIQ�fΜ�P�Zp�]w�fʔ)����Qa��Np_��אlϽ#�{T�/RJ��ˊ����g���Ћʋ�OE��ǜ����G�         �SJ������(����9`-ieV�ϟ��<���NQQi��"M�3�;n�:�5$;�����f�yR��kYoo劉���?gEE��v�l���Ѣ         �Sٌ�H�������X�X�`�iY��GT8ۜ}|��W�}M��A�V���������e���֑Z��������ie}�s��;        �dG��J�^�����߸p��+SJ�FEe��E�z�(�7xj�׀��ǗGevÝw����uhƌ��Vō�r\TP�{f��D��        �%�Kd{M�
n6�����<`z��G�4q��Ê��U�e�y\4>���p���M"�������y~Ƽy��Xoo�P��r3�2**?�Y1�w        @K~�	Qe)�����_��͝;wd�����y~K���|X4����GV���S�|xĸJ6�U�3gμ'`=���y����1�E�~QA�~E��ǣx��        �q7�l`NT��;�S�O֛����.\xqJ�CQE��G~�a���5��p*R��â¾S���)`=*7��������PY]Q5�Z�9�D�/        0��Z�Oe��˚���͛�X����G�����C���C���W�mu�VOeϢ� �kz�m&GE-I)�]�O�]��h��(��K���C����_�       �X�j�{��QU)�7������������q���ewT�6�#�cZ4o�q�zܟ�l�QU�����ޟ��G}�7���r�{TLz��H���O]�       �X��O��������-mb``�����+���2*(|D���jp_]mY}������{��ܹs�X�h�K���7���GĈ�;        �Y�!�m�[�yӦM[�F����pfT�qn�?'����({4Xu�);�Ј����������m������+��D�dD��GlF        0�6͝U�R��^�W�1)��<.����.*��KQ5��E�}p߸.Xu�)?谨�/���~5�M5��<?����*imFD��        [��W�i��f�yq@����npp�k�􈨘��ã)�Z�WC�v�H��4\Ņml``��r3�?�r�j�߁�p       �1'�}PTԻ����
hc)�WE���V�.���.�����_�F�}5��iUM-7����<���h4�*��E�d{�i�IQ��         ƈI[D�u�����<{@����mpp���쨘�N4���`������VAO����%�fΜ�P����^U�e���E�"        0f��ZLG����
��7�ufY�B��p_�(�qJ���G�E�Y�fy��1aw/Y��e�t˨��܌��        0fd��
���'��������X�p��RJ/�
I��i�Q��/��'ྊ�@%��?�h4�P!ӦM{tpp���ROH��iҖQ<��         :[++��L�
z˜9s	���ҕ����6�
i�Ӹ�_��'ྊ�
���Gf͚u_@�L�0�K�,yU9�<�"�������_        ��e�8����.[��S��=88��r��lց�H�}���G�frT�HJ�}���p�����%Q!if��;        t��g ��(��={���
j4�����Q�t�v�H[o�}�+�2��v�fԣ������y@E����k���;*"�}Z����k@        �Xli�ݣb�6�۩������PNO�
I3z������p_y�EQ�7��f͚u����g�c����Z-�i3�9tS         �)�gfD^�fQ�le�*��l�#˲J��}����/+�Zg��i|wD�+s�|���oA@ŕ��{RJ�	���}��        ����5�-�<_@����/�~9�?*"�Oĸq˖ON�}%��1������҇:@__ߏ���n,�bvTD6�/        ��R��=Q%EQ|����'��Q��{+ܞ�9=���''ྒ��ި�������ceU&������Q��        t�l��#m6)�$˲�t�e˖]5nܸ���͢"Ҍ���"ྒ��3�b��^�?�!j��U��í�h����O��;        t��O�2��[�t�5b���K?[N_�M�F�2�W�&�E�zۨ��(�iEG�1c�c+6�s�"������_        ��d�O���T+�A���G�,�L�=m�m���D��M�}%d��ss__ߏ:LQ�N)U(�^��X        �ɤ��Q%Y�}*������288xk9�FX�<w��{F1tS�	���V��|@���7����U0q�ѧ?����ٻ�x���~��3soH��P֢Ո��M���B��Z��U��V��Vi�Uq��Y��RDܢ��,�ɝ�!@P���� ��9����b뒄 Y�3�~�^��3W�{g�<������         zC��ƻ0g�8�Л����G&�n�m�{%���:�+�E�Z��)��m���Q�p       ��a����U@*���f3��{~M��
�{3iR{�����Ȍ3��]s#��{]�~|n         �!��{UUszԁxU��Z\/��{�Y��`��X�~����ϣ�w)��)�tJ@�1c��v�}C��=2�x�c�        �W4�
�_3k֬KzXJ�EQ�p�b�GE�ْ`��Ino%�>����_�3zX�Q9�v��� �&2P<��S�F�Z        @ފm����\Eqz@��';���Dc�GG)�A���{FFn�<�ǥ�ά�,�u��{DZ��         �V��x&(UUi�Kϛ1cƢv���z�����>�	�ߋ��{EF��v��q�W�>w���k���@Q�#�        ��gdduQ���nv��j�U/_(�j��U�oHs ��?2rq�#��t�Aw���z9'2�       @oȬ�����+�@J��$:��{��xF9�N�n�P������-Jk֬9?�����Mm        @����\����EQ�SO���	���a�t���e���2���ٳg��?.�L��%Eѽc         SE�G��&c����Vki�|Td��+p_?��,��W֮]{ɤI����I1�M�6��w�t�o        �S���FL��X�bŊv@I)]TE6���G��	�o@��"�r~@�={��v���.H3#��)�        �)S�R�3g����m���@��G�'�!�>$rQU��}������.         _EF�BMs�G�Fc~J)rP���`��7��O1Z1<<�4���7a�F&r��        �a׬������������rۘ�v�)����v������J)]^�*�����e��9p       ����q���
�3�,m�ݾ���g�W�.�����O	��GNa�F��ї��]�|��Nd���        ��]�X;eʔ���{wL��{WcׇDu�5����Э%��V���о��j]U/\�`w        �Y����
2}����)�Lm�q���:	��Ϯٜ���,��_K"��{L�!b�6k�        ���S"���XЧ��UUE�]5�]��h�s��2^п�8�TQ��J���        ��)�La䒩��`ll�f�Y�q�`���g�����k��榀�u]d���w        �д")����ʕ+1mڴN䐑�.���7�?��%�bt��^���(��o�"ӲyD        �{�����4�k�Ԝ9s:�V��8z����i��#���n�7��u:�k�y���V        �����UU]�ߺ�Z��	���v�ERJ7���+W�0-���        d�ȧ�{�:u�\!��ȁ���%�>�v�E�>6gΜխVkE���R2��        ~O�I���|���k��-���O�}]�(�n9��jY �����+F        ��|�[�B.߃nV��膁�?$�Ŕ)��葉<���y�Z�=b�����        ��L���)��EqkJ)&�n�}򔈕wH�}��`d�� �)��       @���lr�2���("�(�'m�E^!��}.�t{��S'        ���lF	�.�B��#2�D��Ż�.upo6�k�\��X���D
�        �Is˔��>WU՚,��F7W8���:H[�KF!Ժ��s�� ������        ��\�[v����n�6��{�Ӕ{K�c���2�X�a\߃bP!       �,���)��f����.Dtp_7�u��m)�2��հ9E�G1��       @�������r:��
�Ż�.E#r100P����:Y<N��         C�<r�EQ�}��tR&ܣ!W�.��Rv"#y<�6��m9�d��         ��O�G���WŤl�O	��CQ�s���% ��B        y�$�^UUY*،ʲܦ(��B'��3[���:��B��NG1�凜�(F
        d��+� ��m��M@�˩yt�'��%	��KFK��P��{��4�6        ����2�,lN�lmUU����D
����:���=�4%��u�:�        �M>ٟ�}.�lmG�p]�ס(�����9P�         O�4��)�ϥ���֦����p_��fM��hd�%�ͥ(�,n���|�        ���epϣY(l^�dk��[�(�uY�귝��x{#��5r��         ��32�O�6�<���p������"��U�}W�;�D��c`s��E��΢���;        djE6�<���u��EQ�D��Z����ztO[�k	�c_|�&M��-�        Yʧ��6�Vk���a�Y�VQydkW�������s���Ƕ�f��RJ��t�{F        �Q�in.����
/�S)�=����Ͼ��	��G���Ŀ����Ǫ�ʢ�[�        d)��OUU{��;}�(��"��%���x��ŋ������C����#        �Q�in.���3�O]x���i���
���p_�"� jY��ǉ\Їry�HW��M.        �{��*��O�P��&O��gd"�%�>��n�%rQUգB��>Už���q��        �'ݶ,�*#��@�*���R� -�'���	��G�����~��n@z|d`��LU        �����<82�E�
6���_Ed!���%��-�ܡ��Z��FnQ�         k�P�G,X�`�<pY@�)�"�I�p��ףX���v[n4"�|a���W�         o�P�<��E�z� ���+��H�n	�M�}=��X�;n�b�]"�j����#)�<�#��B         $�&��F��p��,^�x۱���"��e�N�n�r�o"��7�1T��HJiV��w        �YN��(f��5k�7j��[d
7D�}�o~ţ�xR��fG.��        �W�(�RzR@�i6�O����A�)� ��~q]�q�C1��\z饻u:�="u��n�!        ���x�x(�"2�w��z������A��nF��p߀���S��R=y=�hll��E7��}4Ѫ�        �+ݽ"�e;�9H)ͮ�S�@7C�n��L���O�}C~q}dd����?���F��ͣD�On        ٫n�6���ݬ���v�q��Sd"��A��n�5�;#�m9H)���z?42Q]M         �K��6’���(��?�L�;�G,�=X?�{�n�>���9H)�e=��,X�W=��p�
        zC��������=�����q)�gEY���`���E�q"�L���i�Vk����ʀ�h4�I�        �ܚ]����z��ŋ�;(2�4ͽW����k"#��b��z>=��E񗑋5�#���         �~uS�ڵ�&E�]�C����t��m"U^��B��^TK��GQ���;=lɒ%ۭZ�jNd�����?�         z@��5���3�ϟ?e��٫zTJ�9��j�O�p���V���Ql�Cd���͛��9s�tz�ʕ+�S���D�ْ         zGZ���|���U=�ЃZ��`==/2����뛂p�7)E��O�:02��;���z>7�E���H��'        �tՕ���(wzTJ��5�sd"��ckp��S>�(˲[���9�\r���th䢪���G�        @/�VUD��8l�������w�Ms{���F�ꋩ�����k�Zo�!�f�o�ird"�x}�J��        �K��+"��(v{ddbj��9����C�.]������&2��
�o��q�U��Ƣ�L�R�s���=���_�~�Q"        Ћ�]�3
�GJ���p���y�ϭ�E.֮��ڥ��p��p{��Ϣx��"UU�S��CZ��>����H���        ����+"�y�E��<�������T���Np��7R���Q��(�CFGG��>�7tQ����._        @�)��YU�Fd�Q����==`��{�������`��o��v4_���H���n1:2 s�����U/�����4��        ����t��Q�od�Us��}��^dn``�SJٜ0�.	6���FJ�_�ۢx�N��Z�dɇ�O��6 c�o����B���H�        ��nX��W�}������|J@Ɩ.]������1r���H7�l���R��F�x�3"#[�z�K��Ā�������        �]�La<�%��F�qD����˗���)e
����Xm�p���^�/E�2�p�§�Ӂ��t���>         ����g+��nZ�"�4s��g͚5? C�5\���Ff�e�`�	����EuE*#����FGG��d�(��GfR��UU        �ê*��G��O��ܓ�p'K�v���鱑����O��>Hw��t�eQ<��IJ�!�N�.\8���zvd�q�        ��ZxQ���y�̙3��n&���#'���VO��>*/�qdp�\��������4��v��I]�*�       ��P]ڊ�zU��DF�EQ���_�����g���S"3������}�^��R�sy�u����tP@&Z��~����Lպ8bl,        �>�vM�E#Q�Ev�����Θ1㲀|�?2��Ƣj_�7y��'�t��HKG����̓Z��!���gd�{(#��W��Zuɏ        ���P#��{#���z~A@Z�ֳ��/"7��F��;�o�.F�ܻ>P����H���Ȭ�Z}Nd�{ ����         �G���jeĔ����Z�����р	��,��n�/2T^���p�R���G����Y���/��LPu!*�B�zYDf����N'        �>26e��htpd���:>��d�s��FGG_^O�u����jtAp�	���.��ґ(fΎ�ԅ�V������P}}���Y:(2T]|A         ���~���'�Z����&�%K�l�jժE���%�}������T]pV42��Q�#�qd�3��)EQ|$rt��Q]yY         �']�(ҭ��b�Gn��8��j��q.ѪU��UO���~�?��S����ֈ�w��ctt�CCC�L �&M��z�#24^��*        �>TUQ��h>�%��G���Z�Yvɦw����]Oo��rs�+�����U���F��/�M��ѧ���&�<���9���S        ���Ό�s_�hDn��xw��:exx��D}]v���#C��gi�� �? ���}q��(������Ϝ9�k[Y}=6����#�BT-�t��         ��mˢ�l4O�mS�gRJs�9le###/��C"G�&�?�4��p �b�._��3"Gu:~tt�����[��v���zzrd��wf         t�D�ܻ�J��j�^U/�����.������ґ�e�����T�{zdp��R���������K.yD=}$rU�jq;         �х�n_Ŏ;G��������CCC��z��Ǯ��j��F�������_F�G��b��###�͜9��[XJ��n��T/w�L�g}o�q"         Q�Q���h������:1�thQ)`��zzqd*����vp�p��*�3O��+^���Ч[��������v���z:8r�z��V        ���==sx��D���j��R��lA.|dQ'D��ӿ�i�& �	����4b�������s��9���ˀ-�����G���Έt��         ��n�����h�ב��(>2::z�����- ��h��'��#S���Q�����p�֮���ӣ��Eƞ��>�Q���.���i���zL�\�����^         ����F�E4��m�����ŋ������FGG�]OO��Ug� b����p�D����g??bp0r�R�@���1cƙ�I}��u��z���Xuɏ#-�%         ��-7G��h<�ɑ��N������hdd�)�wG��Ƣ<��`�p�D��;��h^4�vHd�Qo_�>`3h�Z�(�������        ����;��{�������3f�,X�`��(�^/������D�yG�i�oB�w�����լ��]�������g�VlB�����χ"s��H�]         듮�*����x���YJ��.\4k֬6�y��Mn6�߬�;E��Nt���`��:�=Ѥ�#E~|n4��{¤I�>W��E�6�E��[��7"�}'�(O�J         ܛ�['Gc������4��,x�xm�&�R*Z�։�2� ����"n�9�t��N@�w��AG18�{i��>2��olv.���r��\՚�{;        �Qƻ�/Z��#sn6��_v�e������ ���E�����Xt���`�p��Ҳ[�Ob4�������̙3?p?���S��"wU巿         ��{R4�03�ш����5k��t��C��w�5�����?�ӿE(�==�e��%�Tߛͧ��(���Fr�̙3���RJ�v���z���ՂG��v        ���~q]T���1+�UQO��;>�Rzy�N�Q�������L�k���7�MO�}3H���9�E�Yύ0X��,\��Y�f��Hu*Z�֧�����U�)_	        ���������^�����}��Z^/�p���'��N��/�g� b������DT~�k�x��#��=`�F�q����Ӈ��Z��^��od�9zDy~uS         �W�����h�94zAQ��9s�[6���R:�^N�^p��(��{��"ྙ����F�寉�}UUg�iN]��؀�:yo]��=b��|��        p��<)1u��EQ���j�6<<���y\}��S/w�љ{RĊ���C�}3*�>-�e��#z�.�s����!CCC�֡�a9����R�򕈻�        ��+-�#�S���*z��[�ֶ�����.�^�Y�r�����:��`�pߜ�2:_>!��C�C\U���v�Y3f̸$�)���.>^/�=$���(�9=         ���S�9�Ј��=䈑������EQ��{���WU�M��L���<�s�a6��,]qiT������!J)��n��zƌ�}�p�q���c:'�PW�N         <`�Nt���xۻ��E�v�=-���z]}ott�)UU��^N�R�.����`�p�ʓO���P��=�vo[���x�̙��ּy�&�Z�뛒F���DZ�        �M�j_�EQ<��1�m�Z�-Y���O��6�[�v�yUU�\/�D/��_6��J\OT�W7Ey�7����F��Zŷ������ヾ3����S_O�^�vM�'}&         6���2&}��#����(��_�z�ޭV�o���o�N�ٿ9�tt�lD��|�k�n�e��	�o!���F�O�b�ݣ�4�q�����+V�~Μ9��/ԟ���������у:sO���_        �&w��Q~�k�|�+�פ�f��ŋ-��8`i��Ν��g�}��?�7DJ��.��N	��-�Ӊ�玏��|,��s�R����y��{X��z�����՟�z�[�]�������        �ͥ<�;�x�S��s��AV�兣��/�Q��.����ƾ�RzV��������e�oAi�O�<��hrX���(�����󆇇/zN]|�v���z��zF/���|��        �fS�Q�pl|���fO�9\Uչ�V�?���?������׮]�mmޓ'5��~/��l9=�#Nd�7N��'F�ܓ��������� })�K�,ٮ�n�^� zX��oE���         �ܪ믉�S�q��Gus�G���'�z����;��V�%UU}�^N����շN�,�-m���|�1���v[�G��R�GFFf����c��٫��՟��V��j����a����        ���9�����(�[���ҋ����k��/�1c�eA�Z����3=�^�s�������V��ni�[A���9�E㙇E/+����&M:xdd�3g�\d�.@E}C�z�}<�6����Xt����        �Ŭ]���h��舁��uNO)-l�ZGΘ1��EQTAvFFFWO_�?����Ug�������;�D���b𱏏b�ݣ�=���.�һ�t����K/�t������3��s���k        `KK�]巾��2z\���Q�v��V����ÿ
��Rj������?X��=.�pm��81�:ܷ��>�:>bp0z\� }��؞_��2���]����u:���;GHW,���        ��R���(������R�+���CCC�+�"֢E���?���Ӣ��E�ӟ�T�l�[Q�����R����RJ��qi��:z�v8r�}�]L(�g�O=>[�,<=��]wF�3�t/�         �j�*����>��v��R�l����V������?&��s�vp~[Y���6;��W??����G�}+�v��?����Ot7�#�/_���a֬Y[����L�4���ߋ���"�;��H�/        ��-�vkt���xӿGyr=F�����Σ�̙�:��FGG�^U�'��c��T�F�<��`�p��R��},?x\�>$�������V�)�7Ϝ9�`��o
�S��˽��T�};��         �(�Fu���q�s��LI)}hڴi������/E��-��j�^�����e�gҭ���g����u	�O+��'���w,����3���3�t��5k�:蠃�
������ ]�<9�P�dqt��         �h:'>��;�GO�>�Ȣ(��n�_922�3g.
��V��C=u��6�o֮��1����`�p� ��WEu�g���o�>4�.H�<yr���'˲<��O|�b3}lUU����/��G�n��>Q�        0ᔝ;��1����i��CO+���j�N���ݳfͺ4�,/^�������;�S������t���� �>����>�����>�S]��xm��>j͚5��={��`����w�ߺ�^�lD�Jcc�9�Ñ�\         ֝wD�����HD�/����5��j�Z_+���x�U�&Q��S��ucccG���ǪsN�򂳃��/w���{��}�(��7��CRJ�L�4�]�����q��ÿ
�v�=���\��/�G3�\�I	��?        ��.]uetN�|���Ǻ]_�l6_�j�NO)5s�̋��etttת�^U/�\��E��~��(O�\0��O0���c�| �wt�>V��uOuO��.J_*����6�ܹs�{��s����b������Ɵ�         ����G��^јsh��n����(k�Z���W_}���~xܫ���G7��VU���� b٭Q����.���Dt۲�|�=1x��#�n�o��m6����R�.J'��N^��K.��/�������J��Q���         �M狟��]v��~C��'������{���j�T�O�9s�5�X�t�6˗/��(��~��^�"��ի���E�}Y0��OP���������h�kF��vS���җ���ʬY�F��-Y�d�U�V�u���z<=~{J�ߓ��::�$�rP        �PUF縏�7�-�g�V�#��xG��:;�t�I�������}�b�ߋ��{��˗/���G;�?~Oىα��zg"&*�	�����SW�~S�'v�Ǜ�ƛ���z��z|sƌ�ǎ��N<o޼��o��3��V�Z����]�N��Uc�x��i+        �l�Z���'�L�N;���Т([�j��I)}s�ԩߞ>}���.�^��/h��/��}���tBT�����W��a��-��~~�^�ף{
�M��|u]�N��u�:���=�jݣ��g�˿��3�q�`���<B        ���~���QL����zV�a�V��T7�^��H)�9<<|C���ZOs��Y�����ܫ�{s�:�`bp�@��#v�1�ܫ}���z�~�I�V������UU�Ѓ��w�}�D&.\���wR�<�{���l������H��.         zE���(��p4���(�ڮ�M)=����j-)��zy����EO|�o�L̛7o�iӆ�ev�7<���S�1�^���9Q�=)���sPUQ~��(��&3�l���C�ͼ�ؑX�|���8����럏���w�}���̙��ڿ�e�]�c��ٯ���cV����Op�t:�9�CQ-Y         ���|4�G����=�)
zLO)M��t�?��E1R���q�p���%��k��=]/�����5���뱍@��S]���|���Ϯ�����},���(���/���I�tE��&?mڴ�u!��~����?��.
�5��k��7e���/�6y��=��^��g�z޳�U�W��]�����QU���G�h$         zUվ$:�>:��_#��~���H)�"�|n�Z7����륿�v�իW_w�Aݵ�������:u�#��f7K8�-��6�}lw�?�lբ���������t:1v�c���1��D� <��+PeYv���Bu[�������b��^�Y�Wt�7���<��P���L�w�v�_�T�w�׻ԣ;O����?�	u��'Ղ        ��U_�m���W��J6�ݻ㏳~�'O�f
W��n���)�fo���빛��'W�;���
����}�_��;����a�U|����4:�}8��d����s�vm�}����D����f�Sw�~}}��?�� ��������        �/��ϊ��������{�#?����B����?��F��yp���5��ؑ�|�{�������F�<�sQ�yj         ����D'�x�k#��~W������"V�
�#���T�:o��?���P@ߪ��|���.8;         �Uu�iQ�^�׼%���WՕ�E����gL�=g�N����x�ј9;��|��Q-�0         �]y�y��N���MQ�O�hat��p��X�/�W�:��T��-�8���~���S��G�j]         �Vu񏢳zu��]���b����'ƛ�7�^P����11��D�i���U+�<�Q-Y         ���.֟x4��(&O	�u�ygD���^TA��{E���|�h��h����F@/J�/���/�uW         �V]>����x_�λ������W��C��ǔg�: xݿz�='������n         6l<su��b�_��b�}zI��c��~�[�{P����mY���Ql�C@/�&����U+        ���m�����|��8`f@O�{E��| ��\������.Hw�/�?4 g�9�E�K��e         pߤի�s���������t�/���F��MAop�a�7�ػ��G4?# ;U�ܓ����        ������'#��y4_�ڈR��c�S��N�;��wE�cGF��G��WD49H����GE��'        ��Q�wFT7^o��(v�9 )E��S������
z��{?�~����H7��׽=�m��Ȫ�^�㏊X~{         �i����λ��7���Lh�VF��D52?��}�Z�0�{�o�Q<b����{:�<�3��         l����9���<���|��LD�7F��F��A�p�3��7E�ȷG�寉�S�0a��+:�?�	+        �-�*����D��h��MQl�]�D1�0�˟�X�&�/�}(�^���Ƣ�x�#���5UKG���#�vk         �eU/��gW��k������t��(��SQ]���?	���j�X{���VTv���7������        ��d�����{�y�_G�ů�1e˫��4���an����;��$����|�c���:         � R���S��ْx�;�x�n[����if�� ]qi�ӛ���Gl6U�٧E��/E�Y         L,�ڟ�ػ����.��}aDSܔͧZ��(?w|��n���ҍ�����5�O;4�/�ǈ�S6���k����Q]�4         ��֮���_�Ծ$��~S{��I�]3~���}[�v���;�� ��Έ���h��_���p��-B�<9�3��        dd���o���6��{iĤIT�h$���T�e��1w�)�rst>vd4:���ܷP��Q-nEy�#���        @��2��+���c�U���qO�?��Ey�磺����pg��ϋrd~4���h�����#���(�Ղ        ����c������&�G��Q:�(�==�o~9b�ʀp�ޭY巿�E�G󅯈Ɓ�O�{ET��fTg�il,         �-�Kc�]o��3���4b��S-Z�I����_lw6Z��U���D㱏����9���
�_U����/D�yG         ���N�g���E�y/��3�h4~'��(O�\T���w���ˢ�o�����<��Q<t����ե#Q}��Q]M         �GV�5ޝ�:�h>�ј�4A�>�n�9��}3��8�<�+w�n��Fպ�.FO��߾8��<,�/���t���H�]         ��t����'�����;�7f=)�(������w���gETe��%��Sv���QͿ �O}f4��EQ�K��ƃ��81�5K         �?{��������F H�9S�HI9
�P��v4����sv��U�r��7�/|c��|c������lm�(iG��H�9� �  "v���ѬF"����y�>5��U ����~�OUN���������Zynq����.����L��ߦ2>��ܹ5J)�����z%m�<�����e���K)�Nʿ����        ������?���<�����7=���yT[�K���T�y]��[J��[k�T�Sz���?����{�jp����}#���s�s:         �UU������&�����\/$Ӧ��U9�'�_�C�۶L^�n5wn��X�]�31�
�ݟ������tRl��r�?���Keh0         ����M���~��i���S��/R�=74��D�[�M�7����C��I��ۮr�`&�����s����)>��-u�\Neώ�^�]��_{B        �[fh0���Zн����R�n����I���Sz�夿/p'�s�\�X;���
�֤�ß���?L:����r�/�w�H��ߦr�7         p[UYwm���*̙����K���,X���x*[?���Vv2yC%p'	�sWT��(�?�)������s)>�l
k�&�B�C�����)��fʻ��~Y         �;�r��Z��o�)��7������'����R}����)�����}�ִw��;w��@J/���2w^�6?��}?��v���R޽=�ޮ���         �B5d���)M�rGG
o�e
���L���[�r�D����ۯ�r�'Pܩ�Sz�_k�z�H�Ϥ��{ך݋��\Iy�֔����'�B�         P�*��l� �ɕ�))>�)�j������*�R>�7�m[jE���z#�N}���Y;ndr�����6<���6ך޹��;؎Iy��ɵ-�=;kOH         А�FS��NmUs+�K�;�M�)�{x�pc�˗Rٷ+�m[jo�Ꙁ;u�22\����U*RX�*��7���;)���wbU*��>��=���Ykk���        @ө��=�RuUKtg�J��)>�p
�Ka鲤PHK��)ܿ;���R>~$�H�i,�0���ZC����vSa��\?���P�L^޳����J��8��'���         ��ʕ˩��zʓ�f�V?���R�e�%��if�KRٿ'�{R��ګ��r9Ш�ix�s=���^M�zô�),�7�{V$�V��jMRm}FS}�ɩ)�>Q{�Y������x         ����ʮ�)UW�z�-�%���lE
�L���v�`Q��NL��s&�c��>�����\�h&�4��C�f��䪺�U�=�.O&/��'�'o[\�^��}w��գR.�'�{S�t}د>�         ��ʥT�%����L�NqŽ��E��_�x��3��;�+���'��c��7雼<s�Z��R	4;wZC5H�{��jW?��j���y)t�H�gN�)̘��������))tt\����������i}b<�}X��>��88�^�\�U�|��˗R�x!)M         ���S޻k�]_�\[{
s�&�f����j��cư�/lkKa�k��2%i�L�pl4��ש�T�O�^��)�������+��a�B��Z��;TU[߫+         @K+M��w.���� w��;           uA�          �� �          @]p          �.�          P�          ��           �w           ꂀ;           uA�          �� �          @]p          �.�          P�          ��           �w           ꂀ;           uA�          �� �          @]p  �D�\�>#��gfdzwƦN�ؔ��M�^n�H�X���eU�\J��D
�r:�F�1:�α�td�Е�唡�    P*�ktZw��?��Ψ�?ǧte���6-���\l�ݿ}b�6-N^V矝�9��P��3u�J��}�v  �F!�  ԭ��)��`q.�[�+��gpμ�L뾥_�}|,ݗ/dƥ����͜��L�r)     w�ՙ�si��\��0��e`�ܔ::o���:X��θؗ����}�G�  �[�  @ݨ�����_�<�'���9I����Ott�6��+k��n�μ�ә�D�=�)#W    p+�vMKߒ��_�"����x����5��!�u~����B���/d^���?{2sϟM�T
  @=p  �j��o���,�/痭����R��5�U�}�b�۟%�f���     |�Ӻӻ����V�q��=�Le��ΞW[��>���D�;�E'�V[i"   w��;  pW͜�ӫ����26�+�lp֜x�|�{��{:����S�R(k4    n�XL�¥9�z]z���]�W���Z�{u���t�<�w��b_   �4w  ���_�<G�o̅�K�h��F����֔�ܻoG�ڝ���     T��;rr��[�HƦNO���R�W��sg�j����9  �;E�  ��*���{sd��\��(�`t��������iCV�Y[c�    ZS��3'�_��k�x��Z�UU�J�k�žܷgk�8�B   n/w  ඩ�{W���g�K3�nT~��_�h�ܕ{�}��ё     ��:#<���Z�}��3�h`��|��O2c}V��8�� ��H�  �-f���M��҂%iՍ���6֎^��,?�3�J%    @s�N�ήz0�{2�]S�
�s�O�$s8��>z+ݗ�  p�	� P7�S��h_��r*�O���ޑck����M�XL��蜒}�Ι{Ⱥ������R/�'�����v���
�����5��@�9[?/� �>)2��~]�C{���s�gO��c�ⴢ��佟��,?�;kvlI��X�Şr!�[o6�m9� �zRO��  hq����	C�kY{�n�=+Vg���2:�;���������ve���b������]�&���	 �;����'�����m����?[�$�C�lΉ5�bk��*�bN<�pz����m�fщé��sP  hp�  ��V��̞ǟ�ٕ��S��y�[~_}�����    И���<��Ϙ�M��䓧��+�;[�L��h   �w  �[�5��y14kn���i������;�d�m���)    �k8�z]�mz&�f�9�|u>�=/����t_�  �7%�  |cgV=���?�R��_���~��'rqޢ|��ӡ�    ��DGgvo�AzW�_nh���������w  ���B  ��r{{vm~.=+ׄ����Uy��lx�%-F    P��.ȶ��4#�g����֖}���y����S,�  �u�  _�D�l{�\\�$|3��3����:���R���    P_.,\�����6�9����L��o��v'Z  _��;  �vM���<s�o��ޑ�Ͼ���5�O    P�-[�O���Dηsq��Z�Ǧ7~�)W  �U�  _I�u���~��ݳ­Qikˎ'��ή,?�;    ��u澵ٽ�/R)í14kn��诳��_g���   |w  �KΙ��~���uM�X����?��)]�o��    �#뿛C�l����������t_�  ���  7Ukn��υ�o���Y��xV��    ��:y�w��o�����"�_�M�  �M	�  74�55[��vM�߁Oe���,>~(    ��ѳrM�}�����t����\��  \��;  p]�����Ќ��Ψ
����16�ygO    ��.,�';����l�;�vj�s���W�5�c�  �<w  ���b>��Ore��pgU�m�����k����    �W�.ȶg~�J[[��g������o�:�R)   �%�  |��MϦ��pw�::������Α�     ��X��l}���,����¥ٻ��Y��  �,w  ����\�ӫ
w������ԏ��_'�r    �[�R(d��gl��pw�^�.sϟ͒c  �)w  �O�Θ�=��E�ݓ�k˪=[    �G�mt�e�����y�\�_�  �*w  ���֖O��Q&�[W>�xf��fn��     ��ŅKr��M�~��;���?����'&   �  ����t�.u�X��'~�'_��t��    �fƻ�fǓ?J�P�ep�����T��  p  rq�ҜZ�.ԧ�i������w_	    �����Tm�F}:�f}�:�ygO  hm�  ����b�lz6)B��Yy?����    �z.-\��+��m�������]�&�  �.w  hq��>��YsB�۷���9���D    ���Rl˞M���L���o���  к� ���L�Α�Cc�>^��m��    �j��}$�J>��β�{3�ʥ   �I�  ZX�����ѵ�e�}�:4    ��F�w�����Qm�߿�lx�  Z��;  ������=���Rnoϑ�l��^    ps�ެ��_�2,ɜ�g  �w  hQG�5�3�ޟջ>J�w    ��j{�ٕ���tt���y�7  Z��;  ��+s�ѲИ�G�{豬��     �w���)��1�-Y�+�ff��   �E�  Z���lJ
�иN��PV�ޚ)�C    ��h״�^�`hlGڐ��~)  @kp �38kN��74�r[[�?�H��^    �?w�GSn�ht疭�ହ�|!  @��j  Z��uS���N޿>��ٚ���     �LtNɩ5�C(rt݆<�ޫ  Z��;  ���)]�]�:4�R{Gά�?+�
    p͙{���h�+�d�w�12  �5� @9�jm�mm�y�Z�N�    >��}kC�(������w  h�  �BN��i:�������y�|    ��]��0�s��R�m� @�p �10{^g�	ͧg�w    �ԳbMh>բ��Ys3��   �O�  ZD�ա9�,_�����B    �uUb��z&��;� �� @��]v_hN#ӻ30oaf��    ��+�edZwhN=����  h~�  �����Ь9�y�_�B�   ��ַxyh^C������uu0  @sp �зdEhn}K�g���    ��o��������=��  hn�  ��ʅ/�O��{Bs�<wa&:��}l��)U    �T�Bo<��Ʈ�]�[������
Cs  ��	� @���
�����&W,�ҼE����2nc   �U�����/J�`���..X������  ht�  ��J_Z��=+�]�B�`�M�6v    hT�BR��|뒒��0�5-��33u���3  ��	� @��������Bk�<���x    �1�UǠ7���<wah��/�i��I�  ��� ��~I)���y�5\���z�bc   ��4�%��+�-c`��ܬ��A�  ��� ���8���??{nh�]SkG�v�\����   hP7ip�:�6�5~i�G  �'�  ���h�fi.j%���fn���C   ��t�������YsB���R��   �N�  �ś�r��ŌN�Z���3r�흋�   hP�nR�1<}fh�����X��ɦ�  ��� ���U��]od?2}f*��V22}�?w�Ѽ    4��7	-�t�x&F�μG���ԁ�_�\5�~�  ��;  4���u�RȬ����ӻCk�i�ݛ    hL}7kp�f�j�op���K1 �F'�  M����)SCk��c~Ns    ��M�ƺ���r���9%  �� �	��$^���)]����`cgdr���   �AU�ˣ�d�uF\c�SBk��c~�l
  �@�  ����о틷���m�T�G�   Шʩ}r�uN�4m=�78��  h
�  �N� �\n�+�)��1�\   @�;U�_�ơd�r��  �Լ� �&p�RL)�}ns�\,��Rik���5   ���y�:㯊9h�)]�1��\'�A �)� @�$'�ɪ����[O�x���A�E    4�C7/;ɲ�\���H���   ���<  h�ʅ�*~�x^��Vs�G|`�ۢGs    �t���J2��J%���<�J>  �y� @��[)�ǟ��X.��r��|�[|    4�r���k��iWu&Vh)�r���+;�  ��Wx  �$v�
)u���(s�:C~�[��ŀ��E    4��bk��X���}�1��\��b	  MC�  ��p
9TI���X����:��N�E    4�O�S�P����V���w��}�1�  �4� ��l/�`���u����1:�g�O�鷱   @�8_)�l%Y�{u&6<}Fh��>�����  ���;  4�-�B�����?�w�����񹍝-e;    4�Km�w�-�0m9�-���{|�K  h*�  �D��E�ʅ�*^������j>��X��   @s��\ȿ���N'Y���>��b	  MG�  ���bV��u��2u���B�T4�   �\N�9])�µT�ggb���>�ho ��#�  M��R!�M{!m����@
�J*!�V1u�ʟ>�Ä�    ��ۥb���kES��R.���P�É���9(  4w  h2�*�|R.dc��b��)�C��Zô?6U7v�-��   �9��T�h/�B�-}��MJ�|���
��  �G�  ����l�,�>�tA���t_�P���T��   @��$�K�lj+gƥ��:>��V�YV�  �H�  ���r!=�kq�R���[�"4�)#W�12\�����   hr/�1�^��u�\�X״��������J��  ���;  4�jw�K�b��bI{Q�tc�@����    �پr!�+��.\+��_,��
f\��������  4#w  hRo����J)��{Ck�}��v���"    Z�K���ϝ����M�������ɕ��w�� @�p �&5Z�����d����N��mv_oN��Z��   @k�R)�o*���S��
�����D[�  4+w  hb/����r-�ܻB���*��so��Rѱ�    ��r%���b���I��rRT�����ɥJ!�jo ��&�  M�������|��TzW�ͫ�&�3���Z�2   ���A�����eօs�<qh^�zN�W��wu�  4/�  hr��(���Ǔ�C�w�d���v    ZOu&�m��gO
�7�J%�������v  hv�  ���&�?_�c��38{^hN��Ndg��    �i{���8u2yX�G��ԟ�<���� @�p ��~��M'�&�Mi����ù��    ���{����+��Oۉ#�H�  �w  h�?r4�?�)4�+��lE�   ��v�R���#)�,4���  �� �E�x9�.^Ha���\^;|,    @�ڑc���{�)]���K�  �w  h!�Ȇ�O��1�>�/�    Hz��r��/����c��  Z��;  ����э�Rl�R�Y��oc    >kׁ�����{�(ML�ȑ�  Z�T  �����;v4���?4����?jc    >�ؑ�ٰis:::B�;~�hFGG  �w  h1�v|�U�פP(�ƶ��ڛ    �S��ط'�~44�J��=�v  h-�  �b�\���ǏeŽ�B㚘�Ⱦݻ    |��]���C���.��N;�K/  h-^� @����,_y��v�����    ��������yp��иv���  �H�  Z���9s�T�Y�<4�R��=�v    ��ݻv����X,��s���\��  �z� �E��d��{�:r�@�    ���������������I  ��$�  -���ޜ8v4+�]���xvl�    �����qV��/����q;z$}��  hM�  ��>��~�޳,��1l��Q��^    �冇��s��|w��Bc��?  к� ��U��ݱ}k6>ns�\�p!��    ���߻;��Y�9s���c����  h]�  ����ٝU�m�ԻJ��-ｓJ�    �+��������~�B��ץ���   �M�  Z\����n~��/l�Ա�����     _߹ޞ9t0�� ԧj�GuV]V�  -O�  ȹ��Z+��u�C�ȶ��    ��>���,^�4ӧw��s`����  ��;  P���2��ɵ0ԏj[�;o�����     ����h��ګ����*�b1ԏ���lU�  ���;  PSR�፼�W����P������    �����g�֏�q��P�������T*  �J�  ���+W��;o���w��'�w��     �Ξ�;�`�,_�2�}ՙ���@   >%�  ��ǎf��=y�u���;o�    �֫���Λ��ӻ�ݳo���L  �� �/�x���1#�,[�ꑼo������    ��FGF���_ʏ_�E�L�3����  �y�  �������y��/Ԏ���)�Jy�՗s�B    ����ŋ����~��io����Ο���R�E  |�Wh  �uMLL�W�����̚='�~�͜w��F���    ���Ο��o���x����p�\��7^y9��  �w  ������������*ӧw�ۧR�d�{��ı�    �S'��w�ʓ�6�B!�>�W�敗~����   ܈�;  pSW��j��>��2uڴp�U���>ڒC�    ��:����lشY��6���_}�w  ���  _��ŋy�7���?}!3g�
�N�\·ￛ���    �{��ڙ���<��3)�������\	  ��p  ��j��K��U���O2����J�����9y�X    �����>::�g~�ô��T�
�}}�SBGF�  �Ux5  |e�##y�������{��o��I��/�\oo    ��q�䉼��okeS���7�s�L�|��  �W%�  |-��y㕗k��޷����]�r���s�ҥ     ������������~���f���Ё����;)��  �:� ����!��[o��w6?�T�;:�Ws������266    �~]�x1��տ�{O=�{�[�����|���ܿ/   ߄�;  ��9t0}����~�9s�+�J���ٷ{W    ��0>>���|=gN���'�N{����\�t1o��Z��   ߔW^  ��r������M����ዮ\���^-/�    h<ղ����y��g��9ዪ�F[�7��  �6� �o��N��不�l6?�T�N��r����vf��6u    ��]�t)/��yl�w��C�R,C280�����S'�  �Vp  n��Ǐ���l��x�<�6�B!��g�����߭mz����\�@Ŧ*P?@�{�oo�ɱ��,�;�ZdQs;z$�{��̙;/��Z|�g���|LL  �Vp  n����|��;9�6}�,\�8�dxx8�>�R;���J��  �Y7� hU}��巿���Z�&6m�ԩS�Jz{�f�{�(�   nw  ම�ߗ���,_�2�ytC�͟�f6:2�}{wg��]    ��*�J���ԉ�Y��;Y���tN��f�w�|v��6�w>  ��E�  ��N�8^[-�#�m���������޽ٷgW��    h-չ��m[�g�άy�����#�:mZ�ɹޞ�߯�  ��� �;�\oo^y�wY�hq���cY���
�4�����ݵ3����D    ��61>^;����}��{�ս�{FU�����ٵc{���  �Np  �j��k/���3ge����5u��4�r���'O�Ё�9s�Tm�    ೪����΁}{kEk\�e˖�P,��ȡ�9���+  ��� ���ʕ����پ��,^�$+Wݗ+�M�)�'�P����9~�hN?�ё�     |�ZaƩ��5���6���A��\�,�^�{�<q<ǎ��C�v  ��E�  ��*�r�����w�`��,�gy��h޼yw��hhh0=g��Z�{&�\���    �������V��c��{�t��,^�4ӦO����\���=}����;/�  �w  �nT7U�����'[?J{GG,X��fΜ��=�f̜�B�p˾fuc���s��������ɯ]�    �c�����ꪚ>�;-���2{���,���~�T�냃�t�B.^���s�r���L��  �	�  u����i�������=c�䚙���tuM�m�T[��L�j��8y����nЌM^������##����@�k�    �j��Б�;r�O�U�ӻ�3cƌZ���sЎ��tvt��S-���˥R*�׫'QVg�� }u�Y��V������}   ��;  �P�1�/]�-    �fT�WW��   �w           ꂀ;           uA�          �� �          @]p          �.�          P�          ��           �w           ꂀ;           uA�          �� �          @]p          �.�          P�          ��           �w           ꂀ;           uA����/��sn�tG��H[{.L��z�x�r��r���/������        |�.^ͅҝ����w����ԫ%��R�T�=?�ѕ5SD���ix��<�}#�w�kΘ1#�.��z�ک�LLL�{�v�	�       �/�����̜93+�o��gR.+����vw��F           ꂀ;           uA�          �� �          @]p          �.�          P�          ��           �w           ꂀ;           uA�          �� �          @]p          �.�          P�          ��           �w           ꂀ;           uA�          �� �       ����M��Y��gf�%�~MM��&4iR�=�@�K���V�P��Cp N\�p)N= = "!�ĥ�xS+�DD�hej*��E�����ή��zgwvfg�-U"��3�����#���3�l�����  @�;           �           D�          Aྏ\��x��d���v���/��Y�w����j�M�o���      �e�����Ǟ�q��T�.��O�8��z���¿���I�Y��;
��3h��~�7v�       �4��=y�=90����uju�E.�;           �           D�          A�          @�;           �           D�          A�>���~���+Q�۫�`0�c5�<��л��F�g�7�r��L055U�F      ��Kn�ݝ�['��W�Q�h����߯�Y���^}suc�Ǭ�2�������ig��N�b�}�?+���~���f       �ګKo�+�=_�����ƈ��ڎ�	��o�Z��uڪ�6�h�N��ɚ��.��;           ��㧟�F���fh��u�굡�[���s�2�����������g�N?����77�Օ�����muj7�g�]5�j�V{���e~
      ���h4���<��glll������3S���/��Hg����^]y{�> �vx����c����+��ZZ]z��_\��v��{�U�٬͍K�q�B�?�'�c�?ykq�K�.�ιsC������?�ёΘ��?����r��GF�g���u�̙��o��Ǟx�vW_�      @�F�����/^���������Fn�f�P%p����#�;Ο���g��o�Z�������}�          A�          @�;           �           D�          A�          @�;           �  �8ب���^%�<\�9]���~��*    �q��q��V�.��ů�XSׯU��u�jcP  A� @�����Y�zڙ���G�(���G����|    ��v�]W�/��{���5�κi�� "p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��  ~��++�7/�A�9v��*    �qо�^k�����뽵��Q  � p ����֋��N     �����U�Jv  ��n          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�'���;k~n���        �iq�]u���h4 ��	t����_�(�       �P7���_�:���O����]}��N�f�C�O7{�?��h�lw
 �������H����:�Wj7u��       	n��}O�����~���u�n@���Z��+#��f���;���:�'�	wa�+�~�ѹ�g�6���Fz����H3�W矿8�|������K       &�`0�k�������������H3��?��?����ﭣϜ�KoK�          @�;           �           D�          A�          @�;           �           D�          A�          @�;           �           D��#޼T�ok��0���l�      01�~�=9��:r�|���g�;<��}i��5�� ��      `�4vܓ�+;��&p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w�ޓ�3�0ݼ�g�f�վ^�><?]�A����8�5       �����Խ3��)�Mg�NO���`P�޹K�D�;c�7�}p�NnW���        d���������H��%p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w�ޫ�^����zf�Ѭ��ܗ�B�[����5�鞙V��j       ���O�W[Z�wX�ٮF{��gZuT�D��?�`H��ֵze�{[�<t�P�w�b�z�嗫���w~{�p}��\       |�g��j�s{��Ç׽��N/��R�����g����w��          A�          @�;           �           D�          A�          @�;           �           D�          A�          @�;           �           D�          A�          @�;           �           D�          A�          @�;           �           D�          A�          @�;           ���ֱ#����j�������o���|����'j�Mmuj����       �G�<~g�>1��䛝Z��{r`�l�u�V���t{������L�}�wp��>to����-�;0�����~�O_o�      J����'_o܁��9<�;|���=��          �w           "�          � p           ��          �w           "�          � p           ��}���Z�^{�������͑su�_ i�����`���7W���^�'�����.       �ko��^{�R%jmm�+#�N�Z' Й�vm�����o�]WBZ��}ꡚ��C�7~G'P��]kk�����Tog���#� ���~�VF�g��n�n����4       :�nn���uڑ:�n~�f��ikk����澆t_�O�>^�����z���aM�X4�/��/�ݗ���@��<Z�<�������0��~��|��w�S�3���ި�-�      ���h4�����n����o���Q�{�6��c���U�� ���O�#'z�Z�ꭩ�������j7:zOMO��N���}�=��_���o�\�t�Ν;7����l�z晑���o��q>��:��O=���\gΜz���>y�d��+K����      ���h4����q���ZZZz~nn�N�:5�����q����ԧ>5�������ٳCϷZ�zꩧj7���Z�����          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "��ٻ� �λ�㿻{��V/���Vb����$5I�	I6�	����$&��R��0�RZfh���a��?�:S:����B���e�L�X�]I�dYﲴ�7k��{��鞫(F�%�c�s���dV�͎�>��s��>�          $A�          @�           $A�          @�           $A�  ��Z�j���[z�ǂe��)W��V{Mp}�p1�؃��;f/K�;.W6�c�����)�����^�����P��pe�_�&��Q��1��9�qo�.K5W���n�u�e�X���V[�q��\^�gůw��kbs�r���0��1�x�n��5�����׵.��\ߍ\/]K���s]��n�j������e  ��;�  p�M��Ͽ���Y�_��{����z?��(Ͻ�����g/׷�?�4���/��c�?�x���������m/��1���ߋ���@pm�����?sc�rwL��o�7��ߏ���=涟����엂�;�̧c8�;�[�!b���چ3ۢ������l�����_�������?��7���?�����V�9����=f�}������;�;�g�Ʈ	ƿ�C1��_���w<b�Ċs���*Zs]����Z������c�>�H��������ÿ��=f˯5�}�o�68{&?��=�u��b�o�~p}�?����W  ��y�	          �$�          H��          �$�          H��          �$�          H��          �$�          H��          �$�          H��          �$�          H��          �$�          H��          �$�          H��          �$�          H��          �$�          H��          �$�h��q�=w        @�n�<9j�Zcc 4�����}���j        @���m�/� 4��          �$���K���[���,#��<\���w:�������:|8 RS�޿�������c�m��>���~��9��S�˟�      �-U�7�s�2��\.����/��O�֊~F��� HM�;��������w}�C+�Z'VB��p�a?R�*��W���I	HP�Y��V��hq��?����pe�       u6�"%7�:	0��Z�|���:�V�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�gd���➯�e�Y�?�&Z?{��sx�       ��gO����&�g0�w{A��i/,�-{ ���9      ���99@}M�/���"p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p��ֶ���M����p8�TM,�>�o�����A       ����I�t���1�Y���'Hb���o�{������Hփ��;        ���ܧu�»� ��	�  ��s'b����k��T��x��k��é�a�k�p>�Az����Ͼ�gpr.�� Z�����Oé̞��;��mpr6H�����9   ��   �T��c����3�� M��_��O=\[��NU�s�,Ŏ�Q�Jz:;�G��moo_�p�\��S-���9&����ڊ�{�T]Ol�_W��N�h������  �Z|   �M��.p�����̶ M����ҒU��eщ��u��uiɪ�o�gW�}����3�5b8�T���k럚�ޱ#A��k���y:��j�ir��<~O   ��;   7�ݿ���ѳ�u�4������۸)xs��]3A���(���u�hpuŴ׫�u�����Yh��j�ܦg���+�L������h�i�=4z~ڷ�\]g�\  ���  pSu���bl�-��[�$���5�����u���A���R�~ue��K;�tU����WgQa����ױ�(i��mq����:}��T�?�D�������   �� p  ��*��1��?����󤯊U�Wg�Opum�"����UT���cc������� ]�3�F���7xs�O|m��W-�`_�1  �j�  p�U�
ܯ�����p_S!�N^w��(�h�{{�͌�i�6�?�C�c��wW���{Aڪ�F�ojx~~t�i_���	���c  ��|�  �M'~��ޱ#1���V켸�skb"x�o��@�.������d��z��J���3��
+7~��+u.��@�įW�?57��#m�W��Ԍm�\��    �U$p  �+�슲�Dk��rv����׋���
.�;�?g�髂����� ��ۃ�U��g~ ��i��u�����_U�B�z�ر=�?���r�=]�ȡ   ��"p  �+���윎�~$����>��J�~�δ1\ծ������]��H_g���M��Q�	��;z8��b��;��9�F����o�5q}T�u��F�Ye   �Z�   ��j�`���:SB���B�[�����:���-����V+x��F�1�����W�}�;���w�Nʡ��{�'�וEŞ�A=���ܢ����8M�MYh  �j�  �*|�|���S�?��(f�F�V��ǃ�����v6z�Ě�^'橗��������YhT/�.���uvn�D@=���RuL�����/�D��Fkb"x�E�   �6�;   ��:ʾ����^\$H�������9&����j'����>��R�~�b�TP���7(�iub��+Y,W/��+u��-�,�z({�(���>\4��}eo   �j�  �*��bt�����"1O�Ta���uv���j��M��BpQ���蟚�ü��atf,Ҩ�j�����۴9�Ȏ��2��w�ĺo_b�Q�T�u��U>���   `5	�  X5����׉y�
+7=�|pQ���_�I��;|0gN������/�bij��&?�� ����k&��*�����D�T��-?|�1  @
�   ��Q��^W>��\�n���?�j�g�G��-�࿖�2��m1��ǃ�;�R?U,p��:�ixa!��QTʢ�A�\ڱ�5>8�   �4�  X5��p8���+f^G��'��P��7�n����:�O�4��x*��Uu���"c��:S��K
c����F����q;/�D���ri���{�MW���   ��;M   �����Q�����i�U�X�Q�~q�eP?�� p�����z4�A��,RO�=��,:�Z�.����Z.^�޾�1��Mי��Su?#p_���5e�   ���   ������!橳*�������3�뫚��Y��=1��c��������\P?e�Ů�X���F���h'p�i�]O�XQ=w_�r4]�  �D�  XUU ����ɪ#���^W���\_���cp�L����h�B�_[��]ӱ��E�u���:����^����n�s?Mv���z�l�z�D�V+��"   R!p  `Uu�^��sx���^�1w��;����F;(SSՎ�;�b��M&橷��k|�n�Q����(Rw���O���6�����-�ES��A;�   �@�  ����F�x���Me�������|��h����+���np�><?����w;Q��F���^��k��D��6|�l��5��M微��yhc���+{G��   ��;   ��
�O<M%橿j��&��p��v]m�Q<�U���~D��oyN��(B}]:e��>M%��j�Q����F�W��O}_4��   �����  ��*�����}tx�Qk�S����ݻ;�blrC4�1\eQD�gg�}�C�DŔ1��*�nj�~�T'�Z0��s��T�Q�l�駡.  ��;   ��������ށ}1�?c�6G���Q�	�����<�{��h"1O�籩�{���rR�����?M�����L5�D���18s:��ޱ#1�=�w�MT�
   H��  �U�;�?g����n���kp&����L���?MS��e�	�
+��W;w���zM���W������j�v��V+��B�<�O�:ډ�}�h�u���l��&���`�O�   �B�  �꫎s�1����h1O>��72p���(fuvn�D@�����0bl,��:	�:I���v6z�Ě���q
A>���OE�Ӯ�sQ��51pw_  @j�   $�
��;<M
AZ6�z����a1�5�Czw싉�M�Ͱ�,t�om\�~)�'�5��vp�GS��a   RӬO�   HVwm�vxN��wFYt��v]4�p��4rQE{v���?Mұ�jV�(�q�� -+����s�$�y�,�<4�npr6�Ǐy��9���bl��h�   �F�  @�{^�ᅅ��MQ� 9+e�Ů�X���FS����:M�I�{9�Gw��|�N���/F��-��Ig�h���;�?g����n��g�,�3�-&?����E�   H��  �$\��=�h4��'?U�Ҥ�]̓��9���W�)F��/�(��5/]:y�|�f�?{<�wn����33eE�h���F٩�����   �H�  @2��Q���';M������cc��ic87�Ss�;v$ּ�[�	:;�/�G���T�w����	�EFݽ���T�M
�-��O�NG)\  � �;   �hR��<uwn�F�o�[.;�egx~>���ă�&(��,�/6&p/D�Y�^_74$p�t�D^�47����䥻gW�E'Zk�Et�\O   ��f|�
  @-|s�v���v��ӥ]H׾������185�
\��e;���T��?�t4����Ӥ�%,��Su=<��c�"wť�o�J��Eg�t���#�;�4   HU��    �QEt��u�(r'��W�ce�BT��*����"wU�38{&�OS^c�]��;��������1~�m�;�>�4��vMǺ�?�3��U��5!p�H  �T	�  HJ���F�"[�n����#�;1O��������9�SsѾ���Yw�K��C��7N����c��j��b�L��j�Q�b�E��j�))��   H��  ��T����W"g� ��(�(ˈV+r��d�
�{ǎĚw~K���[����Yu����'rܻ{vEYt�<5!��ty*vl-�i��D�,�    Uw   ������"W� ����;t ���@�jp�d�
�U�S��Ŵ�'gU��!��]���&�2љ����Ɋ]�Q�z�Z�o�ٹ=���Tv���X��D��EFi   �*�;   I������\u�����Y�v��_5Om��ӑ���cџ=�+��ڲ�xb�����16�!rU8� k����=;c��=rU���^���wvX�  @��   $��Y�N�U�����\���}W]c8�W��͍m�9�Ͻ����k:�=����p��� o�5q΁��F�����_��ȕE   �L�  @rFq��9�� /��
�֙z!rV�y��?z(���}��#c8�`Ů�X��wD����A��k�\�ށ}1�?�m�K��X���"�� o�Ee�jE�,�    ew   ���κ� o���l�g�G��-�������9�_13�O?9�ح��88����o#9�U�S��&�Lo-8j��Gn�{w���B���kg�wp����ȍE   �N�  @r'g��X���3r��樞��OEn��
��_5�7d��B�����v�TgF���)�����>��L�&n�����n����ȍ�������]1\�   ����   Վ�3����2�;b���u����W윎�ۍ��D�Z8�=�,�(�쌵�(rS�l��X���1p︯k��n���En,4   uw   �T���\���͒k0 po��+{G;��m�9�5G��E���?���Igjk����g������l�յ���Rd�,��14Cg��Q�  @��   $)ǈ����;�?gN����E..Ţ4C9D�c{���qp�T�Vv��E�RT�~��"'�1�(�"��\�Χ�9���ѾsKd�Z��$   'p   I�����;� o�o��8���"���(�ݠ9��F9��"�޾�As����[��b��&�Lo-8j��G.:�p�N������~�=��u�S����x*r�=�/��^   H��  �4�v{1&?�ݑG�7O��nV����qr�)�ZtR�As�Ξ�ޑCAs��G��+����D.\7O���Ɯwc�q��|CF���r   ԁ�  �dU"g�;��r�<��}if�kkb"rPÍ3\8��/�Ļ�9�l�:���Y���M�>8s*�G-�h�j�������E!n��v�w_  @�  HV'�p�{�G�7Pw��^X���Qw��Ů�Y�^/��fb�C�ti�TL��M�n�F3Ua��g�9U6S�щ0�������wpΜ��[o�tf���   _w   ��۷'�8���4O9�Gw�t�{�cQw�����A�T��f���Q��#h�jaæg��X��L݌�p;_7S���������L�4Pu"ێ����cQw�W��`�D   @��   $k�c��������[esU�}������1|K�_�}Yt����5x�p>z����jn�����;��U�@1�ؓQw�u�ՙ~1���<  @]�  Hڙ���8�_�S����7h��?���;�?ꮻgW�LU3�O�A�]�[%�48}2f��ߋV��o��ύ��L'헣}�ۣ�z�_����~5��kQw�mvpo����If�G�u-�  �&���>   �뾼{�u5�������������.��?��b��(�w����U�`�51   �<w           � p           	w           � p           	w           � p           	w           � p           	w           � p���Ρ3����ԟ9�acl���H���{b���z~�������       ���}�t��ܮgr��r�=���_��p����-���MZ'�!p��:e������gll,R�Y�}�o���\��7       \n5Z�5�v�T�>�Z'XU}�$F�          @�           $A�          @�           $A�          @�           $A�          @�           $A�          @�           $A�          @�           $A�          @�           $A�          @�           $A�          @�           $A�          @�           $A�          @�           $A������X�����V�����m\�Q�9�׏��       \���꫷i2.ly{��X����I��������y4ꬽ����x�m���ל���      �eY����N>�sr����=��|_{v^��0�;           I�          ��;           I�          ��;           I�          ��;           I�          ��{�>{>fg�F�ƻ�X��]�c.�����~l]�|�pj>f����wĚ5�       ����s1w�\���X���N�a �ٿ����Ҽ<�H���w�#��Z����̙�ػ�X�h�ߏ�+�]��9�ĺ������x-����{��      ���gΧ�:u{qJ�d�`�_QP�9=�����.�{���fb"ZK�{+���/����b�M+��o�K���HK{b��|6���/'7Ě5+���[3������v����n~       k�򟱢�)Z+o����ii�]Y�4�:��7�O��/�e�Fevv6^y�e�ڥI�{�����g��矏�ݻ %��S?�=�ܲ���W_��[�.������G������q���       �mll<~�g~�-�'N�����/��ׯ_���߽�����>���|�g.�y�e��#Gb۶m������x�G��ک}q��L��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;  ���1q�Pp}g� A�IcxY�� 5c�����A\R49�j����6X��sA�֟-����*·��4���b�1�,�V+Aj�J��˵�t��	��2������B   ��	�  �`���M�Xp}��Ǆ	Z39���R���G?H��x�^��3����Їc얷���'j���u���������6��4?>�gb�:cx���_�􌍵��e:wh��  ��           $A�          @�           $A�          @�           $A�          @�           $A�          @�           $A�          @�           $A�          @�           $A�          @�  �� e$m"      ��>�D/��n  !p h�ώ      ��ɶϑ  H��          �$�          H��          �$�          H��          �$�          H��          �$�          H��          �$�          H��          �$�          H��          �$�          H��          �$�          H��          �$�          H��          �$�          H��          �$�          H��          �$�          H��          �$�          H��          �$�       �{wd�u���z��{�0�	b#� . E��"$AR H��%ي#Q����Uv�8��8��D��8�����N9��6+.�Jd;^d
K/ӳc0+0����[��G�pt�x�s����JB7�������w�   	w           � p           	w           � p           	w           � p           	���+�         e�Z����  �A�^Cwݱ~�Uj4         Io������	 �C�          @�5wp߳шk7���j��K�����h��o-�5�@r��D���K����+��-�%-�ï�v�t       @��k���h���%�X���[��G 9���:�k��><�"n�e�S٩^�sx�8�C�^sgN��1��~~�ӌ�w���8#����:�;�������gY�q���       ��8}b�5�e�N���N��������۶������e���'�J�          @�           $A�          @�           $A�          @�           $A�          @�           $A�          @�           $A����3͸n��� u4zz�����"       `)FO�����NU�u9��K���������� �zV<�      @mxNP]�^9<��kE�          @�           $A�          @�           $A�          @�           $A�          @�           $A�          @�           $A�          @�           $A�          @�           $A�          @�           $A�          @�           $A�          @�           $A�          @�           $A�          @�T�_�eM���_��l5��șÑ������迾��|w�       ��/7���׹uj6��Xʭ���E#����N$F�N��;��:�{��Qom        H��Z��� � ,           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;��;�N��v�u}���x̯�!R5q�@�{��|ẕ�ت�        8���W:�oדz�4y��h����<}��x��рTܩ��ͷbs�������hܽz"R��w�N�������        xտ�o�����z֬��n���KE�z�������;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�  �����;s:��~Q,�����9�^��wEz�ǏF�ԉ�����'�ij���#n����+��4u�_���?��΁W�4u�-I�}��$u�-U�ؑ =�ӧ�{�H4�ǃ�+��   ��  �Ҝ}!�_=\���[Az���14�bq�o�9�ӧ���� =�ſM���@py���4[6��Co.������4�tpy��51ij�<C�u���cktO���zq[D�C������h���)��w��<\^��  ��<�  �!�-��jEcl,��BT��~ьbkV�%����T��� M�����PN���z1HSs�X�ԗ��s=����j)��:ij���cGc���K+D��*�*�D���|opi�-���0����+p��~���&�  �0�;  �),�fc��.��Ri+c+�������!��S��֜y�$�������{�X�����ڹ=z�N����Ҋ��D����Ϫ�}(�4�����l$p�<��f��k+�fm   p>�;  �E�����[�o��U>D^�����A{��}^�Ii�9��{c��ۃ���~��ſM����xpq�{�{�`��rR����\s����ks��57�N;#���5��   .$p  ��A\�-��W�+��zCC��l������ٷ;Fn�3�81O��s������+Wv�_ZaG��V'����=�=r(HW��\��scl,�����@��{G��[c��7W�&  �(�;  �E�H�U�ÆMc���N��֮c���x5�������EŖ�A��8x��Oל�Ze�Z���j���WF���31�jup!��7���x�7��G��^���'��������v���   .���Hh(�c���6��.�P79�Ç��_�H�G��T{Ƕ��M����P>D�_\a�F%��O~6�P�i&��	������Z/n�Vl����������WNZn-~f�x����hT�5������P͙�c��_.��qv"@�yNP]��\k�>�8ϙ;��K�z_T��B3��?��9u������D�������w '�Cd��E��2��j�O�UC1��t)V����]�9r(Fn\���n9���iGsn&V>���|��Ǣ�ow���O�~q�����;����"��P�彤h4��hP>'�5v≨��S����='���o��}WT���Sq���� Mw  �K(������?���E[�W� ��[���_����=�=r(����TG�q*F����|���(W��_�9���X��&������ٿ'H_y-Q�a�������'��w�x�w�ѻ�	��4�  ���   �P�<g���(�.U������p[���ۢw�TPe���^U�z�2I�2���_`p�E%�.�0I�2;����~Ps�y�*zgN�0c�=���v���x�'p�!vH  �,w�   .�{�X����;�^e��j)W�����*��R����km���3A58�\��nG�i6��b�t�;�h����ޮ�~QD�u.�zk�*�p������sWKy/i��/�*�9v�   .N�  p�S���l^-e1��'�WYq�Z�+*�N*�ܮC��Y�ͳ�o��j�7k���ppֹՔ����O�~����2������W�a�Z�S��X  ���   �Q>����烳:��x�a/Tl�
���Ҏ�:C�k���<���v������|op�c�z�3�	�@y-Q����2"\��׃�ʉW�5�a'��VK����x9Fn��e�  ��	�  .�jJ�������݃-����!�����#��
���9;��x_���7I���(M��*��3����g	M�g0�f�"������I�=v$:�v��mw�����c]�����观��S�   �&p  ��r����Wbd�-�ե*�������	iUU,���ڻv&�P-�1�Y��7N�2�� ����S�X�ziG��s_�����s1!phN?;�R-�9��Y�V�  ���   ����G>����RUU>D��e��j21�UMAZ%�f��jEcl,���AhJ��N����b��{����v�7�S^O��rmUM�կ�s��w�r�e^5��  �e	�k�Y�b~�)iq���m1;Vh t��[���t�G���\�fUY��<����w[�W���Uv!��b����h�����USĶ���<u�t��2��G�6���B�V-���Qw����ֹ�z�e^e�[M�d�r7���o��3�X�f���4�b����:u�N@�N,�u:��N�t����h4���kh��#1�yO�h�ӉM���3ǻ� H��|;�K��#q�ߦ�`��x[�Z9 ����t`���ZI�V����:�>��{�
�t+`�x��;�I�U��w�p��!��g~2��$��jN9���M3��WTO9��:���G��Μ�q��~?��b��>ugw��۳�plޚ�ݡV;��:��z����3�8�Yz���s(N&�:}�Ï���h��;  �kh�z1z'O�К�QgV���~�;YV��=Qg��j+Wi�{�^M����T�k��Qw��TPMB���\]�#���護G�9��m�cQg�Ʃ��j*'��=p�:9X�  �����O~����ۚ�ĉ�q���%���H���²^���_�ûv@J��W��O~b���ر����^���ka��14Ԉ�S/ǉ#�����V��ǣ΄�V��u��PY&(�+��qP]e�]�X��ᨫξ��9r(���$�/�����z�(6N�U�</pwMUi��1M�w�p�������zv(�RCCC�/��k�Ǐ��C��~�b|l,����,�5��7~)��9 R���6>��/��_9|8��^z��X<����{�Z�n��h4q���8ytg��{�ݲ����Z9�O�^������Mox�^cdŊ H�����u>k�x9��/}%��ܽ��;�Zj'�W���h�x����Uך��~������rW[���h��c�>u՜�YTue�5��OE]�^��ӧ���2ꪼ�jm�	�k�g��mŵ�o����Z�:�0��J��9����8q�̒��ʕ�n���� 5��oY���9:c�>!hxx���Ë�cA>��D  `���F��+ؗ1�U��D�Պ��X�Q��^�TW9Ѧ�!�x(��E9(W�u�n���+��:��{�j��d�ֶ-����j/�iz�N��䚨�~���Au������X��QWM�4   �D�  ����q���UQGM�KU^��l��<u�,�4[�W^1�lm�މ����RPme�=��3QW���{�e�F�u��ΑC1r㺨��1\}�c������G��Nܦ��	su��ͅ�d#   ^��  `	�n�>+{gԑ-��PF޵��<Y(��5O5�h0I������ʠ��oPm�D�1|�QG͙��+6N���?u�4�(�ئ���c8u����i   �M�  �DeP�����("����F�B��I��hD����=z8:���ȭwDݴ���x.ʕ��������=r(���pu����q*��:�m��'�0X��ݎ��hԍq  ��	�  ���۹�6�F�(��+f����Fcx8�<~��sA��N�<z��n�i��9�\L�0po�&e�U���|���޵s���ںiq�ӌ�����r,[�M��o���ec�?�Hԍq  ��	�  ��Y�v��,���5���T>zgNG��m1v߃Q'��p��.Y(#ٺ�hm��+'>�٨qp>�f5i�(��{�O���dԉ�F��wڋc��X���Q'�޻�\��n�{��m��   KS�*  �*��@7��Ŋ��u"��K9a�n��c8/���1��/D��榣�5I#E'��1Z�AZ۷Fo�L�ZuR�����*Лfb�;�uRƤ���-p7��K1�t�3Q'�v_   `i�   �P���
�{�(6�<'�UW?��1O^��8��1����=�=r(�o\u1�f�<�n���X��Qݣ��]�Q~��-p/��Y���a1�8'�٩�����pԅc  `y�   �P�����G]�l����e���d�t���Wbd�-QV��Oy.^���E]8��SZu
ܛS��ܜ]9�>�]?���?�v4FF�.��SA>�{M��c���.\  ,��  `�s+�Ex����#�ٻ+Fn�+꠵}k���y)W ��OD-t:Ql��R~��)p�Ze~�v��tM��bn&��V4�Ƣ�N�z����o�:h���#������j��zќ}!   X:�;  �2�+L�^�c��u`�<�+O�$pw�i��uM�b���� /�	s5�/�(��y)6�D�ݎ�h=V��{�.�㷵xn�����T�u���婜@6��3Q�vD���   `��   �T���	�gm���!��O|.�)H�Rs�>�KS������IsC������`'�R�|=������]�^-�4�S~��%p�ӵS��c�5O5���.Ou�,L9  ,��  `��2��ӑ�ξݶ �TmV!����x�ڻvF�������]!H�S��٩X����Yq5_�8��{�^�w�A~�~��L�w�x�w��g}/�y�ш�5]Od�{�pt�[�ܙh  �|w  �e��
S�i+�媽ot��u�#ge��=v4���'/���F־A��2��C�n��|��/��ȝ�F�:7y�1<9��eMv�M^�������yy_����s1Q���p�  `��   �T>\-��[o��Y!-oep��C��Y!-o�1�{��ڹ=z�Ny��D�~��M�A��3/�$���ZW�ӧ���Y;v��3��V�yr�ݛ�[�����g#g�}{�k�D  �e�  \�b�����C䬕����[!-ou8G����g�_4�1�"r�ں9z�g�<���v���\�����x.�W�Y�{�^�e��L~��3��V�1Oa\  pE�   W`���ǟ�\u��RO��	X�/o�m[��ЪՑ+�p�:�(6�Ŋ�=���F�qpƁ{17�V+�W�Y;��3����|��o����"w&i������7��\�  \�;  ��=nM�?�]k���:C�k"G�C�s�� _�n'Z�fc����j:g�9�lց��4�7��?���U�%o����L�k0�9�J���%rT�Y[�^�V^3����"WM��   WD�  p:{wV9�t�)+��@���b��	��9�|������[����LV���T�׌� -{ݣ���O��zG��1\�
�#���Q�SH�zA��{P��ϙ}�  ���  \�2�y�G"GS�:(W]�7p��A��V��[Y�1��m�����=~,�[�qp�ۍb�l���q��<��q]����Lw�z���c  �����  �uR���:���w�T�_��/�1O-4�#:����nq	�꡷0��b��7En�Q����[���9�lL|�3���k�b�� 9��ִ�\-���z�N���ȍq  �����  ��$ׇTM[��Fk���h������[�w��E[�b���Fn�SB��(�'���D��r��������|U�@P^듿s��_w}�<~��1+5��Es��,w��3  ���  \�����:MLFN�<��ﴣ97+}G�0I�VʝrܻGGg���ʰr�*r#橏\��I�Q~�v����EN�5��G�q*V����b��wk��{Q��wn   ���  �
���(�c�;�9)��RL?�]�.橗2�X���#'��z)f��i�hD.:^���W�z�2.c�Y��:iμ�?�������(���M��j%�{Q�٩��C   ���  �*�bN�{�(��:�G��@S�S+�s+�E.�Q/��Ǣ�ww��qW��1\?�5��~,rQ�'�ǎ�Q���
���ʰ��hN?�)\O�Jk���h���\�h  pu�   W!��U�9[��M��{�ӎ��h�| ^l���`���v��=�E.��U�Mp��v!��A�Q�.����>{[;�����ֶ-ћ?C�VG�1jsn&���o^l���<��3  ���  \���[�Պ��X�@�S?��� ��Ñ��F�4�ha�l�A��s{P/�N�z*r��*�\^nqp�D��i��m�<4190���~��2~��"��r�J�4���&p/���  pU�   W��nG�y6V���ȁ����3�e��y�<��<���Asv*��nP/͌�]�ǣ�gWP/�V��%n����^o����w�7r���r<�M�n��Z��T�if�  p��   W�\�2���܊o�� x�k���I���(�)fiu�yy_t���7G���~?��^o0Agջ,��{���=I���l�����i��I�TN4�w����s  \=�;  �UjN?k**��mK����3x���EE���Q_�#���o��z{T]s�$��jξ�?��:�ꫜ��C��<\_���:��Dw�ڈ�i�M/ ����?�����8�O����[c��7G�م   ��U�  ��^�������Qu��z�:������Qe����[����o�z�ܼ!���ecPO'���E���E���ѿ
������<UW8�Vk�l�΁��z�E���C�'���Es���DPOǾ�?��wGՕ�W  �:w  ��T�����Pe�����*[�޿	��ֶ̓/��2�uML���m�0�w���gU֜zv�   w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w �č޴>�n�%�׋ց��}�HP}cn���bh�ꨃ��|tO��林�W����h�~�-1z����9�];��{g���u�/��7��7.(���/�3��)�W^�:�x�#1<��?��s�X��������X��{cd�u�9q<vl�      ��&p HP��������|-V���y����^��oš���G���ch���?���Xq��QK�~���'���������ߋ\���%n��/�M�z*�WO�+����;q���⹫�14�>����.&~��OIsϮ����o}3z�7��o{�?���������ּ��q�/���?��������k����c�o��q�       ��; @b�o�#��k�zࡋ��re�7��o��/~%�|�g�}�`���o�/��ߍw���h&m�_e�{f�t�������G��}Ϗ����7cd����V���������_�-��s�>r(rW��O�k��c���tǟ��c�矉���1�}K�<�������*)c����_L��Կ_�����'�{��oB�r�      ��&p H�������Obl�ͯ����<��?��g>�G�t�a����?���η��o��G���;��/G��Ѩ�2 }�����^��c�����W>S����ܱ����IIU0~�����3�+O������l�韋W������J�o���1�}�K���������_      �kM� ��r�����-)n?gŝw�}�1�3?�i�w��-n7|�1��#���g�f�*Fo�)����EܾL��S��W����+����/�ze��s����o�ԓ?�f3X�r����D��w�
6|�O/-n������S��Q�       ג�  �>��WC�/&�  ��IDAT}�}q�>���Aznz�����6vˆx���?c��Ӄ��
n���� 
f�n��S��o�N�&4,ժ{�ӫh�w�-?�s��o��`yn�S?_���<g���_�����W�R���OD�       ׊�  �>��U���S��nxb2���o�Ư>g6o�����6W�ш���|������~h(������7��w��[����G�n�ēW<1g�}��J��      T��  CC1���W��k��� Mo{{�<Ók���VL���9y"R5~��1zÍ���|���{)�������� :��_�6|�OǶ��#ek���������!p      �)�; @F��!�W~iv����N�������[w��w��_����"U�7�\���E�r86FoZ'p�7~�3�����u�H���[���G��       ג�  �����bj�{Z����W;#���������v�z��G��F�]����U�����w�q����ߗݦi�۴�RF��AD��M�  ���Be��
��R���" �(��ޅ�4m�Wv�������5����|<H�y���os������o��4r]ACwH�;��y�#[��Y}YY       t&w  �,mm�P37�F�: ���όW�;8 r�Ѓ����]��W       �p �N���ǣ��G�o���txu4̝ ����_��~Q{׭      @�� �ͻ��z�aA$1�3{F͔� WT}b�������        =�  ЉV��j̻sJ;���c*��N��)����Œ'       �#�  �l�/����D�v	��k܆�k��<^�      �� ���57�k'#�87��:1
JJ��+>" rM���o���       �'����C�K�w"  t������ļ;�Ġ��}��6J�VEa���w��zE�!�OEAYY���G>I>'�Ή\�((��#����n~��^�Q���Q��vL�}�9    @Ǎ9$���DA  =��{T\\�z  ��k����z��w�56����z$����3��Mu⟻o����_l��k��5�[_�ŏ�>�[??#
JK��5x�b�?��ŋ    ��)))J=v��Cʹ�[�x暟�:�ƕѧ����
���'��Fb� �6mo�������>��e�/�+�̌�T�J  ɻO=��s��    @�ڢ�O�Ҹ"��ݗ$V��uZ�* �δ7��:5��u*(h��sx���A�p���j���m���m���h�|bz����cEӳ����#��sۥ��s  �mءG�ܛ~mMM    @&�b��v�V��:/_M���:-�u�O�ÿ��������q��<�;�/�;?���   :Iɐa1h�/Ƃ_�"       �h�    ����      �I�   ����$�~r�X���      �'�   �ɪ�� �      ��    ����?e��D���      �p   �d���v��1�G       L�   �9�И5��hY�,       x�    ]���O�����eR       ���   �H��Ǽ�n����       ��   ڡ�fN�V�ȨG鈑��ӟ�E?       ���{>ii�����e�9�� U�Ғ���� ��j�#O?7E���:b��;    ��%����E��� U�y���&��G�̞���  ���1�9  �5ί����?�OF}�n�M�������    ����Q��� 9��۳S�,�    �Ts�ܓ�vl����      ��&�   �N+^z>�?�����'3��ϼ��8�&       �w   �4�L��q�=QTC�|D̺��       �?�   Ұ�w�GC͜(��Q�a�s��*Z�W       �"�   ����樽��u���)�����/j�-       �w   �4���֨>��(��;�>UGL�ڻo�hk       �   �ּli,��z�Q�����o��b�_�       �   t��[&��/QP�Q��#'�      ��    P?}Z,~��Ӯ����]���q�zڛ      ��	�   tм��3�G"UGo_xn       �t�   ݠ����]����=ݒ��1V��J��`|F}���y��y��       ���  �AAIITn�c �o��7Ǻ߽4�ee1���cΤ�      �'p   ���_����F��Q�a�so�6ښ�      ��p   �@k}}��uk�8ጌ��?�����/      ��p   �м�o��ǜ����?�Dw      �Gp   �P��y��w��A{�Q��7��-����>       =��;   �Z0���2�'U5A�      ��   ւ�/��
�''�gb��{D���Q?kF       �4�   ��� ��f�����v��1��o      @O#�  ��K��Z���0{f�V�ʨϐ�Y/���      �'p  ��Y3���!
JK�]m--1��)1��2�SX�'�|��Qs�      Г�  t@��U��Ϗŀ]? ����o��SΎ�����:rB̻��Th      ��p  ��W_v�LDAA ��y��Xp�]1�У3�SZ=*��9�,�Ã      �S������[��t�6
�n���V��+
�Z�>�J���+_{9fM�<F�vN �_5S'ǰ������ww    ���Oe�X�ҵ�����X��Y���D[[ �g]Y'��g$9o�~��i�M��J{ �{
�zE���E�[E�:c�dȰ((���:CaEE�=ښ�#[��鏣�wy?���)()��M6��6�ґ����O�Q�������Q�DQf�q��4�6j���^�e�>-˗�W?��X��G��Ι}/�n�m���f���    ��w@����ds֩< ��p �n�k��1��Sb�{�±����hm�����3.�n,��1���lԘ �����1��#c�n{�.NY���Kt�����>nki�eO�9jqG,��oS�ђS�3�';��x��      @O �  ݤ��o�:�v���k�_�
�g�E?��}T|b����m�xАHF>+R�w�-z���mc�����z��I��Q��N���w���Ώ%~,�pK��S�z���������K1��qAm       �;w  ���7����!�F�>��wފ\���˞~2��	*�۱����:�}�7#QT=Y��pg��uk*����|���n��߻<����z�1�K       �	� @��f��`�(,�|���>Н�E1����}�c聇G��7��N<<��,�_ݯ�Q_�z�Q��s&]���      ��� �Un�}l8�(()	�g�	�.������b�g�
ޫ�㟌�o�'^>b�h^�$x���ƨ�붨>�̌����_̿��       �g�  �E�F�\s�p{�O�/�3���s�E�����c��nM��ۚ�����cJ�8��Hgԧ��	1�wD��      @�p �.����A�͹񧂜t��_< �|T��*6�2F�{aL�����F����S���Q�펱���       _	� @H�d�|l���V��Z,�����P<pP�9�{A�UzL,���X��߃���eR����ww       �	� @'+(-�꓾�_[Ks����F[sS@w�>��(����� F�u^�|ľ�{�|��X���E�On�Q��;~:z����       �H�  :٠=���7�L���$��C�?4H_߭�Kݭb�K��5o��#���Î�����       �G�  ���e�q:��vc̽�ڀ�2p�/FAYY�1���_��,z����5#�F�Ψ��/}9f^yq4/Y       �F�  :QAIITd:���3骘y��S��v:���;ﯭ�%j���vaF}
�z��[sμ:       �;  t���O���p-+�Ǵ��U@w��'����zQԷ2��-ޫ��ۢ�����OEF}�zL̽�hkn
      �|"�  ��l����hm����|7���n�`v�A�(5&V��|�^�z�wW;�،�������+��7       �;  t�����j\P�u���X��[٢x� sE.�P5So�a�QP�Q���Op      �;  t������fό%O>��uժh^�<�g�+_}1V��F@6*(�q�ڻn��K"���������z�~�;���G�O6�>}>�YTl�e,��3      �/� �3%2�Λ��}�9t�D"�57_�ߙ��ߧv�l�}���{����3�'U9A�      �+�    ]l���+_{9�7�8�>v�|�V�J��       �   t�y��c/�"����v�Q1��      @>p   �u��'F�u^�Q���zE��X       �N�   ��66F�ϦF�)ggԧ�OE����wۍ      ���   �ɼ;n��ǝ���~�	Q{�hki	      �\&�   �M�����������Q�o��b�      �\&�   Ѝj�N�8��Tu�w       �	�   t����˞�k��rی�Tn�}�o��X��K      ���   �Yr�{�������~z       �*w   �n�葇�~��(5&�>���R̸���T7?       r��;   @wkm�yw�c�����$��c��GƬ�/      �\$�   ���}{�<��(��Q��s&]�      �k�   �@��1�ޟG��gԧx���׾1��;       ��   d��[&ŰC��DaaF}��:!���gmm      �K�   �DÜY����ǀ��ȨO�qF�6;�ҿ>       �D�    ��L��q�=����     ��#�   �E�=�d�|��(��c��Ӯ�k��b��o      @�p   �2�)�����̚$1����~=       r��;   @�Yx��1��oF�!���c�UG��      ��   �Lkcc��ljT��Ռ����!�so�       �@�    ͻsJ?��((-ͨO���E͔I���       �N�    5-�����!��Q���U1�{��u_       d;w   �,Us�u1�K_�H$2�Su�I�      @Np   �R��|-�>�dTn�}F}�|l����'       �	�   d�yS'gpO�:rB       d;w   �,���G���Q6jLF}|��Ѵ�.       ���;   @6km�y��c��^Fm�EQ2dX       d3w   �,7��;c�i�DaE�       �g�    Y�e�TȽ�       �	�   䀚��c���E��0       �;   @h�;;?�P�}�       �W�    9"9�]�      �g�    9b�3�/>}6�x       �#w   �2���b�]       �H�    �����u�7�dhU       �w   �����w�#O;'       �;   @���sJ�8��((+      �|"�   �c�-����2��H       �w �<1��k���5�YkC}4�-�e�x*�>�x���G�����=��|ײje4̙K��D,���ѺzU��

b�_����bTl�E���e��{����hmn�\V:lxF�m��A竹eR����D"       �; @�����S?��hZ� f]ui��|j䳢��Q���#l�m���}ηb��߉���d��1cc��L��7�|�8�6�%U����A�ʕA�[��k��o��m?       �B� ��T<pp���K��[Ŵ�Ό�����.���m3|Q����o��"u�E�k�_���^ا"�ƚ�Aר�:Y�      �+�  ��{���o}㌈�� ��pZ4-���)�ݧ��_l�ө="����T�ͷ:���!�g����?>�ߙ��       �@� ��7x�c��E����e�����G�3��cĄӣdXU�$K����{�?��hkrW�.���n�)�9�/      �� � @^y�9�y(Q\�9:��� �%
c�~GO�<�T�|V�1�~ �Z��3F�vN�       �N� ��P6z��=n�X��kA~��n�ݤ�㣨_��iVO{3�>����n� =���c��]�u�����;c��'      @�p  o�;N�=�V��((�hm�V�Ъ�fM�<*��TD"�_��o��E��7�����#Q��       ��o= ��}���(*����hml�X[�^T�ڰ:���<~uw����}���쉗G6kkiά��)�U��ٱ葇b�g�
      �\&� @�h�[��eK�ۻI��ڜw���(�x��=n��#����|5�z�fM�eV�0��gjn�,�      �<w  �Ckk�|�� �,��{�z��h^�(����K�~2�Y˪������&w?E}+�6��+S�óݪ7^��~�C�m--��l�����5�}>�Y       �*w  ���g���{4S��{���.�ﮨ:��N��u��ed��o��^;5
z�ޫ�g���+/�\�������3;T�l��LӢ����M��]rM       �*w  r_kk���EA�Y�ʋQ��}A��}��1��F�!k�o�Ϧ���`����{Plp�MQ<pP�/ɋf\�ݨ�eR��t�%O<�>���
��b�՗F.�{�W1��Gɐa      ��� �y3��A�x�� �4/[o�yB��O����)G��[~e��J����#f\��%˟}:^�o�X�WE嶟���q��x�k��ҿ>���ΉM~�.V�3��X���"�55E흷��3�       �H� ��������8<$�4�̉�O=:g&|�d ��������e��ͨ���~o�sJ�64D�i�W�s`��>Q}�W��:c��iY�<��~S̙tu��\�(y~yu�!��5S��j�G�O�̟�0rɼ��#N8#
��       �� �{��b����~�T���X[�w�57_-�V�c�k/�s{�C�?4���'"Q\ܮڶ�X���c��ɱ葇"��9���o�=����f�ԟE�ߥգ"_%戀�^������-˗E�[������E��g��������Y=���B�ǝk�/����C84       r��; @hY�,f^����%ύ����>Mu�#$��+^z.�p�DA4̛��~+ &;�55E�SR������>Q\��}ּnk���>�Jkk,}�O�GRaE�(12�*����0�ArZ{c�ԅ'�(�~��1��?�ʭ��ґc��W�hZX���|�z���es&]�3�Y�}W��=      �\�  Y�e劘3�� �4̙�z@>JN��(MDO��j��rO�i]�*?�H��Y3�l      �$w           ���;           YA�          �� �          @Vp           +�          ��          �
�           dw           ���;           YA�          �� �          @Vp           +�          ��          �
�           dw           ���;           YA�          ���U����QZ=*�*�EA���Z�:Z�/���s�i��)��_��Ǣ��W�Ϛ������_���FQػw4̞��z�[��l��(,/���a��h^��۶_X�'�l�E�u�ZV��%z4         rU��8z�Y7�����>���-+�G��E�0k���[�'HE��6�⁃S���/?����K����7����y�X������m�S<``�T����eŊ���vd�����t��s"�ܨ��N,���Z_ts�=����S1h�/F�-�M��?HS��X��gb�C��ŏ�>^�7���};�O�d��d8|�/�%�cd��5'��_�N�m�5�P����O��/�N�{��~��s�'����c�ݷw�v�?D�>��1d�C#Q\�%�&��?m         ���z��=����|&z���sX��W���^�E�<�u4̙y'���#����E�������so�.�\U��4G6K�A�j?�����Λ:9fM�<ښ��|�~���?��d��W�9��w#*>�u��Υ�k�����M�b��.����=]�ܓ��A_�/�O9;�F�nWM�!1`�=S��+so�5�ޘ:A�d0|��_��G��j��w���;/j��*�B�x�/R߫������Oo��?� j֜��Oɻl��y�{��        @��o�i�:���o�O�k}A��Q�����賾u�����<{&Tg�� ���U1x�����1��s�b�-㵓�薀x{$A'����=-�]#N�J�Y��{m�!�:͝�� �������q�N����b��'��{I��w�Č�i'C��֜��xx�y�I���D.K^����؇��ל��9��X��k�왿E�I��6������gQ"�|�;����b�_���z_-�        ��d�����Ĉ��L������+f^����������eɩ��n����K��ڷ��3�Ѩ�|��[oc���x��_�[٨11~�]�5���c��/��m�ܓW����Qԯ�Z�WZ=*��zo�y�	��F���Q���>r]�kԙ��K���f�HMi�Hk�D����_��K�M7��;�         �Or
���N��mvX;�JKc�yߋ�n��?+��5rQ�1b�i�Z;��#c��a���&E�İÏk��!so�6�gN�׈	�GAY��^�H��3�&��R�����k�oAII���I��i����~�h��{�{m�V"�[4-��l�N���&���C�qAm�?�}�}��         ���,6�|G���6k���}J�{�7���I��vܵ}A�����;��n�)�I��vL]p����f���A���n�^[��'Rś�,���K�E��b��n\���w%��c���Ƌ�6V��V��-�-�����Yp/1�����0r��{�)Z         ��:��S���J��W��b̻���5e#G���zTd��r��f����(.�⁃�(HDi��δ��פ�BMWa��wٵ��������%ɫ�ґ(i�=]��4�ch�U��ի        ��6x��=e�3��ڷc�3�U���$�Lb��$�MA�Y�t���RP\�
��#��]���v�#����(�I���� ��ʗ_         >\a�����d[ɩ�c��^�r�~�+:5��(*���^]i��F�o-�V�u=�P4-Z�         ���3�xА.�^���G��w��|8 rA����(5&�R���1��#c�?�봬\�|�����O�6         =A2�8쐣�|�#O?7?����� �v�pOƈ�N��0���b��7Gk�� ���o���:�0
{�         �1�ؓ���W�o�|�&��O���	�����D�a�D߭�O]��T7?�����w�MѴha��O�����^�C���X;7��Ց�lj��AGD͔�:�u��hmjj������~�hm����ڧ�>k6T�n�}wŒ'�!��o�z=&/x�Tayy��         ��x��v�Q+nm��ښ((.Ne+;b��g	��am�MѲjUZ5E}+�Z߲rE����{}AiٚGi���;��.�6
����se��D�[ŰÎ��O;&�=�d��S���EQ}�i�%��3.�v��u[�55�B����7ֹ�Gi݇{r��9%������Ƃ_����a�]���5s��]�Lk�6��(9:rA�º�3��ڳr�b���O         �I�Q'FA��i���枘q�����&�q�F����q�o�iZ}*6�DTn�S,}��t-y�x�#ڽ>�\���o���W�90V<�l�׏:�1�����n�mlp�M�(*~߯U���&�/��X��]�_�p�חҟ�����vt,�ӣ��TKK,��ݩ��F7ܙV���Cc����F�         t��~�cءG�]7��?�i�<3��|��W_�W�> 6��Q:bdZ�F�r��;��D��w/��p��
�zŸK&��{�m-�]�ok=��<�'~%���������ג??��?�gZ=Gwj̿��hml         ��0�����OZ5�jc���_��w5/[3.�^�Ť�zV|b��z�X��_��*��1z�3�]k{�}?�u��;�z�}�_l������)fO��C�̺�����[R5<頨���          �j�}c�!�Oo�{��hY������Ī_���O��p��&Oo�f��р{AA�8�����{W4̙��kV��z,|���ٽ��=��3b�/����jmlHo}C}d����n��9        ����ۋ�V�UӴpA����_�����"����zWn�Cj�?�\���*�[���I����w鞗������V�?���=nôj�ZZb�۵v�՗���?���Ҫ1x��c�=w=WÜ�i���5#�Mc͜�\        @�INov�qi�ͽ��h�_�������Mq_v�AA��07�\e�왑m��Ms�\�I$�[������9���H���׿��o�kmr���G����6F�ٯ��m-������z�a�Z�<i�|���6�c��n�v�mY�,�?��         ��Tq|�S���,�ڟMm�����~�_1)�m��~��b�X���Aϔ��7/[����G�l��GS��Da���K�x,�k-�>�3{�}Pjz���Ҫ�uե1`�=Қ�^6jL�¾�ྻ��)_��?�Ϧ��ڙ�_��٦��ۢ��	Q:b�G��3����        @OQػ<�;6������+ڽ>5���W������N��Nl��X�O2c8�+c��|��d�}�?��l�8�&j�%���u���2���[;�D"u�KW�����w��U����RO��>���ό��ܓ
�����_9>��rO������L�:���F��ͼv�1�滣x��\���b�        ��3��㢨���j��.�y�ߔކZ[c��WƸ˯K���λE�M>+^|.��N�.�7�8}a�\���b�7Έl5��D�u�E�v;~������3����Ǽ��p���|�M�+Z�$�;��mo�Ov�#�o��Q����흵�e:_�����������������q�Z=�͘u�ũ+ٲ٪�_��\����G�]>�_����S�d�݅         ݧ�W�:rB�u5�LJkz����u�8�+�{܆iՍ8�x�ԣ���5�<��X���Q��PZ=��_j^�4j65��M��V�����C���3�ꘓ�+mm����c���O���k%��<��k�C�IMc����]*X����Zs��+0z���m�|８q�l�����"j�FÜY�+�����^2�*�l���c��jb��O�y�         �W�a�D�iմ,_�n��cLNq�.9��ڴ�R��o+_y1���b�ݷ��a�%C�D�e���m-͑ښ�b�5�Ŝ&F�[E鰪h^�zZ�����9*�{r�t�iY�b�}��mw���c��?���^c����?��S��|�+v���sYcmM,z�&         ����G��v]��ɩ��� <��3қ�HĈ	��_9>�~�;�G�JN�_���A��8�^}ҙi�$��g.N^-����G�d�=է��f���         �u�>*�J��e�ʨ����w%��O�:�]:1�����+z��Q�z�� ������������Ŝ믊�!y;���t���^o���f�#         ��RPZUGMH�nޭ7D��Eo����Zw��%���pz�y�I�2
�W����k=��X���6���?�����i�U�rvj?�a{         ��a�AGFɐaiմ�^5�LZ+�oki�9��$ֻ䚴�~n�}�e���i��:p���Q��Vi�%O�kӬ�.��;����񛬩�5��         ������Ǥ?}�S�i�µ�u��#�S����Daa�8�x��@w�p�}�I�Oo_��#����bm���G��λ�UW}�Y�         �Z1�âdhUZ5�Q3�����)��_��誴�}a��}�O�~��Н:p���S���ۤ]�<av�YW_��Ȟ��>�m��B��/         ��Jwhz{�S�qA�Zߟ��ܓ�Ȟ���O�i� ݩC���?y%��˟}::�ʗ_�%O<�v�tZuէ}U�         �Ȑ�����i�$��Ͻ��Nٟ�Nq��1���D���]��Wl�U��r۴74��+�3ͼ�G��S��5Ž�㟌ʭ���O�%          ҕ(*�ǝ�v���o��ښ�,�)��'�ecҘ�<��O��/<7 �K������Z��?ǲ�?�)5��/�~;�V݈��p         :dȾE鈑iմ55�ܛ��Δ��>������U7d��c��WE�����
��&�o�C����GW�}�eiܓ��n�M,{�o         �^���NK�n�=wtI�|���'�e��mwM�{r����;�py�9io`�?��eO?]a�������wN����3�g�          �5���Gi���jښ�b��+�{��EW�U7��Ru��5���p���Q��Nio`�՗EW�}��iܓǕ<�d@         �$
c�	g�]�����}��U��&�ٳi��=���Q(��t�-EdoPE���YV�� SP�(@fW�������[���7�~ޯ����9�i��=�|���r�5TJ�Zg^������OpX��O>SY�^) j���u�ܲ�x����P��������y�����5�&              ���d�"�Mp��Ө~��JNc���j��7��/���sǍj�� �~�ÒS���r��{����@ɹ�����Tx�X5��              `K�N8��>�/<�ƍ�5�J���2ϸ@����OHt���8V�+ J�
��,� O�����Ǫ|�u����(~���ǖ
I����}�o              �9�'+nϽ]�c���ܪ��mq�t��\�z����~��,s���wޤ�s����&q�	�             �-�x��j����Sc�:��g�T���jq�7QQ;���> ���CG')z�ή�a�ZU�񚆓��W�������}"'O�<OPcv�               ���`��}��K��Z���[q���F-ڟ�;�!�Հ{���Rp��-z���#a��[����
���S�؃              �)8,L���r�O�'�Q���p+y�I�������{�U��s� `�l5�9ew��ѡ����/����*W��ݵ�             ��1~�rw���g����T��?+��c��O�3�� �(>�p��2���}�����l9��w�P�A��{��i;
              �/����ާ���WT�����{HL���2Ԕ�+ 
[��L#7j���|I�'�vp���.�              GĄɮ�o��TÆu�����>���p0d�p��%�z��5_ʗ��|l�Q�'�i              ���j���}+W�\R��=��χ��J ���Cbb\=`sI�|IKY��}B����7              @WV��FKI�|�e+�܃��eI`{l5�������K��j]�c|�             ��B\�*�%�8��jk\m�!�`�l5���֦���~?`PX�|��?$���E               =Y��_�U��(����*���m�Np���?��%+��'����vf              ���},WiBF�ڞ\%�����{]�B]�#�O�/������mfU[C�               z�\��&ɗx�����j���j�P�j����Pc����w�!_��LW�7��H �ܶ76             ���\m>v�B���V_'_��.��q�� �T��)�hm��M�j{ϨD��IQs��c��j��~���ޫ�7g��BC��Ңa�Q�.u�K��_@`��駞��C�TxZ�s_sa�J����U��U            �֯q�}PH���^��"_�6W��v'K
`hM��V��1����+��;T���A+�j���8$:F�s���5�bg��4W�ԯ�R WĄɚ~��^+Wر�B�������            x�~�z������{p��ј����z��?I���Qq{�պ�_�����7�p�����4���D��>��?|_ �MЙ~��]�Ǧ���>=jM�            @ j.)Rsa�������^1왣����9��>�*�e�aG���P�7�f�{�����9�z���������~���I���p��}��jU��? 0��x�"�M��v�&8m��7]#             ����)�{������J9�D��{���e�ܪx�/�����L=����r�q�p�hkUջoj�����(���g�k���vn��W�T���ڛ� 0%xx��=��            @��tp7�'���GW���N�!v�=���"W��75���o ��	U���*x�}\����Oϸ
���C�T�=��a�:5koO��	��+y�	PAA��8�ߛ��g:�*�             �T���Z++�I��}<����*���4ƞ��}��������'�c�+�n�K4fg)b܄~?���g�q����g�q�������x�uL�aa�ǭ~7	��"�       #ЫՍj������RGDx��B��$�em�*�[߰GF�b#º��\[�����1)�e��'(8X�����
�n��v��GHTt�����Z��  P�76���*���\��óU�؃j���P��mO��[�z��� lI{sӀ?f�Ҝ���Aj¥W�z�C�P�]�W���*aɩJ>�ݲ�����'         ��M�5�i�POsS�U��PO�BCC�o��U���B��{����n�mܸQ����'��;���Hxx�&M�
wdd����r��ǣ����Zr6���o 8
P�?<SA���7Y�{��'y����ܷ����C�~�_����ŀ?f�늿�it�BG'����9�����iow7[���\�O�          �,�����^��SN��utt�
��,^F� LsA�J�Z�G�j��nq���}_����s� `KZ��T��������7�+���4��_���9�9�5lX��6&���
��������         �������k� � |��zN���;_��{G�  �#���k��G;���5�-�c/���}�>�To�M �%���	���Q;ٌ����r����3.���3/TpD��}Z++T��#         ����D��޳�=d�hE����O Gc��oZ܏8��~C������$,�rn��I[ 6���Mٿ����ybP�U��Z��[�.���?2-�aɩ���0�+��e>          ����>����w #Aπ��^���;  �����|��}������ ����&5���T��}����A��\�M��(�3}��=�mko/\��          ���p�7����������;���U='���_���  �4fg��?j�w�q��`�����K�{��z��;n��`m��p��%�~t�R�;����~PY��RC�u��iq����e������t�9r�������v          �p�����kjj ���޳��3&E�g��O ,�wݬ�C����q������T���0�:�7�VWɗ�����뀻)X�Ri'��3-��j�֪J>��     ���V���*55�  9�s��E��jt�G�BC�wx���KA  �/.W����+����, )z�M̒e�  9-�/>�1���~���n��qs��/�Λho0�)��K-��is�q����n��     Y����J56� ^m�kGƺ��v�~�9��9��x��Q�:'&H�!�� ��g�����R�����^���`$ioow��t�`�J���  ����I��-��^�z���_��o� ��6܍��~ҙ
M��}��=�ݷ�WW�h��    �� �^kk����;��Vp����hYl�Έ��  �h��N�}��poia�5 #GG�a��>y��֭  ��J�{�����so����z��� �m�;-�Y���]�7�-��ޞ��c]�g����    ��V鼼*�� ������Z�TIOEDh��X]��/2  ���UWW����(!!�������������p� �-��l[{{�__ ����T��~��tư��g��#���ڧ��Z���     p���nqa.W emsv1��ڭ��F_t]546굂F�S����uB�   F���Xax����
�6v>�lkk �$}ܣ�-Rٽ�
 x���=~���s���ro��� |�vܝ���ո]�j��hqO�T�w�q�_~��K{;    ����cƌѸq� 蛅ۛ:��֜YSS㌦ͬ�aA����|B���ɞ   ����N�� ǰIMM�u_]]� `��k�x��
���� O�7[�{���ާa��*{�%����Ճ����Ӈ��=s[���O    ��@� �MPP�"""������g���2����vϯ���B���Q:%��;  �}��'&&F�������l�% �D�Z�;���.]�rr* ��7��O�j�aG��o{[���-ܦ���;o���O��{[}ݐ��[{���;LA�I��    ���
Wzz�3�ѽ���W���E�胤Q�31t�_|  dqqq܇�M�LHH�v��C	���jq�^���; ��;nR�����̳�z��ukT�ʋ _2 ט���=�ܷ���8w    ��#�/k͊��r�u�Ƃ�7/�DGGoھ��M����ޯ���tq���-����Xg��DAA����-��ߙ�����8=���  �*[�&//��P"ׄ	�7w���uB� 0��+$$��};̐'9U�Ņ �����4�У\�-�	�,R����s）�v >g@�N��#�i܅?s�߶��;��.��`��j��    ��}�*��W�-ܞ��D��X@�&*Xß7\�������3,1,�n�^�vAa�����Tii��-))qn[[[�#� 2e���<''GM]���U�:��M��(y�  ��gع-�CoҤI���� `���{�ף:ߎY�U>��  ��iq?��!iqߖ��ƍ�U�� _3`�>r��O<]�Q���g[Z�3Ͻ�}{���    �������m2BJJ����7ݦ��:o�5JAAA��i:���/��(..vڮ����m�Ys<0�y'���uQQѦ��j��|�ъ��_  ��X�;��e����ޕ���a ��Z$f�� �,@>-�	�+v�^�?���oT�( ���{C�c/����ܴ�G���1��oo/����r�,��{{��6`�N:P�u    ��#����b�я?^'NTFF�F�=���vQѻ���z/2z��~�p���y�}>�P���2���9z�����ݭ�݂�66nܨ6(;;[���F
�����t�JYYY�j���N���(��q  >�&��j4L<:�'O�u��
�W0 F{��^?�*b�
�KP[u�  �i(Z�3Ϻ���՘�Ae/?/_��2W�:�8���\m�A��d@����W�Ig���37-�g���A޴7ԫ��{���\m��!_�	UؘW�؄    (4��.k`�d�[�����v�������v}�n��m���k��n-��maaa��vk�o�y�>����ٳgw��Zӻ��mX`�F�vl�Y�}�w�ڵk�����^e55:)4D��	  ������&nO1����W����B �l�N�ׂ,���;�z� &kq� �������}�lS{��}9Pm�O7�},Wi�~N�*�oh����F�3(-��ޞt��?��U+�R^&_���Śĥ�U�����@���i.-    ��}Gxx��M���v��	�ڈ�����v���M��K�mnnv��mo�p���mx�k���<��F����HOOw�>������J}�����/��_:!b���k��ێ�֭Suu�s���J]1FW��J   !55U���4�;o��qmў3�y ���Z�c.%� .��5��ÝB���o���s.v��4fg��O�ʗ�V��U��<q�j���/S�����i�</�����jq����{��s�:�s��}�~(v�9���?5�lY�q���>퍍j.*    l/�ۇ�5Z�}���Θ4iR����"���-�m����v�m��+�n�v��o�=22ҹ��{O			�3g�3���[����m|��*+�����f���׫��
)*���$-t�*+�abK(�M�.l��ο�����R�B\.�=��s
��r=�>ߖ���_�z�~X�ڞ�ax�sq;�����6�'�� �I_��]�PPT�:he��崸��y%��wk-�.U�.���|r����vӘ�������<�be]������]��$W���	�ox��iq�^�=�'���wk���^����9��[�|FK��JG����4�����G�a�Z� O��\�{EϘ�j��O�kgt   ��A�}�Y�c��w׬Y��`{JJ�V��>o��h��hE��}-�m�=Y��v���}]�S�8蠃���������G�|�x������`� �M~Y�f��sh2~ST�}���� \HR��nH�v��w_Ps�F���R����m��w�e����	��իW��ݷ�aथ������Ad�-=W��牬J���ߒ�+���+v��T��� ���~����=����s���>f��.����ᴷ���|]���?�N^���N8Uk�V�Vi8�^~�ƞw���j?�� |cP�#mjq����>vО��{��Y?PÆu���v�e����������HP�Ͽ��'lL�f������W�m(g�v������B����z����    l�/Z��򪺅ۓ���0N[3��ٳ�1an�z�v���z���9�6,̊m��{ۯ���QTT�x���v�������ጃ>����]�V��3>��s�nˇﱟ�)S��믿v���㲪(]���>  ��f�*��>x�y�3z�o� ����=f�R� ඵ�=��:�ݠ���&��)$:FS��MQSvp�y��s�Ϸ����� 8r�����IWݠ���T�7�1�]��
KNU��+u�ɮ���~�Wj.)�oJ�����icw��1a�v��۪��j*�SxZ����k�v��
�xxD������pB��'��/$&V~~��]�5t�Z++4؂��>n���Ve/?'�7k�s�Q����7����o��K�Ԭ?���\>�   ��}p%$$h�w֜9s�a�ͱ��7�n�������v���6���w}�Է�z�����5�o�{��o�.RZ���m��������������݂�6�144t���u�6m�3�>�h5u��X���?��￯��J�ͻҀ5���?J*�.&I�ɸ  cE�92�u��k�lo����� ���׉"g�%�k6 @@˽�f�-�A�?,̞q����S��+n�}\{5�f����5R����2�������=g4f�Ssq�:{ź�`'S9i�6������ |k�V.x�>��x�<�	���wܜy��o�75����5��<��]t�6�kK�D�4S#A�������bO�&^��|�a�;�3f	   �����a������^{�弽9h���q���@�P��[x���֤h������ �7�n�6��a��@�ݭq�����ykc��2v��!6�M��u���u�#6I��N^���N`8��3��g�����>��
,�si�[Q�����W�-zdt�   |��w���+''G8vnҳ��΍��� ��[�еX!8*Z1�,R�  p5�[��W^P�A�u����� �vȽ���h9��J����w3!�++]���:ZZT����A����8!���]��V����TC��(���iV�Hb3�࿦\�{%r�   ��@s��;v�j_�`��v_�"��-�nm���>�v���ٽo���,`o�k{z_,�n!x֦n��~� 5��cY��x���t�v��`f͚�SO=UYYYz����[o���@�@���Wrr�dZ_^��I����   pع�=���00��s�M�jy�sB���3+C�y�Y��  ��y��8�i�JMy*y�)�$��Y*{�E%t�������[�p7N��Ns��=����N�4m5���	?���U�_�����-��Q�n  ��!�>0RRR��v�O�>��m�-�h�p�@�,��kl-�o��QQQ�>fw�H�s����mx7n��{\\�s۵��ڵm�����ֻﾫ�_]EE#�H �-##C����D�����@⠾D	  �������W_}�L���?~���+�<`�	����7$z��
򄎨�\ ����җ�S��G鿛w��NS�H�}㯕�t��#"召L:���A�zd��[���+��P�_y�ZJG�Rv��V:K����U����B~s�࿒�Z!   `0|�*��W�-ܞ��D����k�h�"��}ҤI}ncjdK�7��5�n-�#��}���-&&�]Y����� ��m�|`a���*g��þOv�fmk���߱+V��c��g�}洺[��5���&Y���֭�ڊ*5%&)\�  �o�����ӕ��'l;;��3gN���\&?�fB ���6����=��� �6��j%.]���(���	�DM��ʹ�w�/䏲~{�����A�G*zr��=J���1�����
���H��֪�t�f=�y���/:�ڴ��粄����qg   ���mc�љ3gj����{�{-�l,(mg�7u��n+�[P�B 6�}�۰��}߬e�xߖ�	v���FAA��}KHHp��{��y�q�g�����o���>�h�����g�&V�Ě���ua4�_  ��IMMݴ�ܳs	[A�����{���\ 0����E�!� Psa��o�^~��!�������'�T�ܥ���Q%�'%�>��?>. �z����_�w�f��U�%��?�ޮ��^���:�dM����5��'�'a���+����Y��ּ��das�=�
4��
  0�hnwϾ>.���ݓ�-�n���ij��~{�vk��Z�����o-�t�����[�{_Kao���9#22rS�=4��s>�>[@�FYY��|�M����*.���axY#���ެiԅ����,  �&N���?��@�6�m��z���y�M �@a� 6᧫�y���B��f ���{;kw�>��A�w
{P�Ｎ��o��?:C3yF�;͔?�z�]�����v��w��_�җ��z���gH�>7�髳O���O��0(�F��ר��o�T�����M��}
���:O�l���U��ߵ�����\\$Ә����t���*����  0X,�~���b��s�jٲe�5kV�F(aTTT8���	�GDD(66�h�ya�Ϛ���#c�wo��$n��- o��m"�ݭA�;�a���:��#u���_���^}�UZ���\��kiM��R�ą}  �{���I��f���0~�xM�>��}v~RRR" $V>г�=d�hE���  ��oĺ�~���I��3oP����~����R����F_�~������w������o�s���f����&'g牋W��bb�4�۾0OCe���j���>?�H�x�c��s��w���'o�U��t��ݶRacR4Ҵ76h����O�(������s��#"��}�����T�������@Q��_  ��A��RRR���%K�(..���좙�"���os3���-|j�mTo�7F������a�,�n?v��b52�����w�Z�Az�w�̙�kr�F�W^y��ؚ��T',�t�!�����  0�bbb����u�\������5o^�p�M������  ����E�� m�uNh{���ըE��c�|�/}q�
'd�/ZJ���	�մ��Q����J����_q�߇۽��G��sp��mX��u�ۧ��o���vU��ʐ�^��g���%�z��J�w�v?���o��
�O��fO}r�RM�����k0��y�O�S�W�+P����P�)go}ۚj�~P���G�v��>��ٓ�ܻ/   <���W�-�n˙n���ɓu�a�i�}�u��]5w>W��v�[�٭���M�vp������&)�5�va���ޙ QUU��vw�϶��}<kr�N�� �I'���?^����~�iegg�;�ر���1�/U  �b�Y+yVV��y6v�����W�\��h�����s5Ę�Urӯ ��2�/����N8U�r��<�_:T��S��9�6c�;��q�9�<��~��7��������zL�$��;4z��~��w���jX������?p�ۖ��G5fo�P�F�����t����K��!��'�e���웮�/�ph)+՗g��QK�i��?��5�K���m*\��:�Zhrn�N���V��6��}]���\����ߴ�����Ou��	������ẟ_��  ����}���{�C=T��K��y�j�Vn�"##��FBB�2E`����o���fw�v�$
kl/))q&Ex[��-�n��E��O>�/��?���F��~v��w  ��lr���me#�f�m���+���Q999jm�k� ����!��4E츳���  pt����ߪ��q�B�.ݦ��_��rn�������Z{���Me�����L�����P����E%�=��[�s2������h㍿��K���v%�>�L���[w�Ŋ���"'N��6u��W]��4<W�:ƥ/=��������4��S���nu&Mc�F���'g�;���_U��u~�h̡G)aߥ
M=ܟ�Ӣ_��?T��3*{�E��@eK�|~�1��+�r��{ͤk�Z�u��X��C��V���5�_;���G[� �7����  `�n�Η.]��?\����>f����2���mP ����B�־M��&:�HIIٴ�M�h��y�]����-�b�,{<'�n�2llܸ�it��inD7���� �  ����Ҝvrm�[6i���]��ڹ�5��9 �>[ܗ.'� �~͗�����L%q��MJ��>VLZ��_T��sέ�5���,���L��r��v����);h��J���K�[p�� O�,�j.*Ԅ�����s{C�r�Ey��&+.��1j�O�t��A!�F�;ZZT���N!�}��Ұ�"��B�6,5mGEM�Q��xGF���Um��j��Q�W�9m��Z����3,89y��&MSXF�<�q

�PB[M��K�ո~���T�(���7\}�������Y����j��w�N�����l���QXj���@pD�F:��	
�?�   xn?7��[�=)))���>?蠃���c֮]ZZ���JWm�d��������l���X�݆�-�n����R�ս��PEEE�ϛMT�\Ə��.�H+V��SO=�7�x�G8lr�M�(l�R}�`  ����d'�n�8Y�蛯���k6u���$ ;G  l&�>�J���  �Ӗl�ח)<=S�3f)t�'[��v��Ԩ��\u_~���j��sn�����=}�"ƍ�'!�ɢ����{Ҹ1��|޵��?=�򿼤���9y��q�zU���Z�*���Z]�u��Xo�J���)ϨD���������zX>'�Y�זa����CG��~��[J�Vdͅ�    �����l9�C9�il����b��c�������ߏgm�h��q�VVM�b?76,�^__�L���{[[�����mg#66֙�b��/�?�|w�qz���ꫯ:�6;����7�H�  `����lբ����
E�?�s��e�-ܾ�� $}M�
;Aa���y� �%M���@�X����7���Ԥ�����&�l��|&�    ,�ۿ�C=�W��B�`��%�-H���贿[+20�g�Fjj�3ᢼ�\���[ݯ�����h͎6��~.�����N�QG��_~�e�1�Ɏ[�m|� ��b�oM�6�	�7���;Ｓf͚խ��V��U���= ��g���e*'�   �B�    0�,�~n^U�p�5<Z�ݚ�:� '�k��^���*++s���֖g�v]��fb-�n�B<t��---[��Zڭű���	���t�ۓO>YGq��}�Y���[},��<Q]����r  ��b�w�i'mܸ�y^��´��{k�ر��Ц=׷U�  }�3�>���]    �#�    R_�}no���l�����+PX }�ҥZ�b����0{ii�3��vg�`o[���֎�f�ktOIIqZ�mR��n���sss������ϯ]ܵ�˓N:Ix��z�)���k�>��S[i˵s  #OHH�&M���egg���C�����ϟ�m��Mf���sn ���߇������Tk^�    |��;    `�Xs�9y�jl����\�����hٲe:�c�����6������ѣ�A[;|�M����sFcc��l͍[
�[K{~~��������[��9���W�Z�?�P�����K�Lj   #�=��Fw����ʟ���n��S�nj������Mter* �O�w+�X�\��   �op    �@����:��S{-�nA����~ۭ-�ڮ-�n!w�Ywff����TQQ��|[�}sl���B�w�k�}�ĉ��+��g����W_}%��g���  `d����;������|KυG
;��s�=�龺�:�y��� 迾Zܣ�/!�   �@�    0�l��ͫ�n�k �����u�	'8K�{y��6,ܻ5"�� ֎mM��H`�0���&dTUU9?�������t�Ȕ��M�̘1C7�p��{�==��N`�)�k�  �gσ�U���Hl8�����n�Ͻ�����Ouu�  ��߃��;ΐ'i�ZKy�   �"�    Tn?'�J�����Ǐ�?�e�>�hz�
uZ��ih���5Z{Y�݂��X�He�2,�c���V������XdNN��{����ib�M���?��z����	�p  ����~n���`�Y�k��9�M4����|ւ�}� ��B��]΁�:�^�,Y��?�   �op    �/Z�s�*�5�[`۟����ԢE�t��';�^/8��-� �5W'''+,,L�?���qF]]�`�R�ccc�����	t����p�X�B���w�j�*�����	�F^�)  �Vy<gu/;ϳ��5��ڄM;�������ӝ��˞��*K[��
 p���B��p   � �    ��~n^U�p����s�}�̙:���5aM�Y�݂��Y�=>>�i�#�gaub��{ee�f[ -P�n�:���7�"�K~��iɒ%���{���-�|A  �oޠ��[#zEEŰ���k[amҤI���r��ؚ�UUU9+, �5��*]EB��V])    �    ������V���q�}H����Ȃ�'�t��-[�4�(9���-�nM�)))N;5H"""4v�Xge�}� ���$ٶ6�ar�]v�-�ܢ�^�=��ϵ`   ��]�ȞۄO���ڪ_��B��|�����v�����4��sn{ 0����}��x�h?U��    p    �@�ϙ3Gg�}�F���>k������-�k��l����,�nǈ��z'�n���XÙ}���\���Nۤt�<�H͛7Ow�y�����
   )l�fbb�3�5���N[��V<���s�-=��wZ�ݞ;''';��x��ذՐ,�nϵ C�����K	�   ���;    `�R���g�q��������|'��%ہ�EEEi�ĉN����p�͑�Ԟ���L&��Iȧ���ꫯֻﾫ��{�m�   ��
sΣmx�
av�i�t{�B��[�L��}��ޏ��ݴJ�w{{�m�E��� `��p��m�����Q_'    �p    �@	����˗/׉'����h�>k���v�n��w-�k� 6��86,�nA����>��I%k֬q�(ǌ�4TΟ?_3g��ʕ+��o   �, i��s���Ցl  |�M8�������`�j^��   �@G�    ��%�n��s�v�e�M�Y �ZۭQzs�=/55�Y@����;+X�dQQ�3��'�l�	&������q�������nSYY�      |I_-�1�'�   ��;    `;B��Z��������w����yyy�����~���f�� �5��=Z			*))q���{jnn����p{FF�<�fϞ����.���;     �}����\k˰   2�    �m�vk]��������A���m��Y�6==}S ���I"ޕlՄ���>��U���l���X��'?Ѽy���&�      �۰��^�Qъ��P�o�U   @ #�    �&�n�@���d�5D��檶�v��DFF:����hx���8q�p��{SSS�mZ[[������Jeff:M�ϟ��w�Y��~�>��     ����^+?�,ڟ�;   w    �k�n���駟����o�}���***�s�`c��1:11Q �M<�6m��YRR�\��B�k֬q&�$$$8���/׫�����p<     �P�����*��QGk�   �@E�    ����ۧN���/��	Ě���	zK��qqq���pZ�[�;%%E�F�R^^�h���ܳ��UUU���z<-[�L3f����_�6     `8X�݆������{����   *�    �~��p{pp�>�`�|��N �X �B���iK�@�����`����i�ĉ[�������)33ә�b�7�x�z�!���     =�&f�2�   h�    �������D]r�%�y睝���ڔ��������3z�h���*$$D |�M6���VAAA���|���Rss�v�i'EEE��Ns��o��-��      0��۝�b�-T���;:   "�    ����p���������	����zegg;ؾ���;����{l��c�*!!A���jii�͚5k��Giɒ%�6m��͛�ɓ'��k��ڵk     0T���g�{H�hE��/   ���;    `��9ܾ|�r�q�N �.";���f$��4f�%''�jT�{bcc�𺵹�����������Z�n�s,HII���_��zH/���      �Jπ��Y���;   w    �f�k�=44Tg�}���o?�}kx������>���vk������#$$�Yq!..Nyyy���-䞓��|PGq���~�i�iʔ)��;���$     �����ޫT#f�B���   ���;    �O�n��K/�TS�Nu޷P���{_�F����Zہ��������WEEE�����j���Z�p�f̘�ŋ;Ǻk��FEEE     L}�(�IIW�3���g   w    @/�n�={�.��b���8�;��}]@��g�[�3���~�m%��嗽>��x���jÆ:���5i�$�|�ͺ��k��'�     `0�����  ��o�����K�O/�RA� ��/F﨎� ����M��  ����A��9�w�q�E"�X�������>����Uff�BCC����ǫ��M�ׯwB�]ٱ�Z�x��xaǂ_��W����ꫯ
     `��p��g�J���0r�%LPmx�������I �<!m-J-�\�FF��4��k[��i�N���ĩ�W+�|�<� t�^?V{P�����l]��U ��u�:'�گ����|���k�����������Rc�����[������" �ˎ�V��^{�����iw蝹����ാ�{2e����c      ��U&��MT؄�j�Z'�L���}�������) �<��j��T��9o^�]s?�׶�    ���g�������?�̙3���������7���_#""���E���_yyy:��#����k�_|�	�Ϟ=[˗/Wjj����:���
     `������r���   �@B�    ���vka���+��eSTT䌾X�533���# ��&�X3�����ӧw��� ��*??_�r�v�uW�t�Mα���@      ������	�   �p   � ���iӦ����\��B`����]PP��ONN����Р'�|�ij?����c6����=������)--�iq�ꪫ�v�Z     kp����	���<�j��   (�   @ ��p��{וֹ.�H���jkk�ƍU[[�k;kf7n�bbb �_���JKKu�QG)66������r�J'䞘�����������S      �B��V�
Rܒ�*t�   �@A�    �?��=�P�r�)����fmذAMMM�����v�����lR�}�ݧ��>Zcǎ��1;�<���:�C�c�e�]�{�G/���      ��H�S��%�  P�   @ �p{PP�N=�T'�n��띐jKKK�m�y9##�� �R]]��zH˖-Ӝ9s�}�&Ƽ��Z�p�fΜ���:K			Z�z�      ��5����t�/b���NRkY�   �@@�    ���ۭQ��s������o����l�BP����ӝ�; lM[[���^XX��:�ۅ尰0���{����ܹsu�q�)66�i~�y�     p�Zܻt��(f�2U>��   �@@�    �?��/��-Y��y���D�����	&(22R �ƿ��o����c�Qtt������������	�|������-�ܢ��V     l��Zܣ�]J�   ��;    �{<]r�%�7o��~~~�B�)""B'NtB� �-lU����ijONN�t�5����ꩧ���G�E�)**J�]w����     �-�
�G��]!��j��   ���   @ �p{xx�.��2��n�r�yyy*//�]ll�ƍ��b �UQQ��+Wꨣ��ԩS7�o!w�تU�t���kΜ9���+u��W���1     �{��^w�
�x�h?U��G   ���;    �9�GFF:��]v�Ź�c��.�)11Q�.��hjj��?�8@{�g��544衇�	'��Y�f骫�r��v?     �[}����K�   ���;    �1�GGG뗿��v�qG'ܾq�FUWW��.%%� 0����K/����2-[���$���V=��Z�b��O��)�^__/      7�
�G͞���(u4�Z   �w    �S�n����5�\�	&8w,�^SS�m��;V			������;���;���斖=��������L��կ~�L̩��     �V��ur}PX�b,V�k/	   �g�   �����vkB��۳��T[[�m�����l[ 
�|�3��c�QDDD��=��#�B���N�     ��W�{̾�p  ��#�    ~����������5e����iÆNkrW����8qb��) 6;&=��:���&�����裏jŊ�a���+��B     �kp�)j�<{AԖ�   ��   ��p���_z��y���ڪ��׫����X�}���
 ����M!����M�[�}���:��&w�[�{��     @_,�n#((h�}�Qъ���j���    E�    �����gϞ����g(���'M���`8UTT衇�~����e!�'�x�ir�i��t�e�骫�R-k     ���������p  �_#�    ~�������9s�8p�������m�� |Muu�V�\��?^����5o�}�]w�O~�]{���     �-������W�ǣ��V   ���;    �p�n?���`����ƍUWW�m���HM�8�iy _b�qV�Z����;v���x�裏:�s���\��o��ϋ�      ^�ځ�@��������   ��H    ��o�vs��k�ҥ���555�>�	&�Z� |ESS�r��v;^yمho�}��Ū��Ѓ>(     �-�p71��C�   ~��;    �P�n?��t�A9lrrrT]]���111NX�Z���577k����q�V����o�Gq�*++���
     `s���{�&��"[���   ���   ����8AP����>����u����r���{5���{w&ey�������z�Wh�d_Ԁ�A1n�D��kv5�8��̜|3��3�̒/��;���I�QcBL\ �A�H ٗ��nz���O?�=,���Z��]>W���EuEu���{?�~�ӟ�&���߮T�a�     ��\0z��+{��f�S�w   $�    0�$b���K.�W��{����B����OII!�`D2!wf�뮻N	�������/|Aڶm�      �rz��\}-w   $$�    0�$b����H���7�v�U]]����S�'%%�P(�v #UOc�ڵkOy����Ժu�t�7��_������\�     ��b��s��+V��_�o   ���;    ��nOKK�����(�����O���5q�D�\.�HfB�O?������҆�j�*}�ߴ�Y�~�     �ip?�;�|S�+��   �DB�    F�D�{�^��_��


��ޮcǎ�q܄�M�; $�������'������ۻ���T�ӟ�x�b��h�ܻNz�     0�jqO]u=w   $R    0�%b�ݜ���W���ӧ+����"�ǣI�&�[ H$zꩧl�=;;�w�֭[����)S����׷��-{�     �G_��eQ��(    �p   �a,�����߯e˖)����ÊF����Ht����я~�|P���v�99�~�z����&�{�W���!     �'����O�wB�BGJ   $
�    0L%j�}�����mېin�B���n�JJJ��z ����E?��O�?IIIv�y|�l������;�6     �G_-�+�U��   �(�   �0������b=��#��G���������������� �AMM��y��]�ֆ�s��'����^G�с C!RY�#�-.�����+��&����N�F�>ZA�M�uj��4���a  |��Z�S����;   
w    f5�����6�^YYiۋO6n�8{ M�J���/��O|�^�c�&��{N��~���/�B_�����, t��]�sh��+�Ѩ��C�,�  p.̼���:e�o�4��
��   ��   �0���v�H���|EjjjRmm�)���󕑑! �v�ޭ�^zIk֬��g�+ׯ_�k���^�o|C�HD      &�n�\{u���:5��   w    &5�n��ŋ����V^^~ʱ��,���
 F�͛7����.��n�6�C�i�ر�9s���>��?     @<?c_�Wp  @� �    �@"�ۗ,Y�;�C�hTeee�]�G ��M ���+���,�O�n�M�o�aW��馛�g����     ���cu�\���͜-WV��� `����"�GÊG���u,��+�};q��c'���'�v8M��}y"�jJ`N�w��r�����I� ��   `��*a��yyy�җ�dC�&�
�z���~�{t�ׄ �v�}��矷m�=����g�}V<��{�1�^ZQQ!     0��y���V.�W}T��?-  ��	��C��E����ݷ!Ż��um��C��t�������[����u�m������y.*�qy�u���2"���|�~��OS��W"yv�7�P\ ��
b��_{C�v$��p�ޙx�0��Ѡ�Q���mW<!��>�O�W���TUWW���������ĉ�h��.�g���?l�?�����wީ�\_�����     ���W�{Ҝ�� .W,ܩX�C1hw�ۡ����}��cfn�����M���lo.� p�����U8��["wJ�� �CSS�ǕHvL�F\��� .Z����6\\\l��&��ô���&� 8�y�|��u�����W������_�UW]e��O<�      N�p: ��2m��`ۉ@{��D�=S�0���~w��r�R���or���Q^.*�    �?�n_�d����:�0\^^~ʱ�c�*))I ��;~��֭[�[o��n����{���/���Ν;�q�F       p.l#{W��]��v��f���F�h��Љ�w��n�~x�<��ſB    )ܞ���GyĶ">|X�H��Xvv�23k�+ (���
�t�R�m���u�}��������w�
        ��5�����ѤX$$�ɜӌ��7W���Û$WR��I�6�`�p   �!V��iB^����y��GmȽ��B]]]�ǒ��mP p�֯_���M�<�n;�N=��sZ�v���կ��_��b��Y2       p�⑐"퍊v6۶v���1f�`�b�#�T%��c��v$���t	��#�    C,��T����x�b�������w����&  8w&���_�R������CF{{�^�u]u�U�������O       0:��AE:�5���6�ţaE���0�:m�=%S����� "�    ��Ǐ׽�ޫH$b��{���q��ِ; ��utt�g�у>(��m�W��ݫI�&ـ���k�       �É�u�]�B���0�f;�mt7aww���Sj�    ̈́�����L^�Weee
�ý�


 �p���z�����}�n�\.���Kz�����|E�=��:;9�       	+S���D���Ն�1t���ю��%�	����ӗ" ��;    ��w�}*..V]]�ZZZz�gddh̘1 \�-[��1�Νk�M���u�t뭷�����O<!       @b���l�=�Z�x4"?�XT��3��ܩ�r���"�\(��     .ʜ9st�7���KUUU��}>���� �?���oUXX����m.,ڵk����Z���ھ}�        #\<~���VѮ6a�0$�*n��+%S��Z݁@�    p��^����/گ�=�X,f�6���Ǐ��� ���B!=��z����x���o�aW�x��G�{rgg�        #�i�m��ՊEB����N�]v�/Y��\�S�̉T�p�    쮻�RAA��?n�{���+))I ��WSS��^zI7�x��6���Z�v�x�}�{�       `䈇�
��)�RkC�H,�`���e
7Uʝ�+O��AQ�A�    .HII�n��&�������w PNN�  g۶m�4i�f͚e�;::�y�f�^�Z�6m����       �b�.z��7*��-*T���{Rs�Nϓ���3p    �7�˥GyĶWTT��ܸq �_|QEEEJOO��[�nՌ3�裏�_��)+k        ��X�S��jE���B�hD��J�[j�Nˑ'=��;p�    ��v��7k��ɪ��R0��o���G ����٩^xA��{����hݺu�뮻t�w��'�       `�����io�En�R��N��<y�r%�S �    �S^^�N�f������YYY�-� ��QVV���~[˖-�������\��q�F���
       0�����`{[=��8�mto�P��F��|yR�tǨG�    p�LC�#�<"�ϧ��N�y�^ 0�~��߫��D���v{��͚1c����/�k_��b��        ��6t7W)�\�x��Z|0s!D���"-5�d��;%S�hE�    p�V�Z��s������N�τ�Ǐ/��% ���F��կ~��~ؾ���/ꓟ��֬Yc�       .��nZ�Mh8�pP��RE�R��*�ӛ,`�!�    8'�@@��w��ᰪ��{����(9�I JUUUz�7�b�
���ب������֛o�i�       /�P��v#�٪Ί=r���+��#`� �    8'��ԧ����Ç+;�����Unn�  Co�ƍ�:u�
������z�!�s�=��w�#       ���G#
5���v�?��T��I��By�87�с�;    �Ci͚5jhhPkk�)��N�  C�\|�n�:=���r�\6��ꫯ��k���/��}��	       ��"�
��!w` �c����1E��3ANo��DF�    �L�	JVUU�����R  `�0��o��V�Xa��9���:}����W����8        /*XT���!lW��=r��ɛQ(9w    �Z�h�.\��Ǐ+9�:��xTPP  ��c�f�RNN�]eô��}�ݺ�ꫵa�       �G���p{�hX��FEښ�G���Mv�n���'��!�#A��A��7��N��Ѩ��B!9<Ɋ��rx����{���d�wߎ��{�i�gn���>�����;    ��n�|�A�B!�����;v�\.�  Ï9��/��otvvj׮]���{��[o���C       �����X�]Ѯ6��P��Շj(���V)�V��Mi��ҼRzz�222�^�n�NIɵ�����K���jk�Wss��*���ؤ�ΨZc���U�+C��q��L��rx�4Z��]��'�is�~-��DB�    pV�_����TVVf� 3���& ��u�����{�?��޴i�~�a�v�m��,       @?p8��-Qg�ţa%�HS�:+�JG��fe8ڔpkla��/�@`ր?��o�Y��466����񼪛��{��˓'��E���R"7W+��jC�N�_@" �    �S ���n[ZZN,�hZ� �^}�UM�:U)))�!��^��7߬�^zI���       \<��#n�����F�8�X��?���J�*W��U�ƤiҔI*(��Z�Cff��g�����TYY�C�~���&UGjK.Tr�"��t��9�Hb�uU�7�H�#w    @�֮]kC������WPP ��# ����٩W^yE�������u饗��;��w��       ����'�H��c)��~�m���8o����״�Ӕ�T�D�t:5v�X;>�_���۵o�F���U�jN)Vr�y2�*��1�*��,�b9\D�1r��    �!//O�W�V}}����ݗ��d�  #ǎ;�`�����_~Y��z�~�ߨ��T       ���I�U��M��FK���J�(zl�ƪV��fjΕs��v̀|;�2����h�[��[ӴnF�h4j��m$�#��eV<5s���Yf��۟��mu�q�5q������fE+v˗;Q.�����;    ���ר����g�ۇ�� �3��w��g?�Yp7.���{�G���7       �?��b�B����4,�c�<�C��oh\����9Eso[l��˄֓��mI���������[3'ݟL�=
�a
����z�YѴ���|�����+�ԕ2��q<�G[�|A��)���T�)K%��\�:+Xu���{���4�    �0���X�B�����HOOW  `�1��-[�hɒ%������u��wkΜ9��       �ON��&���^�c�8~A�qu}O�6('X��sfh�m���,���3��&�n��j�i`,�y� �}1������谷mmmv���AL�ה)S�0�=��[�A��Y���/���Ƅ�C�veoNq����/l w    �)��.;���`��dQaa�  #�믿�K.�Ğ�0������ڵk���       ����c&(XS:��7�֠�]�ۺKK'hޝW�����4��fs3L	VJJʈX�ٴ��<�&�m��jiiQSS�m�?�Ǐ��<����_Z��\/w K#I��I��}����'0p    �2�4�_~�***�d����c� �\fyVr����퉈M�6��Լy���{�	       ��)����)�\=��(Sہ�չ�%MO���׬Tn�M����=##Î��̳6��Df>��u�����3��&��3zV���ǘ5k�&,���]�k���*i�\��P�]Y��3Q��t�w    @/��n&q�d�a��&� ��nݪE�)//ϮԱm�6�s�=ھ}{�EM       �����X�C�����HHM;���U]9�XK��yV%%%);;ێ������_���x7s�ٽ��ޮnm��ĴٯZy�Vu�w�N��u�L����k�p{5��cQkɓU$OZ��ጀ;    ��4i��.]�cǎ�����t: �b��֯_��k���-[��ӟ��.\h�       �#�öewV�Q<��իe��ܯ�-[�I���	g�b+jONNN������QRR��������aa��ӧ�QSS�o�Ot�(�����4������c����f��)0p    Xw�y���`o{�i.0� ���u��!{Q�a����ߴ���       ����ȟ[����5i�V�?R�*t��k����~��糡���\p�3��	&����f��&�
���k̟흷�h�����v���_p�\I���-5�GB��N�~�Rx�ᇀ;    @S�L��ŋu����}��� $��n�hL3�	���د       ���ȓUd[��W��A�|ZE�t�ǮW~���~N����TPP�����;�����Р��*566��Bs��_���am��C���+��;�dk��t4)v|��y��p{'�    ��;l{{ss��NKK�� ���߱c��ΝkC���n��6�       0@<i���ik8��GZ�Ը�ǚ>�;��N�}������Ϸ�����̣ggg�aΧ�9���J���>�o��W^�]�եW_��vt�QʒO��O�pu��r���S����   `�;v�-ZtJ{�YJ ��^{�5͚5Kn�[۷o�-�3f�О={       ��1l�،���ո�y5������rs����ps�/''ǆ�1p|>�&L����ǫ��V���joo��悃׬����/����+6Q��!�����HH�&�^0UN�_�p@�    F�[n�Ŷ����m�ޞ��, @�2+vlٲE�]v�=��?�ɶ������        ��?w�:��Q<=�p�ލr��S}���6m�>ܘ1cTTT�������̼�)3��������}:�j�m7^�������Re�J��J�M<V����O���J�z�   `����UW]��Ǐ��3� ߦM��p�B�\�iq衇TRR���R       ����/�X]Շz�uU�V�k����꣏<$�����������b���3�[�0ebǎSCCC�����փ�ߨ�7���"��v�J4��/��ȟ7YN@�P"�    �ؚ5k��{������ry �����f�ۗ-[f�ܹS�����o[       ���Jΐ'#_��25l���F��}�CWX6m��ƍc%�aʬ�=k�,�������6��eʔ)������^Ц=�.�_�W�EO�ݗ?Y.?�`�p   �Q������Wmm��6K��� �KO����a�{�WO>�����       e���7��ۮWQѥx_�nVߤ�}dHMM��ٳm����öl�t��UW�м�F�����'ݢ�IK4\��1�rǐ"�    �ԪU�l��ѣG�3G �����a��W\q���:dW���,       @�
7U�ȏQ㟞�����[�z�@ ���beff
#�9�:�|����ȑ#���:�>���3ko��m���MJ��!���4����S��6�    0
9�N�p����W,�-fYC ����[oi����"���~[��z�~�_�9�       �0������ӊ���mS@���_�?��<O���n�&L����{#�9;f�����رc����.X��;���^�Wʔ�5��{W�A����M0��   �(�d�j�޽v۴�� ��9��u�V-[�̆���۵b�
����       \�hW����k�}���q̬���SO���&]RRrJ�#�)?~���5+�644�q���nջｧ�nج������k��cQuU�?߄ܓ�    0
�t�MjllT$��999 �^���\�d��6n�hW�x�W��       �0��ѡ'�*X}��y�wt�e�鮻�R ���׬Y��*�T(:�>���S��f��W�Cm����C-����&�a���@�    F�q���K.Ѿ}��vZZ�� 0ʵ��i���Z�p�����Os�̱�        �)��_K��?l�ٸ\.�Z�JӧOF���ledd���TUUUgOOO���U/��Km����E�i�ţa{���`�.V��#�    ���ի��Ң`0h�io �6m�����	�7�xC�]ww    �Ƭճ�   @"�v�����S�>�~%%%��{TPP`���٣y������a�2�i&7�"{n�>�Y���8������0s��Ϡg�ϑ^��v��'���)S��������C׭�FS��_�{�\���$�X8���J*������w    E�Њ+l;������� ��بݻw�U>Lk�C=���,544    .V PSS�   YǑ�t�ߦ`����Ǆ�����t�M6�����
̳fͲ���΄�����0�����j(&�����HJJ��9�0�#�ir_�`�Y��'M��Gss��g�Z�K� _�D�X�C��R�r'����B�    F��K��	3�d�� 8ٛo�i���io_�r��}�Y   �Ś6m��=z�6T  $���O�ȓ�W,�y���3F<��-�����K&L�pb�֛����	���<&<o�Y��d�Bt7�7��Ҕ��n��#EO�{ff���|��mjj��x�'���'u�a��>���h���Bެ"��;    �"�W��m�5K��	  zTVV���L���z���u�u����W,    \�Bj�P�� �����Ͽ��������.ӝw�)�����3wh6+l�h4jC�泛&���5\�<_3�?n���/s.Ԅ��0�F�;s�	�&��B����Fm�ӟ���G���n�ps�n�<i�w    %���m+��1L{��e�  �y�wl��,%k���͛�m۶	    .Fuu�:;;U[[+  �Dw����_o����q�ݺ��[u��W����yfn6))I�%������>��碫�ˎ���m���3�Õ	�ϙ3ǖє���q|���SZ����m������p�������JN���   �(a��{�4W���  N�w�^���9��[oٟ�   \�cǎ)##C)))�  `������?߬�}��z���g>cKE��#�ٳǆ�M�@1�v3l.B4�#=��A�yR3LC�i�7m�f��MI�ĉm(������d%%%�\z�~��o�]������<O�z	���p�����D�    Fh7����v;;;�� �tfBz���6�n�r���km�Mkk�    �B��VCCCB��  ���u|�����=��3g��Vrr�}sQ�	7O�6M��|3��*++m�}42+�VTT�aZ��J�yyy�x<N̊����{�n�F2s���ۯ�����W|I���!y��XT��R%N�w1F�    0
\z��
������Lx  p6��}Ŋ��fǎ���+����N    p��Νk�9����Q  �Te�j��Z�HK�Y�c�T?��O]t�TMM�m/((��2�*;B��pBgg�>���2{Մ݇�J�f����ې{ss�)������}��|���0�3��N��u*XwD����w    V�\i���;��  Ë9�a��/֮]�t�UWp   p^���m�BKK�b����� �H�~h����u��5�y��tꓟ���S�/�����ʜ�MMM����\!�f>�����aZ�ǎk[����Ps�ݚ={����o/z8�؃k?����:�W���C�Ϳ	�/E��\���;    $����<h���� ��ٲe�����i�1���$    ��.i�A=L��������  0Ҵ����㍊v��y����s����O�ޯ��\,�g�{��|J��g.�zNkk�p~L��9�jZ���1�yzڴi�uv���3��}�����~���'�4n��<�pC���$��v1p2�    ���.]j'a��C3�r�� �ѥ��Z���***�;Ｃ�˗�g?��    �\�&�H$bY�%�\���.UVV
  `�i��k���G�}OKKӣ�>�q����7E${��L������#G����M�8��	������\y�}	�z���f'�㶛��w�ѮhX������`�a%��)��x2.�     HpW\qE���:� @��[�ڀ��������O�	j    �0&t�;v  `$jz�:��O*	�y|̘1z��l z@�GS�m�8qb������qS|��e.ڬ��Rmm�]��sA�P)((�!ws�C��=n\�Z�߽����'������;"_�$��;    $�@ `����o���� ��ڹs�>�я�%OMC��ɓu��      �hв�5��mg���vn��M��i��������ڪ��R���+��B��Ǐk���*,,�r1��9s�v��}F���5�Y����}�9��-��$Wk�ܩc\(�    ��.��ruttض]3�f�� �\��a����Z�d�ms7��p      0�����M����<n�_�җ���2��k߾}�7o�\.�[�fq.�Z������R��Ŷ�(�ջM�ٮ]�l��d�ܸF�<�s�9��_0uП[���������A�    ؕW^���f�5�� ����ڀ{MM�n��f=����)       HTG���?�Q�����&L���n7L���������\���ڳg�=;i�$��`KOO׬Y����~�Mz��?R��ays��y��1k+�`�4D-���   @�2�3f̰-n��.W ��24������Scc�&O�L�;      ���>�}�"�}7A�G}tH��=B��0|444��1s�Caa����	��ܹ���~�~���OMK�$wjΠ>�X�C����f�p��   @��������f[v��t�� \�;v�k������w       �(�֠�߾^���>��_�␆�1<�����R���jʔ)���r���!ws���Oܨ'~�/�]�9�Ƀ���MUr'g����0�p   �e��)�0w  .�	��\�R����馛��O
       I<ҡ��	uU���Y���Sr���1������w�����5nܸA-!������ӵg�[��ì���m��������!9�L��#J*�a���w    H@iiiv�b߾}��|�H  .���?|��]z����N�=zT       ��q��Cj��Z��Mp��_��=|.?r�-#�:u�=_;X����\���O�o.�x��K��׾����`��:n��'=_��"�    	h��6�h&Ō  k���vR|�ΝZ�d	w       	����Q����<��z�j�*;GjB�.����aLa̶m�l���KAA���ٟ�<��4��-�)u�mL���r%g�願熀;    $ p7� Fzz�  �X{������Z�b��{�9      �H״m�����y��t�k�QVVV�7�|S�HD�^z�RRR|�Zٽ{����T\\,��1(�׬���٩���S��"�k�6������I�i��b�P���	8�    ����9s��������v  p�B��8��3g��v�BL�       �T]UT�o���m��?�h�ر���	��F���v��~r �Kyy�]�{ƌ�x<��=Ms���?}.��K��د�#9%r��j�D��i����9>w    H0�{�,��
��v @2-3&�nn�I�����      ��(l���Eю�>�/Z�������ٱ�~t�={�rs/,��Ǭ�����y�@ 0��ϴ�O�>�^�a��Ov��V�{?�W�W������j��+%S�e|0^!    �`L��\�o�v]  �˾}�l�Kuu�/^L�      ��U��Sg��>�M�<Y,8��1m��ܑ#Glxyʔ)*))З`0�;vhڴi�����g^��fͲ��h4ڻ�������+?P�G>���En��7{��B�    �	���������  �K8������ƍ���T,       �$կ~W�����XAA��/_~ޏi�Kǌ���;������s�
8�	��ٳ�^QXX8��/))�^x�w��S�����yYzf׫
���K��V�9=~gC�    �Y��:4(W� F�ݻw��S8�I�&�[       ):+v�����1�ľz�j�n}��=O�D�~�z���ۂ��yL$�x<n��vuuJ�NN�]�����v��ïiW�%�d|��0��P�Q��
8�    �@�ϟo��3 @3�vsb���\���#�      `Ĉ��*�ޝ��:�8��xt�5���������ʲ�o��m�6Aw���&��	���S�N�j/�H'N�!����S�_��*�������é��lU��Y��t}�    ȢE�l�������  =������l�̥�^�g�}V       0�?�u����˗+33s@�ojj��}뭷l���[MII`����V�iӦh��<���ӵm�6�:<y�]�-����3J^�)�P�1%%��' �t�    �̙3G���3f�  (���˖�F#sQ�	�      �pֺw��^��>�͝;זz��P�{ｧ��[^5P�z�,����F��9s怆�͜�i�߽{�)�����鵊�򏝩�i��;-G���   @�(((�ACsu   e߾}Z�f�:�Y�fٶ       ���*}�.);�Xnn�/^<������a�Z���m��9ׇѭ����:䞝����|UUU������j̛,�g��PS�ܩْ�)�d�    A̘1C---r:�� ʜp����?s�      ���
5������j�ʕv�s(��*�2syy�v��eW�,..F/r߻w��O�>�!w�bASS����N���軯=#���5�Ѱ­u��
8w    H&����f��9� ���~�ldN�       �p�~h�j~�o}���+�����f��������s�yyy�;w�0:�������:u�}�˥iӦi����ONN�ʂ.�V[*_N�C��R��1����    AL�2E���6l �@3����O(���V$       '�hDe?�L��3����I�&i���ζ��ׯWzz�.\h��]�*�f��4����4�����_�p��}������%tn���[j�I�Ѓ�;    $���edd؀�ph�  $>�dn0TEE�mq7K�      �pR�����#ߜO[�t�����,{�q�F۪m��&����̿��~B(���jhhPWW�)�o[�D���[%ͽA�!�\-wj�N.��	��   @�1c��t��|�z� `��b1���)))I�f�"�      `X	V��_}���C˗/����H`Z����~[�pXK�,Q F���Rr�ࡿ���J����)�333�ػK�5���}2��i�����   @0w���3� �`0�f�{�̙      ������X�����c ��iq7v��a��F��
=c����`fΜ9va�Y)|̘1���;e�UW.ӎu�H�>��n��'-Wr8p   �0}�t��^PP   �	�;�N��      0����O5ny��& l�G2������Wss�fϞ="�8w�hT�w�����l�ɓ'���I�H�w����nz��U�/�Z<V��Q�@� �<   �gB�fҪ��R))) `���֪��E555��ɱ�       0��1����<t��'La�	:��튊
�ڵˮ�Y\\,$�`0h��/��9�~|�z?~�-�9���Ӵ�W�V{��4�MU�a%�;5    �b'N�W�'%%٫� L�Vvv�=yB�      �P�����o9c�	O�0A�Ɯ���R}}�mu����ܹs��c�������`Jժ�����q���.�D?����S.�@����h�+9]��   �7i�$����� G��K���Go���       `��B�x����oZۗ-[�Dg�H"��6lؠ��T-Z�H.�KH���JKK����4ÛAv��}�~��������e�s�_O�j� �@����?ji�W��M�`���-ݣY��c��3Q�3wr�����,�?U��49�y���d	   ��,g��7K 0�L��4�s      �P�~�
5���޼y
-233��ƍ��x�d�y�^!1��������c��|FF�m�?��+�{���ɵh��V{��ӛ,�^܁Q �Ѥ�����}�_��#
7W�s�j�HK�/�p��Iϕ7s��iݷYE��M�/���×3��>|h  �cǎU,SRR�  luuuv%ô���q      �`3E��/������5g��F���x�w�ܭit7�LK��}��u=q�D���3�L�lՑ�*�9���Hk����ы�;�@�Ѱ:��T{�Vu��;��o����D�
���/�K�1�T4K��+�x�R�o�>   ��$�	��  �9)r��1��Hnn����       ��f�}�L{��=���=����{ϞW\�p���������Y���***���6av�j�)�9��+��\/߬�4�"���d��9C�N��]�Lx�u��v�-��nQǱ�m�|$�Ǣ
֔�Ѵ�7��݁,xL�\��?����,5  �L���r)%%E  p7��&L �      `��B����؟���)S�'�|>;8���&͞=[�����t��effȹb3�z�ݬ(>3�E���$������1E��N#�N܁$�X��ݯ�P{K�VR���5�e���0�?SJٰ{�ݷ���&	   '���:;;��  C��ѣ
�7n�6o�,       L5���>��MS���Ne�MCwEE���}M�<Y�&MF�X,f/V�;wn���M�)[���=e��e����W��1�Hk�Q��;0�u��Rӻ/v��ئv���=�;s����=ey��i(�PH�HD�p؎�����o�Q���ǆ�M�{���)s�-�f�  �hV\\�����e 
������       �X�SU/���M{�9���3y0t7m�6l�رc5c�a�hmm������]?~�w�+��m*��$�S)l���)����L<���M[��m�Q����;�$��*s�9##C����ksk~���~���0A����jn[ZZ���h�&7�f�t�_d@���jٹ���O}I���(c���Zz��
�p  F���"{k>� 0T��@MM���      ��T��)����ؿ`��ܙ��~��{ZZ�-Zd�������}�ؔ���a]]�)�W,��=�%��+4�L��7{�0�p�	��^��S����>?p����t{E�	;����Bj7��`Z�͇3>�9�m��愷�j��������:�������3�y�'4����M  �h���7`��  8����*o.�K�hT       0j6|�}YYY�8q�p�zV���� �׫%K��[_&{w��!͚5���dO��2�	m�J�poo�7�Hr8�х�;0�B��l��~�O�y|�=�i[�0a�JJJ�0�>,h>TL������s���7'��;�Ç������5��竳b�:�?l�=0e�rV<���n�ӛ,  �D��x����� ���v)T����v       h��j�1Owr6	Ɣ��7o�Ŧ��=�SCC����\��_L�ݼ���Oٿ|΄���;��>�<��n ��x��M�I<tQeI�c'�d{�$�$���u��ɮ�Y?�>�Lfv&�d��Nf���8�oǶNK�(Q$��&A�qߍ��oy��ţ�����<%P�nT�Bu���_���G\�N^J'J���nJw`L�|Y}���F�~�9 �1Y���;�p��K�|+��ߓ-�=��36::�'N8���ǝ��a�&O�t�_�U5?�Sj�c�^r�   ��u�ɂ�:� PZ��{$q:�p      �}O.c̺[	��M�ȑ#�5`�<�v�����{��Ҭ���������k��8�n��%��;�#6�h�_�Z����"='n�s�`Æ����ի�@x�kll�����,ƪ�=zT���ӧ��*7�~�/|�Y���������/��  ���v�"�} `����)�9� ��4���u�r��]g���L&    �1��S;�����K�@@p����b٭��q�]��)ȅ�155�����������px��������j[��Ԩ�NI��.��S�W-������wO?�s�"�7�y���Ӗ-[�`{gg�볪
������W(rf8p@�v��ވ�ӯ8K�>�y��5�m�w�k  P��т��`P  �5�i�ʕ ���%���7T��(������>��O	    pc���o?
����-x����
�Z��ĉZ�d	ׅ�������nO�����3�֮�CO?������R:�t
����A��Ht�[���]���J'�7�9V�|ӦM�bmrJ=�>����w�}�b�v��k�.����T���Ӆ/}R=_�-�?�Kj���*���)  (<6S�����F @������       ϥ1����q�\Y�ix��QZ�mllL�<��u����V"�ХK���n�����ݛ�Q~E'�i�!�Dh��{�!��,�sBW����O��V�d�-�o3��J��?�� ��i�q3����Iz�����/;3�JbrX=������hގOh��>���f  
�WVV
 �|aw       �����Tbb0c|͚5B�8�I��8�K-��vqܸ˗/k�N��-eeejmm͸��=w���
.�G^J�F�֔�#_Y*�.������K�/��
����i۶mz��U__/ܾ��:=�������������Ty��T4�+���=��{��Z����  @A��� ��.l[u��m      ����Wc�Z�`�0w���v���F�R�H�ܲ�r_�t���߯k����?�QypO�SJ�������{�d\��{3��f�����S<�z��[돷���ںu+��=�b�
g�Ї>�W_}�i�322r��IE&�����B~��kގ_��<(  �|���@� �W��v8v&��Hw5       �Y��+?�LƸUo��|�ܳ*�f���N1�͛7���Vȝ��-Z���*�f��ӑHd����~������ט�{i!�����Vl�*����Z�Ă�����z���J�\��d���{��O�>+
�WUU�L(x��ަ�_]�>��.^�x��IL��W>���L�?��j��  �� dm��| �|166�P(D�      �g_�������V����{��v��s�=jii�gU��:}gg���7o�Ο??cl�]k���]�y\^JN�I�>%��;�֏���N���R�µ��c��8�C����+|��u�g3-������9�c�Xk����Y�?�o}�[:{��u?�����^���vu~�U�x�   �E{{�R���3� �]vgppP���       /��rƘ�;����SEE��tuui�����;���!x����Nw+��lw+ ܙ��y+��)��_N��R�ia���AE�� h��@�*筴���}]�>]�ʯ��$)���yv�� �;��N��	�e�ڵ�r��	}���֙3g����c/��oܫ��?�E�m*9  so����X 䥡�!�}
       ��=�����˗/�������۫S�Niɒ%Z�b���D"���~-X���u�A���k|||������W��^^�*���;�Nb|@ѡ���_|�ʛ���J�4��˺���C�ɡ�>Ղ�����O�o6����կ~U/^����֨���ix�?j��AM��+  �������L{  �2<<��J..      p�Ȟ�f_�t�P8��WCC�FGG����;�>7l�@�/Xw7��^�k�kV���^�%ݱC^�iy�<��pG^�
��K�>�"�F�ꆜ}M��:�g?�P�k�}��$}�ЪU���b�>�����^ӷ��-���l�#=:��S�C?�Ο�C�յ
  `.جxk� @�QY�      �od��3�,lk��P��J�t��q�������;��3��~�n�߹�g����lI�G��?ݑ�L8��c)v�iBް����_�V�µ�����i�=�G����Q*��iv���'�e�f�0{���~mڴIO?����b�Y�?��o4v�u~�sjy��  ȵ��*� ��dܹF      �m�-�ݓ1���)���&���/�섥-�z�,W�\q5�n�K]]�&&&f��5?��)�+��t:�ddR�*&�;����aE�.��sө�"�]�Zx�g�pb����ŧ4~�Y�co��>�����w�v������'~�'�m�6}��_w��ۛb66)��~Z�{��%O���j�  �+vj�.  �����4       ܪ�=_u��^k���B񨩩q>�ٳG�T�)Xzu�Ʈ���qW�/���d�W�\����/������@�s.95��๛���<�`�2׿����.|�J��g}ΪU���X�-���X��_�������e������Q��{����F��  @.Xw*  �Q(��Ԕ       �M���9c�����C�)kÆjmmn�M���w5���ܬs�����Ұ��'���\�#��9����?{KU���{ X���6w��xD��h�>�s***���;v��v�X�v�~�7SO?������*�Lf}^t�['��۴�=��������  �Ruu5� ykttԹ��F       �˲]��^���� �U�,�gKWW�^�u�u�]�뎛����j�ݪ�g���:�ay+	�����E��;�Ua����>Τny���WT�_Y{[_K������td��X��#���Z�łc6��f��_��.]���y�dB=_�-MI+~��U^��P  ����:.� �;�������       �vM�~�ɛ]k�Bi(++s*�[P��ɓZ�x�V�^-��j�RsKSS��z�ٝ+��+gUѶ\^��i*6%�F(^�1'��"���N%u;��Uή\�V�����#{���?Jɩ����,�|�z��	����N}�3��7��M=�쳳v�8���}�^���?�v��  p���wf� ����;w       n?�|����2|���������?�ޭp)پ�f��,Y����ܛ��Us���M22I���pG�Y�=���T�vC*St�*筺����_�5�?��f}�����G?�L?��f>�䓺�{������������e��O�j��A��<%   7Y�v;/  _�������f      �V22����c*:��
ߩ�ҩ���$_��e�����5
�䯪SYM�|~����e�Y%j:�t��H$��/:EW��n!;����-�꼼�����ƻ4r+�Vl�;k��ۑO8���{��m��?����d}�fs=��cz���GpY-_�\���g��/}I{�����T<��?�w
u�U������L  �'��~���=�F��i2v�Ϸ�;f  ���7��4]_��}��Si��o	      *�R|�O��+�O)����'Ĕ�zfr�_�}>�U7���]M���ܵ,�VrjTSݯg�ϟ?_��p�ٹs��{˖-
��L�pX�Pȵnᖭ�u�:߬�&�������/�p/~$w�S��KJL�y���X��r����ϋt������e}��O=��֭['�z*++�
��V��?��?:����O�9����5��5
 @��=�J.�����*�w#>�ehh� �gp�٢��fE���<�Np ̩x<�t���,   ����8��h�҉��0�V"4�,�ޓ*�iVE��7-�L�8��ҩd�8w\�jp{���N�k���N�0����!��!#�zy�~p�*ږ�+�DL�dB� 1�b�+��IL*>���6b�䯨���2�㓧_ՙ?x�_GGG�>������U��ھ}�S���_����%��c?����M����u
  �vXE\*� ����]�  ��n�ۍd�   ��I�'�=�Tlw��yaz���ag	\9��U�hY�TyG~u��:���& ��F�9�T-_�~=���222��N��kV����'c�r�R�M*V ��b�]&�D2<���Ϸ�N���R��;������{��ӟ��5��%��G>Bk�{����������u�С��	_:����V��wUݹA   ���Y	� �Uk��      n�U���R����i���Y$caM]<��@��;֫��"�� ��ZƘMniip=���ݭÇk͚5Z�h�J���	�n��
�ٴ���'o���فJ�Ŋ�;<�N�����f*q*��xcl��/��_�R�V5v�����v��!�vTVV: ��կ�������e��퇵�_U���  p+,�NU\ @>��8L�     ��HL(t�����J*�d�.U4w��㮌B�ȡtZ�������/����ľr�N�8�ŋk���*E��*�nU��	V�-�y�^P�<�������ޚ>:��d"��ML��?֧�y����ѥ���\��O=����nn�١�����/}�K�l�kYG�S��.���ߩi��  �[��������+�������9�` �g�T*��������h�V�     �ͱK7��S�����Ӝ��bC��z�&��<��br8c���V���ѩb��Ϫ��]6l(���n�MmmmF�}i{��EC�k���F"��_R229'ێOo��;�E���ì�ی����Z�d� �����	���MNf�Xg��?����o���~F   U��y���o��� Uq y����c     @�I��:����7�}�<�S5��UY}��[��{��755	����c��?pڛ6m*�{���㮮���NCCC3�:::�8إ���
��F��I�F�������j�b��������O~�xj����ԧ>����o�&�J���?oS���O  �F���;U� �g�Qr      ��t2�P�n'k��,�oA���
6/rg�����V�p��5;w�t�h[�=����a��q羳l���l�@u�W	ypO�SJǣ���U���vЈ����>�y��=��Z�l�~��_�d�y�*��ʯ�Jփ*�6�L��OZ������ӓ�x:�P�����ߙ�ZyJ   7���B  �H$"      �z҉�&ϼ�dxB�.�N+|�|>�*�:����:NaS�������w�^'�}�����^�ʊ�������?�k5�G�u_�T2� ��D��K�8�T������޹���͊+����O��O��U�V����*++���Ą��ۧ�{LO?����3�8�����U�塟  �[��  �;�      ��t*�TE/�p��VQ��������E.g��^�M���r��1MMMi���jk+��w7�V��~/�Č�@��cVe�P|HE�u����Ss�����D;������'��m�\k�\Oj���]�v9�w���y�;ߩ�}�{������tJ����WT�i˓  �*� 
A4      0�������
�۫����"T�T,�����q��X%}�K�3�}�ܹs:x�֬Y�ŋ�XX�V7UWW;��7�_��	y+��	ŉ�;\��L*>֧�0��_��q=����YK��|�3:t�3�
�������ۛѢƂh�z׻���_===�g������j��[T�v�   fC� P�ɹ��     ��<���*�xL:!���ވ\9����e��\����>gEMO�:���N�Z�J�.
����������ymJN�(P���l*A��bE��>���Ϲ0��7uu�z�]�ٛ˝w�����d�� �088��_��]n��:	����3�<�K�.e<��Gt��߭5�}A5�6   �`0(  ��_      �Mrj\���T�R����qD՝o�{�goll�k�5��=q���jkkӺu�
���]÷N�n�{�
��jnnV��eO�Tp/^����E�⹟3yj��N�һ>�����n76Kh���:v��O��?��v�ڥ����!j!����s�=���3�(%#:��?����NU�_-  �k��  �.�      �)��K��TJ���RM�TV�*�/�6�8w̵���b1���NflӦM
`7���V�=�z�gR�>�{g.2��RpE2<���`η�9��_���������v��7��W������#k�l�f����ڿ�"�Ȭ�gco�O<�r?w�\����'���[��G  �P�U   ��.�      o��dhD����k���(��Ň�绬jv__�*++U^^.`�\͌�ܹ��)nٲ���q[�ݪ���~��I�kR�I'���II>��ņ�;n[:�Pt�\η�Qծ/�?�o3B����Ndf��t�RMLLhllL�����r���l��ޜߊ�?���y�]�p!�q��z�߯5�yN��
  \e��  �w�_     ��ҩ�"WN�ؤ"!ņ.��m��.���Ͳe˜§SSSڷo�S�V�;����ٻw����*�[��|�][׬����wcV�uŇ�;n[|��f��P*6����Q��Og��+**�p{Y�컷���I�UߎFiQ�744��7������j������zzz2�8�/:�W��_�s  \eE  �w�     �f��J'���_��*Z;� �X�
�UUUoi��mۜ{g�籰nmm���b��-G�u&`lذA����W�HĵuY7�¥R��eI��[6��'�ņ�;nK*R|b0�M�5����>�N���,Ծ~��j�aT�:t(�
\�ڪ���+�	HSS����vǎ���gd<>��_�r�����S   &�L
        �`�R���U�J�#�_V�e����pf�l�ˁmݺU�t�ɂ���^�\�}Ҋ�vww���Z�f�/ο��Ł�8���*�'�Xw�u�'ѡ9�����޿L,�1nU���f��(kb-k����������m�����������ojll,��_���;7�~�  `�& �X�      ���{���W)8��pwQ*V"4�1~��۸q�t?r䈮\����sŮ��>��קS�N9!�իW+_X��~_�w����eiy��{q"��[�W*:��m��v���^�_��]�b����oz�.����&��ŋ����ƛ�8q��:�Ր��L�!�R�����O�UѴH  ��%�� ��     pU|���]rjT����U�P,%��A� �n�@��uׯ_�,VAۊ�Z�ǭ/p�l߳}pbbB�?��Z[[��s���[��B�[sCYYf$����d����{M��^��㖤�q�G��t���Zp����g�M�cR�����X�r�r�B����={��
[r��#���з����Zb|@]��7��?�/P.  P�� 
���;      ��1'�P
�#�UUu�p��ᱬ�5557��e˖9�Us?~��jkk�ˣ��ޗ^z�ٟ7o�<�����kw��~����1�P��A�I%��C��$6tQ�\��{�꧟z2�!/_���Vook׮Ձ��d2�����y���Mo�����:���l��N]���j�W  �tq�
 (TC     ��J��,���Qb��ݐ�r'�~�O�exxX�r�����ܱܣy�嗝It�9�:,��lܭ�B�°��t���ň�;n�ͦI�Fr�͑����޵-� n3~,���Ӫ�*�Y�FG�J������o�8̵�K�jӦMڻwo�c���=ծz@M��'  P�J�"0 ��p     �IL�T$�ƕN��+�nObj4���ܯjnn����555�}��9�1ݪ^܊�����,ln�1�犛�l�������R�
�E��;nZl�RN�7սO�����sƸ�\X =[[�[e'0�/�ŋ����ӣcǎ9��%�~ս����={����iu�)�,ߢ�� �ғJ�        P�C*���wX���3[w+b���jm۶M�X�`qmm���b-l�B�6c���jkk�|�nv�p���*�����?/F�qS�,������q5�������xlɒ%jllt}�V9{rrR##��R�ܲ�x����l7��GyD���N��͒S�N�}Ϳ�f{  �7/2  ��l�H     Pb�)��!��ddB�"�~�,7����P����t:(:t����[�L����r544�ܹs:x�V�^�Q�M^Wp7�TL��zQ�.n��A >ړ�M���}�����xG�w���2�����F��b'�{��qޘm?�wv²c�}�k_sf�����g5��_��я
  ��k�  �G�     ���J.w���V��+�D�ܖei�����q�F��'O�ԥK�<)�
�(�|n�[���u��i'/i�F���=|���/��o%�FS"�˄�W*��������[�d�����v��yX��N�/^�3g���ԩS���q����f��lV��?��>�_�5������V
  x���;<��M=�Z� ��n>�����4�     r)�T�I�J�{�B:����W�7�l�-������r��^fՀ�}�����I���jii����]���f�}��)�N����{��wܐt*��Xoζ��i��N��}��\�R�`���B!�������Ӯ�f�Y���X�j3D�,����������Nh �B��U����m��d+���q�BF��  ����uy�*=~ϵ�{D      ȕt���Ҧ��={b��j.�W-[��Y._��cǎ������j���>�H$��K/���F�6m��}2'���qo��}�D�7���͊�B�_�TO>������v���y��p8�#G�8o(l�HD�v�r� X���=��C���������S;5������O  ����1 �     �t2��S�߳f˪y�2�E�9���:���e��V}}��q�Ν����͛o�����gS�{Z���{q"���d'��m/t�����N(���`���n��v�1����t��>11Q�۳���o����o|#����?|VM�߯�  ��*�'��9�� ����a)      �t����SW*.�T����Φ��Y۷o��Ԕ����t\��+%pV�ݼ�����NE������w������ip/F������0�-�RG��Z�л3[�r��3�즫Un'�^غ��t��9566���ZŦ��U7n����g�'����_��_� ��g'��Ymm�  �GN�<      �8_	�����.��V,��m�6瞝ex�Z(��0�l��-G�u�#�[�N���7���(��"�[@��7}���]���]_�S?�=c�f�Y��+V������x-`����	��@�p{1��v/^������W�V��<���  pOzxPi�'Υ#7wj�&''�P �[v!����ĢJ�^��R�{S     ��|��߻�����s��W��b�[�nu��C�ihhH�퓶�?��'W�^�����~���I9��~&=�����|^����V�=��VA��z�uR���3���V�Z��O�:��Qx,��ꫯ:���w��͚{��ަ���'���cZ���W  p��o~��m�T)����N�>
� @���{2ys��5���      ��/Pz�R����f/@u��s��7nt�m�{zz����\�|YSS����u��iutth͚5�>�-�Y��$���B猢Ļ)fg����s�9��/k��y{Ƹ� ��W.\���Qx<���1��Ԩ�XG�;��9)~�H�i�~�j��?#  Pܬ�  ���)��     �<_E�J�����g/����@V3��u�]���ݭ��.566�Z!����>h���{�9����͛g����?g�{|��
�ŉ�;f��R:������zrSg�l���j-Z�ȳ�Z�v���\�|Y'N�p�|K1�~Ֆ-[���k�mW������S*o�'  P��� �gp      �Z��@e�}�^�g���FU�-[�,���:v옓q*+#���c�͋/�������}��
�uXH{>�I$ň#&�K���ͶRI-���V�����V�X���H$��ǏO�^���[��ǵg�g&���K���^xa�x22�+������	  �p8,  �Ummm^�
     @n�+*���N�ε��*����+���J������;�b=p��S���\�\ihhp>���+N��C��k랭�{����"]�wd��)���d[�����~xS�xkk�g!f;�Z�=�H��^�ݻw;��ϴr�Jg����|����D�v����V
  ���	 ����MT     @��)PU�DhD�"PC���M(���U�yھ}�ӥy�޽N����Z�\����������k���Zg�<�e�R�J�W'>��k�!��������P*�5�cjk{lưUm_�d�g�={��&''��w��Q���N�Ϊ��ߘ1�N�u�C+>�w  ��Α켙�D �|TUUE�      ���֒	���e*�&���o����R!�P�#�<�X,�Tt�����+��Y�}ll��/���oy�E<��u�����}Tp/Jܑ!�*�M5ȩ��юm[2ƭ-�W3�FFFt��!����8�ɛ�������v-[�L���3Ƈ_��{ǯ�v��  ŧ����;  /Y�ۭ�     ����{O�j�,i)ܾ������RԴ��B[�nu��:tHCCCjhh�kW��۵}��n]���U__�,7#[���Q*=���B#^Ud�U��t"��s���g�uvvz�M�!t��)!�,�W_}�	�[�7�Nxϟ?�T*����'�=_�Z���  (>6! �|dE�Ui     @i*�i���B�DLŮ�a�������9�
Zmܸ���ɓ'u��%56� �sm��'-��Fu��e�������|5U�u�@��U�L��C9�T�������,pf�y�������f#�ٳǹ�I�ͳ��W�։'f����B�{U�l�  @q���p*Tx�� �[e���7      ���TִP��s*j>�ʛ���WT��Aɩ���R�=�5k�8Kww�����<�U��d��������-�nAw�t���:�ɖ����7"O���^�xU1CbbH�T2�i}������V����ÓM���9�3�Μ9�.8'e����}���$�Uܧ]����O��  @q�D"��-w @�����|�	      7/��Q����y���X�k��V�=�e˖9˕+Wt����׫���'�g����z��}�&]���g�|���M8��q�
�ŉW3�'r����g���M�V��F�7˪���6���A8p@MMMN���NfW�X�ӧO���5�/QU�: ��a�R�� (<6�*[R   ����^�3   ��UVӬD�x�Sۖ�*k�'�����R�S��і��Q'ce!c���������u��b��t�	�_�|a�k��H��}�
�ŉWoH������鳪�zhư��Y�h�'���-v E~�V$����s!���p�=���Tķ�7L���w~W����)  P<����Ȉ  �7V�=��A�@  
���mkk   P�*����T���ZUVC�m��e�<��p8�,UUU*���ھ}�����o�>g���x�f�W]-b<44��imm�5�9��>�L���D�oHL�d;�3/�ѭ�3��ϟ��3��70�����>]<xPN57��Nh�,Y�s���~�+Z��o9'�  �xp 䣺�:ޣ      �����	�'BEv��g��Ղ���٫�[����C���V۶ms�����w:>[��V�j���@ �,cccN&0��$�qkxU�d�N����������-T�={V�{�������@��c�֭����	�?��Z���O  �xX�7kk?�{  sȪ�����     �MU�:M��ӭ��E*�i�Wپ"�x�ܯ���[�nu�:t��yX&�YVL�~�ߩ�ͤ*�%��?��P|�Ñ�L(��y�����~O��:kQ�E۔˗/;-i0w��ǵw�^���s"�#6Y����9y}�����=�䯠E  ���w�bA2�  ����3�
      �	T7��u���T|�2U/\+xc�
���BX7nt�}��Q��������qMMM��+�̟�R)�+�) ��ʃBq"�Grr8'�iܣ�{�g�/Z���mY+��/
s�fd�ڵ˩�F�=���.���?�1���=~�+j}�) ��`���B�  ��[[\      `6��PbbP�Ȥ
]��u�{[����e��~��a&�
�r��9�9s��kq�c��]�wK4�S�a���/#�^��CJ��y�6:5}RzO{�xmm�S��m�f=[�x���s^[̍�+W:������	� PD����
���  ��.��B!      �q��/ݤ�S��t*�BlY����;�����W2<>c����.]�,���:v�jjj����,��W[=[��P|�`Y!/Q��xq�Sc�'�I�7t�%m|�]�,p}S�pX}}}Bn]�|YǏwZ�n�[vbj!w;Q}���4y�Uծz@  ��Y����A� ��a�d2י      P�Uu�Z�^SJi�@u�*;�	����d����������ett�)VUQ�m�����ٵuY!�l�����q��
�ŋ�;����v�,��?Ƙ� jkks}[.\P:]�g�jbbB{��qnb[��a͚5w3�p �HX����_�֭�� ����Ȉ��     P�*�+�(r�
�?X���[��W����ܘp�.��nll��~F۷ow~f{����WUU����v���F���E��(S��xp/u�tF/D{��u�3�� �f�co���,De�v����� ��<��Ң����#{��%����WT  6;;��|>w ����"����'     ��U�_�t2�h�YE�jW�/9��s���XT�7���Zo{���Ŝ���pX���B�r�0��W����Ǩ�^����T44}���|;�O�P���6(n���w��Q8��ܞ� ��^�Z���ꌱddB#�S-|X  ��9s�	� 0�l�;�v      ܬ�Ew:���R_^
T֪f�}�S�:����p߰a�ps***�u�V�Z�C��6-=�`P�����/[�T*�PM���+c�Q�"�^�S��o$��چ�:6+��Y`6�lppP���|m_SS�nG~[�b�v�ڕ0z�K� (6�pbb�9� `.Y�$�6      ܬ�Ry��[*R����E5�7�(r��c���K��EPo��ڸ�G�N�8�����%Ī��YD-[��ohT��,/�˃�3ŉ�{�KN�y��ą}�pwf����v׷u��%�v����^s�SnGa��k޼y���1>~�Y��zU��~  �[�PH���Z�t�  �Kv�;      nU�y�ʪ:��R���o��j[���w��#�`�S�?|�Ȍ�s��	��;��~��=ڮ���~�x͟�^f�
�F"����ɴT��q�_A�bF�����Q��y�#ޥ��̀��rS<w�=p��
ٿ������^������t2��]�y?�I ��f���a� �9g7=FGs�-      E+PU��;V��b��GҚ+��U/��To�ܪ[�-#�>>>��#knn�a�m��ѱc�TSS��2"��h���+�9�k]�VJ5�?H���q�)a����ە�������zUVV���+W�d=P�֝:uJ�/_v^/��´l�2���+�l�7��� (�D�9gۼy3�� �9c�***x/���U���Jѯ_�T��o���	   ���9��`s��.Qr*�E|����W��m�D�P��!�?���O��}��'�˪{�222��*:�Qjkk�<�[f��z%��6fC��F������o#ݳ_w޻2c�������N��ԡC���kn��anXȠ��=����]������]  ��uuu9m	 �JSS������ ����F9��J��3�H�7   ��5�N���Ġ�WN*�t{>�*Z��}�|�A!Ԯޖu��������۝ �}��1���"�ܬ�n��ml��Ny=E�_Q%/�%,y���d���Ό�w[�9�.p{��v�ޭ@ ���Q<�,Y�Y�'��������  
[ww������  �3�8�
      p[Y]�ꦗ��b#���t2���}��nRys�*��(�O�m�*Z+6tqƸ�Ὢ�*=��CN>���Nx٪��0-Z�����}�k�����Y^��5���F��D�bS�'z	Ϸ��>3t^SS��L���^��X;���q��7�Ogg�3y�Z#��E� �"099�t4�Im  ��g��      �����YԱΩ��^�c*2��i,�/�P��ez]�*�o����L!�]���_��cV�qll�B�9bŶ�n��t������a�����][_"��Z��R�J���A��Ŏ�{�JF&=�F��Kw���w�z�Un�U�<{��s�A��xYР��N3��?�Lx�5  
��/^��e˖)�J	 �\*//w��
      �ϯ��vgq�RN�!���Q:�pK���K��_^!��GKYP(<�w=�p����c�������t�=�8�>y�.]�Dн@,^�X�@����V����^�~6��*��p/Q��[C�TYٞ1nA[7Y����LÄê��ݻW����`�k/s�ĉc�XX�G�W�?)  P��M\|�G @�ٵ���L&      ��/e���x5��NKV��r�G�%�>�֬Y�,W��Z5}�^���vG�l�p4�њ��Z �1��p/Q6c�kK�������2�����gmAv�����)-.�����p ���<�� s����	�S�       �W��z�zM]84c��v����s�:M�����&555N>�#j�|w+��B�����G�����l���G���G�N&<�F:6�;�g�[�p7ghMNN*7�ȑ#N��:��X�=���/
  ���a�Q{{�  ȥ����       �\����[�s��i����ܛ7o�����������TEE�0��.]��D�X,�,�:3Y%y�=�UT��ō�{	JE&=�F��I��ؖ1n��D��s��e���M0 �^�������ccc3Ƨ.VbbPeu�B�H���U2<�T4���Q��	�SI9ӈ���������N[�@U��Ս���"5>>�K�.9��� ���c��f       x�a�;t�ۿ�1nAj���r��>��S���_w�_Zv	sgŊ��ϊ_˺)�լ���d K���y_Q�-�g����n�j���Ąv������٣0Y�k���8񒚶<)�t"��h��c�JN+����i�O����'���x����U����]��r ��]@�pႶl٢d2)  r���ՙD��       ^�]���j���,�a�����B����Ҷmۜk����w*�S�5��kss����Bc��F���"�p/�KP*6��6U�윙wk5b-G�b�H$"d�o{��qN���,�~�����c/p�S��AE����N�v����u�9�.Qy}�*ۖ)P�" @a���ֵ���p ���:�C       x�(W��j��9c܊�^�xQ�/�Syy��n��\K>t萆����� ��ʕ+]]�ݏ�p?����9e�P��� �+���Q-k����w��5<<,d��roo�������LQ�/@���VrjԻ��R���:KYm���W���M ����ӣ�����=  7��ڜ�      �B�����}��p/ �t�ƍοO�<�K�.Q��c6�`�ҥ��Ӻ�g�/p��!�������E��%���锷�}'�p㼌q�޲��PSS��?kk�c'���3C���ǔ�L2�-��S��tX��n719�ę�T�0OUw�_Q- @�WWW�����;  ^�N}555��*       ȅ��WY}[F�b�޽z�����Q֬Y�,����=N��nݪ�U�V9!w7�}�k��2�ɚ{�@��RA���$cS�o�5=4}��yq3t�H$411!H�pX�v�rn([��k�|�rg��锦�P�m�I�8�H�I���+V9>11���kUѺĦ�
 P8��.�lڴ��; �s�����X,&       �_�LM��G/�Ō���~'(m��e˖9K__��=����ʈ���&|�$7�}�P(�1~t�\j�>gTV� ��%&���{[`r��3��6���ֽ��V}��[_�����555E�v�%����iǎz��3��B�^'�>G҉��.�W|�_��:}L]:��䀪�-_���8 ޱ��cǔLz۵	  cw�>ä*       ��|��2�Ɗ�p/\���s���1'UQQ!ܺ�K�:�d9�k��v��b�jy�&����~?�_�KL:�|�3ojVWW������J�U�<w���-0�h4��|��7N��,Y�����ׅ�KFC
�y-'�nV|�O��U��~*� (�x�/^\�B �	jkks&�      @.����*Z:�0c|Ϟ=�Ї>D����Р�۷+���_w�y���y��\�v������:�7�H�y-`��}�W�G~�H^bR��OO���%�R�۳����U������il�������ĦM����4㱅���\�x|���ٽBn%��4յ[�DT�*	i��˪]q��t� �B022�ӧO;�ڨ� �JKK�r�D���       |~�>�s���o�����͛��WUU�m۶9�}��9����:��,Z�H��ͮ��^�l�o�O5J9xi�5<�  ��IDAT�B� �^J�i�1O7�9��E�����Z��B:�PH��*p�޽۹q|mX���ږ-[6�ɺ�Gvc] �,�{ʩ"�`�c.$��:��ҩ��]:��WU��!�+�;� �aݎ,�c��  �X�X�H���4       �O�#O���IJ�f����K܋�����J�t��a�H�Uy��z��\_o���X\�w�k�=�(�YJ���t2�Tu�Rcbp��U�nVp�������'V�ݾg������`0��{�yC��l�t*�ȕS�^r��TtJ�]�"�~���L�٥��2	 �]�9{��sq�sH �W,�n�Z�}       r-ضT�w=��#��?u�zzz�p�B����~mܸ���ɓ'u��E���b��ŮWo��f������J4x_��_Y'�? ��%$��z���2kK�p�v!nW)�7`{#�7a�I���799�|����ϟ�uܪ�p���'�v9U�M:q��uk� �ut���]�!x p�UƩ��,�k4       �Sۣ��p7?���S?�SB�Z�f���?��nm׭- 覆[��l]]��;�eՍBi!�^B���+2`�@@�m#
�����{�����fxK�rǂkW[�ߨd�
��V��a��{�JE&�pP�K�  Y��̙3���{	� \w��Q,       ̕�M�Uy�<���f����z�{���@q[�d������ȑ#���UYYi�bW�\��F������cݽ��l�>Cd��@Y�RSڿ��?{w�]���=��%˒m����J;qH(�Jvi���vwۅ��v���?-eۅ�YnXh d'��H�N;����۲�C�}��_�ojcy���H�y=����(���o~�����o�IG�{I��{2��M��-x�u�V����(.����
�-[v]��%���R�[hm�xg?���R��Z Ʀ��^�ݻ�p;  %lU0;���       ����r�gt��2b���O���/�a�!;X9��,S�c�W�
��m�@J���wʮA_lWw�T�Q��r
��w�6��g��7�Ǣ*�����&m�H$�r�{�7����Zہ˱��2�����̴�UVV�hG����:��~�5�S����B�^�V�  $י3g\�����	� ��&���婧�ǅ�      `4U��5>�7���,M}�g\�&�ۼ����^�n��X����<v2�c��^Hl�����:{�T��\���/�{�,J�ё�3*��D2�z�������A{��QII	�v\���:;;�j�*$�Q����.����='v+ɜv�Xd��s''�'  9Z[[ݱ�Y�� ��V3�X@       `��痪���������mmmھ}�n��f!�X�{͚5n%��^{��

����={v�w``���.��ɘ"E�o��x}��	ه�{�ES������ō�rɒ)w��u�V7;�B��崴�hΜ9Z�bER�Z�/�u�(:�'o yS0���ݪ��e���
UԹe�  c���ۻw��� �,������+�      �h�p��������F�oڴɕIZ$��5��\������뮉���X��~�D�������ko_��(|�Ŗr��,����|%n�
��7K���O���m��.g��0ܸ��v���kÆ)y���҄�m�
UL�'s��c�?�!���$ ��c'il2ۡC�\�{$  7v������q'�      `���g�x����c#�O�<�;v覛�5d;�׫%K�����߯����
�O�6�|AM2Y{{GGG����z))W:�ʄ�D�=[�b�ESh����7>�N��m,:~������R�v``��kצ��b�pO�Ho�;�(SY3}�o���< ƞ�g�jϞ=n5� �U[[�>f�
{       2�����j����]���ҥKiq�y�g�v7��8p���, ?^Y>3U�8��E�?�X����S$���g�X$��F�(q�=&m�6�Xk�]�\[���b-�---ni�t������H���cVt���v����5s {��b�޽n!  n�]��8q���&f      �X�7u���Km;7�ohhЫ����˗���ɓ�����ڽ{��������H�e�����VF���7��d��s*����lc���m�u�E�R���_�L�N<5�۟u۶m
.�\Nkk�f̘�+V�m��g�pO�XTm�t��'�8WLv���&�Y����iq ܐ��J�c���       cM�o�w��z"�����w�㹥�SUU�n�ޱc�+�������I�4mڴ�<��^������Q:X�?�\�^ܳD,���{�'~nO��.�!��;::���+�r�����;�3�����O8>�~ZH���e~cnl�OC]M
pP	 c�ܭq`���� ׭���}���       �E�u7�x�j{�g#��y�f�v�m.���H�֭Soo�k���bc:�g��o�9%�m�������G:�[��Vu_^�<>"�ٌ�,���{n 7������!��1�9rDG�Uqq���rl���ޭ^�����jp��v
�1�yV�b��w �l������ck���� �����X��/�       �S���Lm;�kq��G�b�
WD	\NNN�֬Y�򊯽��+~�T�j�X��U�R�4oד����hwp��%P�� =�.��"�����p n,�����ۂl��m۶���ԅہK� [�f�ҥ��2�.���#��,C��C�M �M�hԵ�[�}���D  ע��F>��M���       �r떪��y�G�wvvjӦMz�{�#�jX�q�ʕ��o����f��>̙3ǝ�O���w=�b/�կ��J��7�;|���,S�[���-�v�3Y�b��L/����9���\�M��<y��/_���R3��ܓ":ا�@���5��"��� �=p߹s�/^,� �ke�eM��H      `�����Q��G�1���O��nSII���e�d�uVc�b����Z�[^^�%K��䱭���)�䲣�O�)]��	�cl#��-b��<�l�,c����7�t����)�����u� �㎤�N�(�3�-��q�o�@L��.��x cQ[[��9��v���] �ղ׍s�4      ��.XZ�	��wjx�#���O~�}�p=fϞ�nڷo����Z|%�pXk׮M�6O�:��Z��AE�
�V�I���{���>��(�����!��r��I��dx	��r����C��z�rss5Y�{O��٪�>����R���p���NBؒy��~�z� ��v����;��P�        �P�����_~W�'F���ꫮ�t����ĉ��
rw�ޭ`0(�?�q\���V ���I��wvv��+>�t�t���S��*�رS"��C�=[��ddP~�'n8�mգ±��m�TPP0�K�`|� ٢E�4a��evpuq�=:�+ܸh��M�/�B� 0��l�]�v�Ue��!E ����x;Aolu2       /��\ռ�����?w߃>�Z����QZZ�B����ڱc�KU }��媪�J�c[��]O��e6�k�T�<=Qc��'A� C�=KĔ��J,qAًYp&i�� ��_z�%���[��kl�P��e�4�z�`6�E�mbC� �]v���Ԥ����v��  �S[[��7ڹ[�       Ɠ���������n1~��=��S���{$C^^�֬Y���>m߾�������s��q�xS��퉮�|�I]�w+]��.����"����|�ݱ�F�ݖ9{��km.�\��ڵk��rA�%s
F��?Y'JP ƺӧO��^Ӽy�� �h����c�%I      `��x5��o���/Ql��]O<�-Z�)S�H�p8��u|�����Ң���zL[i5�e�����,�b]��ڙ�R���}�V
8��{�Hm8�2���GS������ٳG%%%��qY�����+W&u�]�$���j	�&ɾ�`4BP �:k�8r�Z[[ݱK:�� �KYY�����8       �Qx�U�����G��u��}�{���?�����e�/^��¶5�_O���T�x�;RVb:88���Ƅ�={¯��2����B�f��$�%v��Ѻ~#��{�֭���u�v�rl��-��b�
q��� `�MMMڱc�n��v �D�M��>�����T      `������Z_��z�����דO>�{�G@*X���ev;|���=������X ޮ������Z�ӊ�]�s�IomP�X{{��J���g�Ԇ-�n;�T�L���M�cی�m۶����[��&@lؐ��T!��:o���z� �>kصk�֭[玱iq \,//O��o/j�      `<�B���i�_��v��p���I�&	H��ӧ�ۉ'�w�^t���Vл~�z�����c�h===q�=�}z��N]^�b��Jy|�0R���U�C�����lpOU�СC:~�����R���g�v���[3�b�:.����T��%s<,� �B[[�Ξ=�={6w @���:w�����      �LP0w�*���y���׿�u}�_P8�j6��n---z��7�:�m�C�����������<uh@UuJ�ק@!�툗}�,eK8��/���A�B���\�:�w�A�ܹ�5q[��}���j�ʕn�\&Ip��Swp�M<��{��	�n�(  �N�>�-[�h�ܹ�8;�S �M�>�Td'�       SL�ȗԹ��ֿ9b�̙3�����O@������x�kQ��ܘ5�WTT�4�h�:޷��U'*�P:����HWƳ"[����?��}2�^orB��<�u�V7������X�}ƌZ�b�2Q�&>/�����m|����`����ɓ'U__���jw  3y������
       2�7ִOO{��fņFff6o��ʡ25#��+77Wk֬qE�;v��޽{UUU�9s�$}[V|f׉]���Ӌ�R0�e����
VH��{�Hu�]�r��d��]\��v�R{{���a��:;;���-��I���hI���%���P�M�Ɵ �+��f+���K��>@� �X���i���n��        ���-U���L�?�|�}?��T[[�
��t��ޕ+W�����}ʔ)I݆�Yc|"���l��)PR#y����B�=[�a'0����X	�9rDG�Uqq1�v\������z�j�Ae2�Y�|���S���7���ח��� 0�Y{�������쎓	� ��M8v�www       2ф{���_J��^1��ק�}�k���?�\)�nVƺh�"��k���JF������������W���ȟ_*�R�g	�R�@��gM�9#��C_/��t�:::�}�v��p)6��^��,Y����X��Raܓ����bu�(�쀓� 0�tuu���M�����n� ����������G2��       �Xb���{P��p��G�g����w��O}ʝ7F����磅��ڮe!-�~=�K���9~�E��U��&	��������v�Xp8/��p����ˮ����H�崷����F˗/W6�T��_P&$�?�<k���r Ɵ�'O���֭[玷�� `|�%wϭzg'�       ��&h�g~���A���"�;v�g�ц�&�=zTӦMSAA��{Y�k(��Lf��.l9΋��詮��*����.p9ܳ�'�ވ/ḅͯ�}�b>����h/��o�����Ё����u�+ty���<}��{��ZH�@���:�l,�  ������&�m۶M��vw �b3f�pm�S;�       ��`�:�|�/T��w�O�SUVVj���F���-YQQ�j�f���Z�e�.�{���'ܹ���أo��[R�t�������{��x�p���R���y��ח�>ۑ�ݻW%%%��qY����ӣ�o�Y999�V��TN_N��@��Ne2^���< ��<��Р�۷k����!w �>&LPa���,�       ٢���A�G�����F��u�o|���?�c���	Mt����\���(meV��Y���GfD-�n�v�o&���6�*O�*�������'Ef#��%l�K��{�	���XoT��{gg��nݪ��"n.���M���wﳝ�]$B�{rJj�ݫL`V% �k�O�v�ؽ��Z�t)w �B�f�:����        #y<���7�W�[�#��{��׾�?��?%��Qe�p�����Zi�9j���ٛ��]��ʈm��_���ç���.��7��@A���A�=Kx|�����Xvo�x����joow��Nx۶mn��{��2-�ׯ�f��$(&��L��)�?}P�Ȑ2��P��F ���Nv466�W���[b�w �.��ra{��o      �l��)���������l?=�>+����G�䞬�W�z���j����7o^�}^��e���5��:uJ]]]	��l�~X=��O���lR	p5�g�wx��ށES����5��ܓ��ewc��Μ9����3����m�]����E��5��~"PX)$�M0
���ae�P���� 0�Y����V;w��M7�D� �����̙3��vһ��G       ��Bu���׾?_����s�����������B����b-��|�k���y���n71#�Ξ>m윩h~�����\-iY�B�����=~�7����dܭ���g�q��n.�B��B�jժ�Mt)Q�{��vx_���y�.T9Mg�)ͬw�?�Py�  �g��^xA�-�� �ą��v�v       �,o�rM��wu�>$]T${��}�k_�g?�Y���.1z�=���<�������u�ĉ��_���n(W_�$���T��F��`O�E\h5���P�"���yG.!a�7��5�O�v��D;f�Bl��+V��(��0SH>�?�p�,��ܣL�8�M� d;�QUU�;v��(� �٬�e֬Y翦�       ����������Oq��ݻW���w��\^�W�hٷo�[���N�<�cǎ%�~������V:[�!XQ'��'�Z�J�"���ά�;e�����QI�ȧUoo��?f,��R0t�v� K����t���ׯ.�&�$Z�&T5CH�`�4��+�ӡL��-R��V ��a�6��W����.]J�; d�I�&)??�}n����      �m�����N��Ͽw�+����k��_�kB�5���	�/v�G��*�X�������	�k4
+��Vܳ��L�6Z�c*�9600�v�׺4KGG����\����k!0�}�9�����;��� �JgΜI8Q���>�T���:�KŢQ�g6�2w�R�L ��bK�UVVj�����	;@���+�g����ο        ~m��~Y��^�}��q�mݺ�]G����	�c�X��ڭ���ѣ���'����;5�����5�I�,����j�����uaa�U=����݂�v����p��F�jmmՊ+��W��Y!��Z���k����r&-�/�/ @�ɩ�N���͛ݒv6y�&� 2�����/[j���q>	       ���Q�ǿ�Ho�Z^�Q��Vee"4�c4}��_Wyy�+/K�Ý:X1:�vk�U�Y����A�=�����iж17~5w��j�����"k"���:v옐����4m�4nǵ�T�=D�=�B�S�n�@�	�Gv���J �l'N�Є	�m�6�z뭮}"��/ ���ι���s,�       H��մOW��.���X����nR���'\q�.v���֦M�4q�DM�<y���b_�^/�p��U��p�ثf��4�Ǭѷ%n�JK���488�v�WRQQ!d/[6=''Gw�q����c���y�9
WpO��ɋ�j���Ɠ@q��5 �lv\��ب-[�hٲenU% d�Y�f���b�m"        1�/����}�����Sq��رC_��W���|F�pX@�Y��~��*��k���O��/|���{;P��P�vY�}���}�<�'
�ܳ�5�[ 8��������Fn�.�&b����=�j��Ɩ�H�ρ�ghh�=_V�^��1��9���67#�n��m�Pw�ƃ@A����� �������v'E֯_�VY�% �񭠠`D���       pe�@X3�ݣ:��>��m?���������;}�s�s�a�T���wa�={��onnַ��m7��#�ڞ����-���v@
�$����B����m��V�@L����L�@���m�5t��Yj�p�������R�SFv����K����R�q}}}	��$����S����}l��5��'(��Q;� ����<y�-�h�a%%%nyE ��6o޼��f:::��       W�rw�?�����'���w��?v�����Z���g]��lmmm��W��k�����������Q���*����Fp�2�@��)����fGξ��===���ՙ3g�X0x�;���
�Y���kjj�l�2!y�?�p��)K�4�z�[w����T�1�9;蜦����� ���'N��g�yF������D �삊�O1���        ���N}�[�tz�?��o%�r���`��r��	noii���T��'���EyOR��C�!X\-_N��d ��e����-��8;��Y��`{8v��7ʚ����'d���^�<Y�n��^���R��r���kO̙�P��
�ߩXdHc���W��E
�L  ;�%���ѣG5u�T� 0N�$��s�����M|       \�ǣ���<��Nm�R��}}}.���X��v���}�v}�;�q�p'4�����_���?u_Z�z_�^E�һB�/�@�bV/@�p�2��ةH����]]]*((H�6�û�,��Y,D��٩իW���ơC���<��rj�9:��T�M='^�P��Paa{���� �4a����?�'?�Iv�c6 ��2}����m?n�       ���Ѥ��
W�ֱo�~\���F��?������}�]c��e#���驧��di����O|Cek>��1�_��i�kܟ���/�P�4��${�,�MCX��W9��j�.�9vww'm��]^^�Z����4o�<7y�u�ȑ���i�������)��lmPO���ӻ�`X95�M	 8�N�رCNN�v�ءe˖�r����a�v��c��       �W��
�M����Ez�Ͻ���z뭷��OZeee����~���޽{/�=��R��7�`�ڸ���<K'����R���*\5��d��e���ۡ�b�k>����Uy���8�D��,��555�3��+**�~�z!��w&Q��`�Za��x(�QQI�Z�wꀢ�=)ݤM~�����)���
 �������U�=����
�.�� `�Y�p�|>�������        �Q��.��/�ҁ/�[�'��������'>�	͙3G��8p@���7���~��	UM׬�ѭ"p)��
E��5�լT
�Oq�z ��g�G�`X��%Ot�U�����QQQQR�1q�D�"���.�[��u��_hG�:t(�x��ۄ1��U��V���l?���zv��[�y�
V�m���_X" pi��^\\�_��뮻��5� �6+�I����       ɗ3i����-:���R���q�[�������|������BB���O<��7��/�`�:��7ɟ�UB��MY��嚬IH�Y��My���ƍ'3�^RR���w ���^|��}�ʕI{.���۷/n���)�-���*P\�n��u��Pg����车����/,>�,W��B_rV�  d>;�oll���۵l�2����Œ5�
 �t~�_s��=�uWW����       H>+�&���u���3�~����SOi�޽����UUU%����f}������/�M�����&}�KW���x���ކ��E�{���W��L@�p�Bn9�Φ�n�l�fx��<��<r&QwwwR�3e������`��3fhŊB�ف�$_,w��r�l0x�AJk��؁g��[Ѿ.E���w�������w�|�Ǩ~ya�����n� �~ǎs-��p�}������  cӼy����6)��       ���B����(o�r���O+:_Bk����/�B�Ї�z�jy<!�mٲE>�����.�=�p����JW}����F����?}(if�P��c�	H%�Y��O�6Z|j���$82�n��i�<y2�q�.����k����詯�O�}�;������	LP  ����?~���ڵK�/�����x ��QZZ�Ι����Ϊ       �&ek>���:������Ѹ�������}O/���+�����������?t�^/'\=[3��O��S�{[��B׶>�ڠ�������T"������E&{ɉ�n��Wď�����(9aL�`k�ej1��2�m�ѵgϞ��EK�-  ����ب	&hӦM�6m�


�� `���|Z�h������Z_        ɗ[�T��|���֧���C	�������?�s�s�=�뮻hs�VH�_�J=����W��_���Rjl�h��z�?k��\���@��,�R�P����-��8��r�����NZ��L�2E����0v؋pKK�V�X���alx�7�����ʟq�   ���:tHyyy.�����_~�ߵ� Ɔٳg�U�Ρ        F��rf��OԲ�':��Oi��5�{����v���ê��2׉'���H�����r�5��_U�-N���Smث�ൗ�y�>�'̔'�ܳ��ѓ��iO�����FF�2���r��d�8�1c�����`����:-_�\;��.сQ�⻙Q  �IGG�N�:�>_�p�f͚�h4�n ��e�̧N�z�k{/�$$       ]��>���+u��S�~��L}�_ԪU���~�N!s���������?�명6hꧾ�`IM��RUNW_�>�bW}���*\5C�`��t!՘�|�Կ Db:��S]x�x$Qoo�rss��{���j544��^�C����N���v�ڕ��hɻ  p��9�B�7nt+*�A�. =>�OK�,9���οX�       0���S4���������wņ������_֞={�[��[��[�a�s��ڲe�y�uvv^�{��x҇�J�w~��)�3YHݞ��g�^���s0T5��Re ��g)o(�ͪ��Y8��p_����q�v�5Ywc-��G�5�ٿ�P%��ɵs�θ1kn/Z�N  \+MZ��Mp|��g��w�K~���` E�g�������jw       0�X{v�{>��U�[��}u��L�������jӦM���{�l�2a�ٻw�z�!���_�{�߭�������_�h�;�^��,���*_N��t#����w<6�&�ۑ���V+�9#O,2b�f#UVV&m;������q��H���f���K$___�;`�X����`  �z������I�����Ν��S���+-� H���2�>�Ώ
       0���fh��lR�������cu6%����F}��_ל9s����ϭ����V�~��u���+~o��J��*_s��-X:Iс^E������u��ܳ�/�(���!��w�4%od�}``��n��pR���z5k�,�ڵKH���vM�8�فㄅ�JWD   7����*..֓O>�O~�
�X��` H�����s���>��}�      ���Ps��w����Z^��%�u߾}�˿�KW:����Wuuu��c�v�n���_��=^U���j��^A��s0T9M�'�*�讷���-ܳ�?�H:�����/Ӕ�Ƹq�ؚ�������ݻ544$�ƹ��u�ֹI�n�7��Ur�o
  �FX���ѣ���z��u��w��i��Y�p�[��6V�       �q���懪z�����w�:��%�w�޽�f����w�X�����z�'ܿ��ț�J���ʟy�F��P�r��N8_�C�c�,�	���E�S��c���gZ�4�7b���S���I�N(Ҵi����.�ۿתU����'�lH�;Q��]n  �u��)UTT��W_�̙35c��|>E" RkҤIn��slb���       _�gܬ��e�Z^yH������K~�o��ns������]���*�H�ӽ��k�쭷޺��'X6I5���o��kO+��|Jj4�R�/�����0&p�r��"EϤt=�Q�	iJp�Vk{�����([�����,ÝD���� ���Z�mۖ������  @�:tHK�.գ�>�O��nR��p\ �c������������       �S�JW}@�K߭SO�����u]������nUUU��;t�-���X�Nww��l٢���ꮆ?�T�������CWJ<�Jс^����g9_N�;Rp7{�*4%��.�&3�^PP�ɓ'�رc���Rqq���.a�ڼysܘ?�d�@�  $�M\=z��ko���G>�7� �|^�W7�t���_�ڳ��X       �7�����Ϫ\��:��?���_V������i��G?r��V�\�5kָ@�<�֋/��V����ǂ�����}���Bu��YΗS �ǫX,�Tzk�Dް�ё-�p���tf�e���:~�8u�����z�jJ��u��566ƍ������p�&�   ;�())q�o߾]˗/w�ˡ�! �k޼y**���6Ѩ��O       ���/(W���LU>�v����W���+y��������M�2��W�X���lb�2۶ms��W��y����f�ф{����>ܳ��+_n���[S���HTo��hY�ȋ��hT���#.�ި��BM�:UG����[����Y|�܎��f&Rq�  H���U�6m��VV�ɬv�i7 @rTWW�����בH�        2ӅA�SO���<����ͱc����Ԃ\�}ѢE
�¥�$��;wj�֭ڿ�5����Ty��r��ɟ_* 7��;��+Iy����T-�w+640b�.�&3�n.\���z� �UjiiѬY�܁2CWW�v��7�?{�rj   l9>[E�N�=��#����ݪ@�B+,�����s+�]�d��      @泠{��J�j��C���۰������l�m��B!r_�d��ϟO������8�wd��k]�:<a�*7|F�R� �@�p���E���FR���^���4�32���ݭ��~��,�9}�t� �K�����\mذA�,/��B���)  �T�U�N�<�>��ܱ湐; ��y�^�t�M��}:��׳      �����O���O�m�:��c����P,��m�6w��|�9s��[yUUU�����=zT{��q7����d<^-ܠ��������# �E�ng��-�PWK�7�z�Mȉo��̄	��-k4�eV����N�e���,;��,���_�"nܟ_����-  �T�Ք�����}uuu�䘅ܭ� p}l��W��}���       �R�����n���u��o�e���`Ǚ+���HD���s��������ٳ����˕),�~��	:t�������{]�,�U�;>�򵿧PE� �w8�����u�鶼�D;G���������K�p8�.������l��M&�ef���ɂd�t��*����  ia'��Đw>��ú����I0;޷�e �kc��&M�t�k{�Ғ��8       ��!�v�&��4�w�F�;�PӋ�Q�΍�E�������e��f
ݹ�S��۔)S������Ο777����.�n��G�qe�����x�T~�'T��7��&/��������o,�ڰ�`4�mm�zG�Ȁ�`�E���,�۳�d6�*Q�7�X��:�/_.d.;H{�g�ƽ��*7|F  `l��|�x<׾������ܧO��Z,�
���h�� ��SZZ�y������K       ��*^���6�qV�/�H��~����)hy��_��α���'��UVV��+�k��d�ț��t���:uJ�O�Vcc���믻��Bj/\p�JW~@%��+_n� �w�m��v�C]�)���H��;����5��E�d��y�^-[�L�?�����`[S�w���>��v�ڥ�������S��J  `l��{AA�:;;3*�n�%EEE��7�}�{���2���T���q�5.|?���}CM3       ���/�P�;���;Ψ��Gպ�au�yN���k~<+��۞={Fn��wŶv�����|w�ЮZ뻕`��n�h�
���yo[	�>��[WW�;'n7���_l��3� ~��`��̻]�+[���+^� ��8/PP���{�`T�:��4<2�n/L�TR������\n����>�|͚5	
���x��A�GU��G  c[0�Ȑ������ݻݱ��U�·� �vnҾ��?������io�       �o��JU����Ez�վ�I����:�|F��o�-�f�vo�f�h���V0g����<o8��7�DǕ�9T��B����777�dɒ�˗�%H�����-Z�	&�Ö:v�X�x�M�Q�Ĺ  c_&�ܭia߾}Z�d��y�UWWk��ɮ��Nv [�x�;Gr��.X1 �v       ��������q7�w��w�~F�{_HKI�h	UNS��5ʟ�F���P�j� �M�1�?�L-�)�NKϐv��4�?2�>88��.����pص�mٲE��.tWVVꮻ���ƍ�=M|��  ƏL�����&��s�ꡇ�<�~F��,  i֬YnՋْ��3       �f-�v������x�>������>�۩�`����NZ�ܺ��?�V�^�@q� ��1��[�ES���=5��Y���/~MMM***Jz#ٴi�\��ɓ'�iz{�nݿ������>;v��[o�7^��ʛ�R  `l[3إ�=�Rn��:C�v�___���Zr���\��!�	 �6q�Dp���       �T;x/�����XdP����װO�'w�w�c��=.o��6_��5���f(w�B�LY��ɋ��* �w������+�PWKʷ����-6��wk%+++K�6o��=�����3��F���}ժU*,,��=}���;<^M|ߟ	  �}������a�m���ۄ�����'�xB��{����g�4 ��JKK�dɒc6����v        ���(w�w������k�����?�Իr���c�8�HO��zچ?�):p��-���/���B��J���/�p��S\�=\9�� �pGAyZ�����ZXأX_�����f���%u{�pX�W����??�CB6	`Μ9Z�b���^|�E566ƍ����r'/  ΅ܿT>M��|7�i!w���߯�K�j�Ν*))њ5k\3q,C�� p=rss�|��+���v��       ��Ƃ��v%��v��u��*2<��������,��F�ql�o0�fM]���!��)�"�Ȁ{$q!���ʤoӖ��9s�8�񨣣�5�mذA@�6n�7nz���  �����#��27�n+6�޽[�/�/~�i�.�n��q�B��_�r��x�����E       �x��]�
�����#![ƣ��[i�ֶ�
ͯj���uĸ5�[�%
%}�˖-�ٳg��ڪ��-�v�m����Wo�p�Mz�X��R�z�  ���!���n:tH�g��c�=���|M�:�|�; d{��j�*�/���ۣѨ         �lCJ	��J5�ڠ�P��%]}���9A��#���9uꔦL���m�|>�]�VO>��k���b��W�X����9sF�>�lܸ?�D5��o  �W6���X&����zH��{������M� ��^���o�/d��         [pGb���h9����h�ӂ�bF�F�����v���¤oӚ�֬Y��{n�������]��؃>��������o��  �o�r?~���WUU�?������6�D�9 �i-Z����c��E__�         �lE���/��`k�b��/�=��W=uzw�n�"#�N�>�B.ֺ�l����b�]�4�tuu��ҝw�) �;v��7ߌϩ�����  ��r?x�B�����������տrwC�@&�?�jkkG�������         @6#��K�x}�z��LZ�w�ݧ�U�U��q��9sƅ�Sa��.t���6�Y�b��ի]p	HĞ#�ޞȤ���<��  @�����������&�644�G������\	��Ds���ԩSG�n         D�W(��P�ٴ�fl/vM�GK;�mq_[[�����'}��G�V�r���----Z�x�*++\�O~����ƍ��x���S   ��{�ɓ�y!w���4K�,qa��\��{�����D �b�̙�1cƈ1�����h4���    ��   �	��<����e�lJ���v��D������بiӦ�orL&{̵k���?�y������USS�e˖	��}��i˖-q��"M��+  �˅��ї*23�n��{��qM�;w�T8ֆ�������;�LPWW�ٳg��P{SS�v     pM�^o�X���   d@�Du�(Kυ�m�y�5�\EC#C���x��)O�P(�;�Å�{{{�j===.��nݺ�o<���������~�������%���   cG���mU%��7o�<�����g�����d�ɓ'k��q���e��*U������'4�/Ǳ��Ai,��ti¼_�>ņ��C����):��BmܸQ_��  p5l��ņ�7�_xV   @& ��+����k��LZ�7�iS�}��W����Y�z^^����S����|��i�&����dԷ���ի���+�j=���.�p��y���  ��roiiс4k�,���.�~뭷����0Y�}�q����; �2[�38}�p��E�瞁~y'����XK��������cn�А���=��  ��HT�׻k�"]�]�   H�*��	�lJ[�{C��F�-О����=�[*j���z��500���nkk����5a��bǎڼysܸ7������M�  ��r?s��O�>]�=��|>�n��fr0�L�2%a�������      �U��{׋�	   ��qU\�{a��O�m����5��Fy='G�[X���Auuu	ߴ%CII�n��v=�쳮q�F��������ke#����'�o҇�F���  �'�C�v�o,���3�(
i�ҥ���+�ܾ`������֤O�     ��sQZ,2���   �)������=�����#z��F(j���F���߯��F�Ԥn9W�oذ�5F���Goo�{c�nݺ����,���o}K���q�-�U�� ��!w�[@t�ƍ.�>o�<7fQ#���7��q��v�����'     ��({п�E�Z   d
�j�_��	h9�ti�hk�V�����}�}
��*++K���u�B��r��B�v�zժU*,,p�~���i���q�6�d꧿kS�  �[��܏;&���&�>��#��ٳg����,!w c��>1w�ܸq[��&�     \/O�k�]/>'    �p�5	V�����5�_�WZ�5��ZՑ���Μ9�Z���S����R����Ϫ����o���3gjŊn�믿���J���ǣ��1��X)   ��!�#G��V���j��'?ѽ�ޫŋ���]̱6w +.n��1�v     p��ܣQu=��   �LB����Q��F�g��m��hLO�O�G���>wCC����\�'U���t�]w���wmk�؅jY�;p�������|'a��7�H�K�-  �ez����î����R�=���|�r7f��ϟ��S�ƍ�*t���     �q��a��j�t�   �LB��̟W���BEz;Ҷ�֞A��m����Q���H$��Ǐ���58���Ŀ���/��ӧO�pa�իW�4d����ק�~��	��3n֤��   �䐻��8��+**�J7�^`ժU���:�7-Y�D555q�Y��jV�     �;q���/ �
��F ��	�����G��%XZ����i�l�i{h�n��;���'Nhʔ)	g,'�����mݺ�5H���iٲe*))��;��o}K���q���4�2�"  �����m�t)7ύ�qlaa�Y���������DUUU�M�6���˭�d!w��c�  �l�c�l����*p��    @�$�Ct=�� `��>��"=�+M�}r&-T�b�����x�9��i��)���|&���Z�F���g���--Ѭ�d��7�t�������?�B{~�a�ڵ+n��h�>�&�   \�������!�@ �1!wkr��v;�߲e����;���9	�H�@�|�r�����G�     $S�����8vD   @�!���(��PO�b��G�ј�l��G'*��1����N566j�ĉ)پ�h�~�jkk��.V�۷On��͛]i"�?��ʟ�F   W+�C��ȑ#�g���^z���}��.�n�S�ǘ�
 ����j�*�����g+������gﾃ�>�;�:�$L��  )fR�-�
TI��[Z[��[w��;��u�ݳ���]��kѱ���>K�-�vO�i-�,���@��H1 $ q&ar�����`� ����TO��t�߯���      �����(   �p�����M:9=��?7����w����R��y�[�zww����\.�2===�{577���{������z�w��o���:~�K�z�w  p��=�>22��w�ܩ7�|�MH���>w5�n��<!w ���U�=��{�Y�ޗ �     �[ɀ�s?   P����۔��+[�ԟ;��������r���>?77�v�:;;��g%	���������C��x�]�xQ�ϟp��}�k_���H�Z���iǗ�L   w��C�n;j׮]:r��7}�_t���&�R�Y p�z{{��C]wP�^Oggg��     �z�x<�]��S��	   Ո�;�Z�cH��e�s�M���f3zٷK�S>����33����4�nm�������-�k;�CCC.$t��	���Z����?����d2y����՞�w�B  ��r�m*��޽۵���_��~�7~í�d�Nkv�f7w@u��4���+yP�p;     �(%��_~^   @�"�����l�Wr�¦��7��j��}ޓR�VF�[X���k����/�sh�l�X�LKK�y��:u�j���K�.�O��O�Ů��=��~�i��[  ��=�>99�B�{��������o������>��~�mo�� p'|>�[��^SV����     6J��B��g   T+�X�m��D�MD6�g�0ը��j0zL�_r�����������ִf׳ ̝��ݿ���9s�6w�455�?��?����u�󅛴���A��[�   p;�=�n�X�2΁�D��o~S��k��B�N��@�+�]�pX�>���Ծ��a�����     փ���:����R��   Պ�;�M�c����)��n��������a}~p�zc'K^gnn΅uzzzJ~�B0v����a�~����������Pd��?��?����u��������?(  ��P��Aǰ<��j
���#G���{�u����ӟ��{�1�RS0t!�J�w��^���-侚Mh/��      �Q�}�բ��xO   U��;֍'R�}P��s���Sٜ�?֢/�Q{�T�����_�g7��躺:���o��e-����joo�ٳg]�$����6�`|||K~��K�����%��P�~�o����  ��,���ٳzJ�r��b:|��[Y���YO?����ԧ>���!w������>���}����ۯ�s      l����f��	   �fܱ�����Ɨ���m��N����h���=���h����g�XȽxZj��z�P�C=䚻GFF\�����kpp�Mf�7 ���������B���z�p���]�<�Y  l��\u��-�~��Q�۷�M8}��\�����B����f�Ye2�J�>��m������,     ��fǶWܳK����   �jF��.�>�\"�\f�C��TV7ݯ_��i�l��XX�����������\��.�Lc�Ƴ������~/ڵk�%lV���S�����R<��s�Oÿ�M�<�9  l�j�������544��۷��ɓ��׾�/~�n��Z�m{���yZ���_�<�ZZZJ~�&�$�I     l�R���W_�7?   T3�Xw�v�Pb����H"���[_蓚�J�����������.���,D�s�N�$~��E�"N�}�َ���,�d��Y��&9��������;��/��/J6�{|�η���_  �V�����	���7<<��,����~V<���n�n[-O��i�����ׄ�l��^?lB     �f)U�y�Y   Վ�;6�/ܤ@K���[��b)��h�~�߫��ӥ����Ç���sm���[������LMMt_������n�R�������ۧ�G�n�����/����R���C���W�>��  ��j!�n+(�j:��g����kttT��˿�!m��B��lV j�Mt���G/�^fgg�g     ��޳X����E}�e   Վ�;6L��_�dL��Җ��H"��\h�?أ�詒�I$:r�k�nnn�V���={�c�MLLhlll�ū�5�����n���յ��?~]�������{�������;m��I  ��Z���ϻ|l����Qo��������/|�����.�n��y�܁�P__��~X---%?�L&�k�	     `�����k�H�0  �@�*ԹS����K'���'�Y���}����OI����lyqk�Voo����������߯��Iv��Iܜ��������Iw�n���e���z� �׿�u7y�S��~�i5�|D   �B��I���l$/^���������E7Y���n�	�5��^x��:W��'F"     l{�r���
   �ܱ�<>�����-�$�9���6}nǇ4=�|����\9}��;p�{��3�7�5�[���������lG�����׫y��{�qm�x�SSS��?�3�����|�}H{��Ӫ��/  �rT!w۶>u������v��o~S��ԧ��c���ؿ9�Ͳ�P�����裏������~x�64     ��V�rɄ���    �pǆ��خ���-�R���w6�O=�e�v��%�g��XL���S(�V���Xpzzzڅ�jUcc�:;;][����8p@�������o|�!��iϿ���m  (g�r76���m;ж��~�i�8qB����ݶ�M>�ɕr��3P��9m��zV�=�mu/&�    ��T��=���ʳ
<   jwl
c�r����3[�;�ry={.����N*�+y=�X��5z���������>7�ɤ�ۨ���-X����F]]݆�����������:>|���w���Z�������  ��J�ݶ�m��Mr�ɥ###��?�s���O�g�גݤSktP�l��&��H4u�^�Lh     [�T�}���   �
��4��!��	e[�~s<�����l�y�&J^�ێ=���Am߾������5K�aa������7����Ԥ��6j�Û������l�׿�u�9s��
�����?�����>  �$r��3g�U+���.�Ɛ{*�һﾫ;v��l[��;���}�Q=��.köU-�'�
T�bk{q߾��_����r     �r�:���d{�y   ���;6Oa,ԵK��.辕Nͤ�_3��|W���ox��/jaa���ot{����{OO�������;�Q	�wXK{KK�n/5}3�ڵ�5yZ��f���[���k�+�j����kj{�  @�
�3�2s��C����v�8�w�^�������]�����n"�m���T�խ�������������yo+s     ��R��Ｉ��   �ZA�����+ܽ[����f��w����7����P���ǔϔnj���[o����a����\����f7�t�y�BG��a�-��UlG���^nX���͖��
v[�߿�ح��D"������+��r���G��oU7�!  T�Z	���j���w�Vgg�fff܊=����_��_tۊ���m+�is����v����/�'?�����'�>?�c     PNJܗ>+   ��pǦ�B.䞘8�|~k��Ɍ�{Ƨ'�Ї�O)[(y=kr;}��[�|Ϟ=�ͱ��A�b�|�d2��Ҷa狧~���:k��a���8���Z�W/�V��w߷o��=zM��رc����n�����v�/.o�Q   բ�B�]���ﻰ�Mt5/���k|�'�䟸I��]kۺ���I� ����}||ܵ��>���]f�]      �f�1�|6��?   PK�cKxC
v�Pr��V�*���ze4�����+����^�B�o��o߮����	k�T��H1�c��^na%���f�۰���vj�-�S��ɍ������ܹs�����w��C��0���4����O�k  T�Z
����Ir��{ܿqddD��?�g}���c�=vͶ�zLpw�h�IE��|���~\��i�U'O�t�x      �T{{������
   �%ܱe��ʷ(57�rp�RT�ܡ_hPo�}�҉�׳��l���qm��+�tlTBK�f�믿�?��?t���?����[���   �Y���m��w�y�m)�J�g�ё#G\�{OO���m`�
�I� 6�=��}����Q��?��Ԕ;o�����kll��^�     @�(U(=��   �ZC�[*��-�J-L�,�R��S>=���>�|N���^wyyYo�������cǎkZ�P���̙3.��K_��Q���7��?�7X/  �ZPk!w��\�p�j��mZ��7��}����>���M�6Q���W��`�X�ݞE�dRt���E��n��XL      ���\NK���   �ZC�[.�ڧ|��¤�A./�1��h�>�բ�œ��2%�k�-�2;;��۷_moDe�0�ŋ]����Y��~������.,Q�ܩ���Դ�  Pk�!��4�\�܍���|�M������_}�U���{���>�&��b�����4E���sm�>��S�����=WMqr����\     ��p{A��	e.�Ga    ����,[�]�{ziZ�br>�o.7�#C?��g���q��WN�>���	�ܹS���B�)NX� D*���s`����M��Ylm� _�I   ��B�_����M���Ԕ��٣��&��������z�!=�䓮��B��`�]���k�ua�-��<��D���O��&+/����     T�Rez�C/   �E�Q6��C�[�#2�r�����ٸ�oݭ���y�r����Fu��Q577����]P���ܹs7]�����FR:���m�~R   �͐��m�#G�����5�[c�[o���'Oꓟ����~w=�Z����-���WG(�	$����^z饫���f�v6=��     PAJ5�/?��   �ZD�e%Ա]�甉Ϋ���G�W�=���>�>��칛^qqQ�V{{�������(����9�ؾ��|��y|~�L�k��O-�  �j5�n����q��{�n����������믿�O��t׵P������r��=,ܾ�����3�hz����lⲭ��zE.     �rW��=u�R��
   �E�Q^
;m�Ν�SoY5��\.��]��lS���>���I���n�5vp݆{�o��/(���V�v3��^M�syR#���/�/    \V�!w����請�[���.�k���������Fw���Tv��mA���R�v�����H�N��zY2�ԙ3g��7     @%*��}�   �ZE��ǅ�w����2@�f���Qi{�~}��G-˧�K�o�5��Kss����&l>Y���ؘkּ���N�:�^��Mp��}�i%/�Q���x  �e�r7�.]rm�6��������.���c�������ՠ�ܳ�,Aw`;�k����eb?t�^{�5��1�ܱUlU��e      ��T�}��
   �U�Q���.�Z�P9:?�_��`���h��<3'��fn�5���n��a�������6:�?:X�httԅ"n�j�;�6�d�G���$�be�Q��F��   ���{*�r�v�Tim�J��z��Wu��1=��:p������a!]kt�����R�v{~���z���Ů^n�rYk���      *��D�ZfrLɓ�   �U$kQ��}�!;5?�rd��o]�轩&=��cz�nB����ntO$�ŋ�������Z^^���km_K���ԱH�ތ��\��Û��0�5��H#?  �J�r7�=z��:::�s�N7��&�~���u�������B���N��ʞ>�2{�Jhta�"{n�={֭�      PJ��G�(   ��pG�����|J�^T��'3z�ļ~n�c��#uc�N���~��Wl9u���.�n�w;��;c���'&&�F��5�@H'cMz}y�f�&�h�R3��ֹ  �C�_��T�q����B�fffFsssn[ǎn[�V�������At��AwԚR���&����?v+q�s�&����=G      �E�����Q   @-#�����%�?��Ԉ���=�K�u�LZo�w���u��2S��Ϧo���HD�O�vMt---���T{{;a�5�p�5�Y��Dk;x��z/�MoD�4������19uV�}�x��   V���WfG���v�܍m�Z(׶U-�����.���-����O|B}}}��Aw[��0/�͍��6��������^f�[��J�o�o     PI�����dgg�8zD   @-#����oQ�w��,0����K�G'Rz��E���j���O*����k��5<ڰp{[[���)a�X�ǖ����u�ί�7�M��[��|�f�)�nw����	���)ԽK   �M�H�R:y��o߾�m�k���׿��{��F�b �B�6�6��j��t�Okc�A[����K�Pd����)��D"!��-��K    �����E^y��   P����xC����B�*.w�xJ/�L��@H���k�Q��e"�k�zm[+�۱mnnvawkx���S�I&�.�o�������x����;�V�;ۮ�h�pYj�~�LlA��I�{  �k�ܿ*B��Vo:v����m|c��S�Ni߾}��_�%����0��^v;�>��L���=~���9sF/���[�`%[��V7�F�Bm)�$;     լԾp��	   �u�Qq<���}���:�l|Y� ����ssz���=}�����SJ]:�|vmK�[���m�P(��6,�n竍-?o��⸓�>�?���6I��h@��������q7	�n   �U���g����Z��w?~��;v�p��v;���{z����e����g�w};�e!aŠ{�&'�){��W����n��dωs�ι	ͨM�    ����W�g��u@��շ��
 6�7jwT$�קp��ƕ^�T����zot�0���6=�?��f\�����m}/k3�t����ijjr����%��ʂ9�X�l,//+���7�x�k��{��:��҅�b0~c�.�ߐ�:����.X  �kY����=��4�<!������;卑�U۷ow��v[������ק'�xB���z�����t��Ս��cm���\���=Fm�W_}USSS�|����^�Ѝ�UI�c     p�JM����� �R�}H  ��\���`k����R3��WV�c!����I���hO���ϫ]�Ee��(�<s�������n��թ��A������X4�LԱ&v�ܼ�۸�P���E�S�t*?�S糊'���[��F>�q!�p�=�1
  �k����2sFO凕k���!�ˊ+6������m�k���w��Voz�G�(��d��6�v+����fm�z����'?q����~��.Gm�ײp�v�     jO����~,    �Q�����\�8�N��X�����B�v�>�}]	��+�0�L������̵�yÄ�aw����k�Ze2����8�J��N�]������t�BK��4�j��x�NO���������MF����`��   p=kr��&wB�כ��s�n����������s��СCz��]������iu�f�Q[����o����z���4;;��m�.��Ku)&�   �f�v�� ;�R��+����������)�ڤiv<�x���nj}� �������=�*�ӗ   ��;��7X�p�>%�G��Wn�[2�ձ�:V����o����v�d��."otJ�ً�gӺ[���Z�mo��l�,6En��/s��S:����	��#1�M
#�r�^��7��&`   �z��o�n��Ǐ�U���������m[���^s��������+W��[�����fm��8;s�~�ӟ�ܹs�<��qh��-�n+x��{y&�  ��f�Ͷ�M�D"n���wö�l_���U���n�~�}_���}n?�n ��xJ�{�U)}�y    �pG����
��QzaJp�S�snF��*u�iO�^�ͫ/WfqR��i�Z#�V�x}�o�R2Ԧ�hHӭ:s!�H��h-�@{)��n�0   ��C�_�+�@��F,hp��I��{oo�[x��w�u���M=��x�T0�Vw����]�����+u�Ղ7��kk���v2k�������8�ܔ���o��   [�B�R1Ծ���v���R�MH5��n���j�����]��?�w���` ��J��9��    \F�U'��+_�6��K������ryM�-��r�|}�^���k�#�^߼zq�3�Df�K%T�\�yS�b�F���4�kׅ��fcW��]P���sJN�Q�o��  �zr���Y=����V,<22�.��="���Ƃ
�=����y�رõ��߿�j���n�w��X+�;��s�&]X����߿.���]����c����/_��i   ���-,,�}9���l`?u��`P۷ow����������:���.�ξ9 ���%�TR�C/   �e�Q�,$m����Ee"��6�DZ'������/���=lP��:�������)]P6�d)y�kf�o���Y�@��!Mf�t)�䅘"�v�9U2�d��Q�{�   PZ���)r_BXpxbbB������QKK�;(f����m�e>��MMMW���;n�f�vc�o����9�/+���>o���M����k����  �["�p�@-�^.��6��v�������۰U����@>�W`}�z�%�����c �b�q���taNsY�0�9��O��y<����}��++]�h����we\�X���1 T�Z�.Թõ��f/\�G�ʤ�9]�^r��W���7���uvբ���Q���SB�dL�T�5��Q�q��<���h���W8��ZJ���k!_��\�����+O]y#w�[J6C&�(�[]    �C�_հ����n���7��kڳQlu����/����p½�ޫ}��������(v���];lbD�qp�P�ُ?��G�jll��'�I]�t�� ��^����X�  �[�ȶ��)�^��G���:|��[l�޽n���5;::�D���Y�� p�J�y�Y P��9W���$���.l��̺g�nŎoX>��FH^;�i��e��iՊ) *wT=c�|�F%g�)_V���r�Z���Z�_�m�-j��>�W}�_aoN�\\u���y��=���7/O>#�?�p��>��F�md=~%s>%�>%����^%�u��=�$3�̥�i-G��w�
_��+�v�&\��&\   �4��B����7]�n"�6*>��.\����V�����v]��~��F���O���W��ʀ�}���;���@��o�Zh��ɓ.�~������p��OZȅ�'�=�����i�  ����FGG����J����o�رcnU���a�ړ��m��B����r����|&��� e��ʥ�n�gR*'�?b!{��+r��] >X'o�������QlVV�g�2�Y�f/Vu��Z�2Y�,��X{��7)3+.+�*�^+�Vx}-l�*=?N�  �\�}nDOy������C�6,0jAwkڳ����/^��Ƴ�>�]�v������ߍ��g��v�ʶ��vc��S�N]�g���;�'m�R��f6*��V����%  ��a�N6Զ�+yҰ��ӟ�����M���Į�.����c4 `�J�7�Me�+k2 �JX�ؓQ�R1e�y�W�� �O�
��k�q���}�FWV�7���	@�!����olw��ܘ����$��N��  �[������]��r�c>�Fw�755���ӵ�Y��Xx��mX@a��ݺ�{\轱���u�vw�� �G�Yhw%7Y�saa����/�B�|���������	!c}�J��{ ��I�   ����m?̶�������?Ծ}����}t۷r�ީ�)e2 n�T�=��� `S�1�'"�%��i���e��n��{�r�݂�@H �w�[f$ԹC��V�f/���)�.�P�B�B�  �ڹ&w��w*�tyB�w�n+��l�={�݆Ű�ݦ�¥'N�p�����g�w�x[��^���un'�n���Ą��-�nA�R,�b!�<�9lE�kI��oR ��g�̣��7�Ʈ����7~�#q������M��� �`��6�lV��  %�N*_*�Ś��E.wC�v罁�+���5FS��W 6ǎP�|��
�(�0���뱮l9�`K���:  �;�B�s#z�3�M���n3k׳q������l����׹t�����-�w�^��g��J�@���ʰ��b}���j�Z�ZڭA��-��DJ^�B�sss��ݾ�������>�  @%��lBq-�m�G?����~�w�}�2��hm�?a����R��$�;���  X7���l2�llэ\:!ܞ\:Y�J/M����n�x�o�7��A�5���)�6�@S�R�c�D��-c�{\Y�   w�B�_�&wϰ���ד�v���n�>}Z���jkks#�`��t:���7�y���s�Nz� �5��V`�T�C��w��r�@�㛵�Y�����.`c����o$�Hhvv��S�Luuu.�M����   *�mo�;wέ�U+l�����n��~�箮Vܟwh �*��N��� �ٱ�d�e�l�ia}��+�K�ܨ��Z�kl#�l0җ@�'R�kX�����Ef��ؒ4��Ay�u  ��qM�3g���N�.��r__vZӞS__��6l���auk���k����?88xutvv�<XW��ju�8j�����0�Z��533���1��n�v�F��]�����k��b1����:cv.L��] @��Տl��Zekm���������[�g���n�Ě� ����|^K�?-  �T6���򬲱�s�3�v+Y�0�0!�e�,��ohs�C 닀;��-%R�@��i���Y�%pk��l�w��   `c���܈��+�H��F�гKہ7�ދ��"k+������ykw/�����\��P�j+�G�Y`_=n�5���bcttԝ�e7�ǯ�O6hR�V�����f��Y  T���I�=^�l���O?�O~�jj������o�� ����_�3'��o	 ��X�:�U62�\�I�[)��+ec~\�P�������	��#����(��K������^�d�J���
������7   �Xr�����!�B���Ջ��gΜqau���ncu����O�v�Ȯc��}}}���PWW����7~[�V���]�t�e���N��}��:]}ٝ��uqq�5B����Vv��f��E֒�2ОL&�kn�����VC�5  �������۶9.�D"z�g\��&G��rsY9
 J�O=�  X�|N��2K��&�B��%cJ&/�37*_C��zÍp��7��*��#��/)�8�|���(<4|Zz
"��  6��Ϝ�Sy�ܷ���ۘ��p�-�Z�777���W��л5��(��|�������joow�y�C�G��X�|~~��$�xjjʍ�4��c��"���a��#(W�zmw�M����i  T���~ߏ�c}�ӟv�����ݾ �) j]���g�  7��ڗ�]c;����v����o�p婴����;p�_��~�ut�q���o�v3�l   �F�������7ms�r�:�n�b����<��C��u_��f]#��cǎ]�9�[ �x�a-�vj�۟+A4ucyyمϭQ�B��P��<����c���vj�%P�,�d�	EO̎���v  Pa����߄�<��s��g>sub��#����.�f�*hH�?�Թ3 ��l|I��K��+��+5{Q�1tl�'��!���A�.73.�<�|��mz�|��Mp�`{e�C  T�enDOy��k�ɽ��r9�QdK�[��8ݰ�k)��g�ҥK%?o�u]]�+���ˊ��.����g�A�R��R�E�ؤ�N���e���6���f� �=��;����������T5��b[�iA����  �,69wrrR�9�oy��g]�{q���Æ��t��9�_ ��T{{�՗ �5�ye�s.�n�hT+�M/M��oV��G�p� �w�6y|Z�h齼Q�0閃A���݄C�v  �2��g����r���˙��>�Qd!skj�0���[��۸UC�"l��~wʂ��Yɂ���)��-�n�>�@�}���U`u�=Wx����Q  T[����ؾ�����O~0����������֔
�G��G �����L�v�آ�p����շ@i܁;�������ϙ؂2�,L2*T6�؆�m@xC  @ys!�ٳ�j~��M��e��+��7�P����5���~Ű�k�[���@�ݰ��;mY��7�R����0{��F6�de���Ч�Ϋ#��  T� {��y��LMM����z�ᇯ^f�s��� �
O�"�̥q%N ��Y�}yƕ�l�=�D�o����Z�Z܁�eA���TL��Y���r���X3���]��Ny�A  �rX��+s#��.e./�GȽ�Y��-ko�;0h��5 ڰ���x�xj�Z7���s_k�W6ތߋ����H���t�(�W٭���j������xMKݮ�q�|:"  �Ja��gϞݰI���������V���l_�V�ZXX Ԃ���^ ������+����j].Wr�2�Z���& �p֑7X�`{a��+�Sfy�V�2�B.��SG��MV   @e����͜�Ws4�ׂ����z��Kp�{���n��9{I�26-  �Jr���N��ڼ��+��_�7���Bﶢ� �v��#/<# @��ȬR��4��:�1�N��ς�m���:��F�x]hچͲ��{&:��I���]������  Phrǝ��x �`�%{�]�qaN��<!  �J�����i&��-������D��ԧ�^f����422¾:��f�����ܬ�G� ��Xn,=?�\�I��9t�8)}�m��jw`�Y�:�>�`�N6Q���r9��3��������v�   �:�ܟ��T�&w �v����΍���g����P�rK���?�\0�/wyԛ�)�-�U$}��i��Ϯ������j��g�J��k�����By�	��ގ�q��%�={V���W/�Bjoo��̌ �Zل��"�t� �ڐKŔ���l""�vdb��Ɨ\�-��/���/j�z`�x<n�������{l����B�C���   ��B�_��S�a�//�G� ֟������:h?4=�/E��r�"�Z���Z�s�+���֌��gN��k����-�{�brrR�dRX?o������]���n-� P�VO7�� ��Y,�0���4ǥp�챓^�q��@K�M�.��
��V��{�67��!�li���2����1����p�۶��v  ��B�g�T�&w Xof�`��R��l6�'.��/��  Pi,�n��X_�DBG���?~�2ۖ���-@U�c׫�٥E��|M �*���JϏ+��
X6a�V�,�(�>��q@- �l�+�l�־������7�Z��M�^�0���   �b��W�SyB� pW,|]㦽��P<�ߚ>��\Z   ���ֹ����ɓڳg�Z[[�^����F$ T�R���)���? T�\*���ye�Q�c��7�+�6 ���/��p��x|�GȆɥ�%"�F.Y��^���&4�W��n/   �F,����=%��`�,���������u�>�km���/Ŧx�  T�X,���Ea�=zT��G�������;��Sjųȋ? �
�sJ/L*�8�q'l�Ld����ohP�8��9t��7u����KF/�Sq7�jd�u_�A�pa��-|LC;   n׍�ܭ1�V> ��x���7cl����qu�h�  �mbbB�X�ϟ���߯��櫗��թ���M0 �jPj�:�*��A �OjnT�ia�,��J�+.�h]:�W>�q����`rꬲ�.�NI,�w�¸�w}�E�lF�T�j�=��+�N*�˪�r).����ʩ7P�2*   X7r��s����~������  ������҄vdR  �t�DB��;~���x�k.��. �A��㱟�DJWgq Ժ@k�k�Υ��Ev�m[}H�Am��)�WX1�+�FoZAOVu)����7oo�i�ȫLή�W,S���)��+�S�W_�̣�XJѤ�
��Dm�?���_is���M@5!=
T��궹����da��F�����5�g3.��3�<���,��?�7��q�Vv   l�`>{]�; ����1m����yu��  ���gddD��w�����^�������� �ҕ*Ո���  ��rO��]J��_���P@Mu��VG �vo\�����)�ӗ�Y�Q��Z+�=���l�XÕq����|�zy;�n�r�-��ZȆ4�k�T4��Ÿf���d���X�2���e�.�NՂ�;P�쏕��]�q�?[�
t�]	�[�{>uC�r|�]V���&Ċ�r���λ?��3m�el�&   ʈ5���; �Y6�U0U|YO$"ڗ%p  �O&������9r�������\���J�@UX���O%y� ��7X�`ǐ���T~�zZԻ-�.��C	��"�DN+[P>�A����׃�flU����qwY���W�p������n�l&�K�M&�����BT�\^�*�S.Q�s���JG��uְnM�

   �Ő��f� v�ݟ�FN�|N͙��Sq��&5\��  �������9��ӧO���-���n�-  ��T{{��ו�E �n��v�`�^�V�	���hT]Z�9�����]���,\-I�� ����w�04sޅ�wƮ@H��.i�Sc�:��Ztq.����J���&�LJ�ɓ
4�(��k3�T*�O    j������    0;;+l�X,���iuww_��B����ZZZ T�R���� ���A�1e��?����AC�Yf�k[F�����^�OW�&y.�Tj�T���]^���%�@�&ҍ:�h���eM-�US�mwjaB���B]î��D�         Ԥd2�h���'��ܹs��MKKw ͳ�%5��(�� Ԉ�����s�MgK��i�j㢚ScJ/NJY)����6��������^�rR�����M궢S&�q狗��|.��¸���B���~Ev��L�M��fuqf��Tv��&Z�c1ԹS��m*w          5innN�###z�Ǯ	���׻��FY `#�jo�y[٥ j��e[�=9y���ZGcH;�3��Q�gY��r������k��B�������h_=��v��ga�t:�T*�MR��D"�x<�N��v�����Y
�+��j�Qfh@��m:>�ѹ�����D�D�(�����*	w          5���cA���uuu]���/�/ *R� _��� �_�I��>��ƶ��77�u�-���i�g.)/l_']Y���m�ۄT;�QWWwW�����ܰ�]���-�����\�a��;
��&�0!Ʈ��߷�[��Ov蝉�f��D�I�S	;w���	��         Ԝ\.��:SSS�܍W��D���٬"�?- @m
4�(��*ۜ�<,>�ͧ{���9�\d�B�RSS��m��NmX��\ٿ�� ���v�r�ߋD"n�byyٝZ��m����|��!�O��Ф�[����Rٜ*�=s��+ԽK�@X@�#�^ò�eEO�. �H���xak�+        ʉ��v){ܝ��	�w�}�\v�fF (g���&��1ef� �]֖�O�tr�~F8о��l�QKvF�lF��ڿ���RKK�Z[[��ܼ�����6[H�FQ"������ݩ�*�f���SgԪ3z�n�>q���%:��h\s�	U�\:�ĕ���4 �3�,�W.U�Kf � vl��{       U�Z��������f]KdQ(����	 l�RA��� �m�O��].P�ϯo�wgSX�.��e��R�rDg-������5�[�}��x5�����7�Mz�����ܜ�x���%i��߇����\�~6��ř����[X���olP��         �9�hT�Z�\ε'vtt\s���/--	 *�u�����Z  x�u.H��Y�������u���W.��XnI;;;]�}e�y-klltc�����L���M�]\\\�7���>�3��ޯK}�z}�Q''
�:�Z��f��>�|:�@k��rD�         @ͱ���,Ⱦ:� ��T{{��Ie�F ��7�)��*�4u�ߣ=��#�h�)�I*�Z����]K��[[[K���e6���׍T*���v_������Z5����ݿK?�kѻ��tO-L(�N(ԹÖPN�         �)�lV�tZ�z�#�T����"�^  +�\�=������CY=�;��R.�|��_c������*�w
7g�#}}}n��qMNN�ҥKkڇ�D�*�O�7���Ӆ�?��rιg���[��]�x}�w          5���򱸸x�e�T����  ��x�ޥ��q峷N�w6����y��)�II��_?���[===���ևݖ;w�Ԏ;\����n�u�آ�bo�Z������L��N��~+d��JN�*<Fw��#V���#         @MI&�By ���y<��.K_<���S `5�/�Pװ��+�����c�˅?*�[6���a����`;m����wvv�a��n�r7�y`����7�Ϛ:uq��^hz)�rd�$&N(ܻ�=V��F�         @MI�RBy��b�]���\8�Va �j%��_9(  n�nR��O���k.�z=ڕ���5ϫޛ��7�>���P[[�����}xxX���.�>66�L��32���մ���:�ۡF�'o���r�'��#�����Z�         Ԕl6+��X�}uH��;�JP��=��?
 ��	4�(��*[p�{���X�iu�c��m۶�`5���444��/]���/�r2uz��x/hx�N���ň�*/�C�'��+O $`�p         PSN��t:�P���D�Vd ('n_p�LM(��Q p+��j�=��=�toÒ򹛷y����0�5����
T}}}������䭃��Q��}<4���Տ&4�W9�eR�O�P]�=�ܱe�         �)4���R���D �����9tP  �E��!������/}A�\��W__��۷���C(o�m`A���nMLL����Xu#�dT�ɷ�?���g��z�|\�\����i%&O*l!wP�f#�         ����^^��}�խ� PnJ�NE^|F  �L6����7�9�w���*����߾��J0Ԏ;\X��&��F�.�����A�cz�?�����3��4>S��&���)�{����L�        PS��߬L�����@�+嗯�̟�ȟ����֐��u	�a��	�_���u&�P>{�C ����._���Z�ϟ�\�}"QM��ok�~7_������o �Y:��F��/)5s��e��3�<��|�3�[8zpp��j!�~�_�������ٳg577w���3)m�=����՛-�z�|�l��s���{��܉c��h        @My����o(��I�<�����V<���~Ŋ-
@���<�AB  T������x���u}�����=�#��D���	����{���-���ox����Ϫ�=��x�����;o���=���}�b�K�8d��h	�B��l�-����������0˝�t�t��2�f�ܶ����]��BYI�$�$N/q�/�"��u�&�8�'�dY�~��<NΑ%Ŗe����x�B�1y��+r�;$�;              @��[^��o�!OǁI/SRRb}\�l������TVV���R9rDG�U(�z93ͽb�}��,�0�@�u+��ny��3�^�qv��;              @�m��Z��5�:�ͦ6��nS^^���߯�k�Z�S�	��^�|>���`0h}<��px�)���o������TFF���l�X*0��E����R����g�r�芜~�?�^ϴ9��4ۂ���-ʮ\" ��              b �q��Ꮺ��Mz���r�y�Z�r��}###:|��5�}����r�\��㱂�c[ ����=''��f&����*??���\c���瞫��577O:�=��r�.U�U�_u�kpԫ�u��lWVi��x"p              �!O�5~�4vt珞���t�-�D�;;;UTTdM�N6&Z7�M�~,j7�{"� ��v[���tw����������|.���Qii��Q�C*i��k���b5�E?#@"��dwd)�h��x!p              ���폩��R�;�x^^�5����ϟ�z:t<؞M>��
���LhOF�`P����f���V�n6����r*&�_�v��9���6��ᨗ�i�Emͭ׶6��_*q|m�efˑ[$ �              �D8��_~^�?�+���,Y�D���UQQqʫ3����ۧu��)##����"��ק�������
3Y����ښ�����m��eee*))���'�ͦE�Y�����.&��uq�J����2�^�nB|oO�r�ϖ=knL���B�              p��~�Z�W}[���	����w�=�y��v�����Z�z����rYA{OO���Ɣ��^������|L�>o�<���'U�^XX���;O��'ф���PѢez��TcހfK8���Q95+es�##�xD              ����_�_�Y#���z<''Gw�}�֮]{F�o綶6-X�@�f���N+j��|J'fB��ښ���&r����&�'���Lka��޷��Z��#�C�=��U/�/zk58��l	|��6+�j�Y�! V�              ���Ӥ���>Fc����O���3�����$�6�t��
o���f$�����󕕕5�w�Z�`��P }J{��Uw�����9��l	��?ة���B�              0cmo�����7�5k��#��Lǂ	��?�|egg���	�&j���J�i��L�7ӏ9bMu���UQQѬ�'�����Ӿ}��v��^&c�M��z����j��'�o�����/G^��X p              8�Ѧ:��k�z��+�Э��*����4ӻM�v��Ӻ^�׫��v+n7��1=f�}__���	�&t�7o�l6۬ܟ��\+r7�^�>ڣ�J�����y(����mVn�J�2�l1p"w              �)�����^=#�Lx~�7h���q�m�˥Ç������5��������k��8s�����`Mu_�p�*++g�~8�Z�JMMM���~�1��/9�'�:4�l����6)�z�4K�:�              &1�گ���?R8��8����{�ǚ�O]]]***RUUU��cccjii�&�#���ք�f���E�TQQ���`&�/]�TYYY��9�1��+:����u�/����s�+��N�L�              D1�緓��999����bŊ�ܗ��F��章���>��oM���db{������﷾�K�,Qqqq��Â���f�{��w���5y(�W�sv��n9r
��K�����              �$��-j���Q����<����:'J(Ҿ}��n�:eddXQ{kk��ٙ֝�\.���٣��2k��Y�&h������:���[����y�t]�A�2|��C�޾V�֮��A��3�#              ��C/���R�;q���H��������/��kE�>�O�G�=Tmm�.\(����2�שּׁ,��f���܏=5r�gX�)n�/���6���_��VeW-p&�              ����Wt�ޥ��q���p���c�����`��6������^%%%1�~��-�ө����q�1���Z�`�u��"wۘS�-=���^C>%Z�=(�H�2
+�.w              �qޞ&���
�EF���#9���o��***��=#cfyn0TOO�u=&n�L^^�5=�ȑ#Q#w��O7���h`��G�J4_�9��ef8�               ��{�����uG+((�����Z����&�/_�\�������p�
������i}Nnn�-ZdE�&�?Y��Gח����Yr{J�p8$o��̯p:�             @Z��t�o���1�XVV���~�vL����޽{5�|-]�Tv�}Z�744���Q��v�rrr�Or�����ު<�G{�|��ɜ!�PFA���"p              �+Rӷ�X�C/Gr8��G?j���������ȈV�X����I/��x������g�s,rommU(�WzZtuM�~Ӗ���7�&Gn�l�eL�              ������;~��f���;�Ԛ5k�	3����_W}}�*++'3��{zz�E&N��'�GF�a-4���z�ӡD
V�=o��� p              i���/��ė����u�%��	�744hhhH˖-�N���*(333淗�����:���)�8�=�k}�Au-W�pb#��k@��$w�T�             @��tP�w�N���K/�T�7o+]]]V�~��g���4.q�1������Q{{{ı�ϭk���h`��%����rkW��#�
�;              H+A��~�=
�G3S����200��;wZa{GG�6mڤ�����fQQ�|>�5-�d��a]?�]?�T���^����Y<_�T�Ә9�C�y� ĕ�.             i�Cj�����qh޼y������A^�����z�嗭i�ǂv�ۭ����ڸq��Ϗo�]QQ�@  ��q�x��YU�'��+���v)��\6G�&�c��8���Y              ]t=�e��M�~!�{����0S�v����
#�����>��.��b-Y�$�����ʺ���шc��&�)_�7�7�4
���PV�"�!p              ia�y��>�@�c����p�B3q��Q�۷O���Q��cB���n�*�׫�+W����l6��֪���
�O��u�ի�T��G��QX!{6�I�;              Hy!祥�y���l�ƍ���K�)��e����V�>�pX;w���Ѻu��v������݄��9uM�Q=�Q V���۔S�B@4�               �~��t6D�_�`�n��6g"j۶m֤����3��7�|����=;;[555ք����:���H/�%n�z�;��{P��'#p              )���������333��}H�8}&L���QQQQL�ˈg�^XXhE�'	k}^�ڊW��P@��sv(��Q��              RV�կ�G�$�[o�U���NGgg����k�ⱈۏ1��Ylq�9�(^*++566fm'
yFtUI�~ક/R"�|c
�:��_*�D�               e��'��ؿf�]v�e��D�۷oWnn�����ݻe�۵z��\��f�u477+N8V0֡��s��@⦪���0S���p�;              HIC{�R�K?��_PP���ˊ}�S	�BV�TXX��۵k�����lٲ�\ff��ϟ�����c�v���LݮMq�{PFA��c�   ����,:2��������oĞ���l!y,g�?�       ��
yG��ȟD=v�m�%$T����ب��V���(+++!����>//O555q����"���hxxx�~�LW����C�y��?ة��2���8w    i�%+W��-��f���Ft�p��_�6��Կ�/� �4��Y^��r�)+���         ��?�Ky{�"��Y�F�ׯ0���~�ܹSeeeVܞh&r��u��W���4.�a����nk2���]:��B;{�>d��e�;& p   ���ۓ�Kfe�8"���'���<=R���       �Y4־O=��׈�999��?�c��z�z饗���������~����?�k����ǚ��Puu����&�ti�Qʩװ'�D�v��8w    i��=��O��=��       0��~��
#������q����o׮]Vqq�����~,r7Az������w��>6��y���R��{tɑ�<_{�w    i��}� r���}� r       `v8_����x:bMM�6m�$�d---:t���ʔ���d�t:�ꫯjÆq����*�\.�B��Z�۫7�+�9���w��B�    m��=&r��lz�P�����""w        +�������f����o���{��ofj�	���=�� ���\˖-��ugddh޼y��?�����v�d�Va�_plD!���ɷ� �E�    -��]��u��t�܉��."w        ��ɯ�����L�^�|� #��_�����31|ǎ*--�B�X3�;44$��3a�|�iyi���y��?ܣ�y���F�    ���}����}D�        �_�=���|1bff�n��ƛo����i�	�ڲe����Z�qK�,UUUjmm��?
����jZ�`(�s܃�N�Kke����;��B��#}�)>B~���G��q2G^��/4�d�ˑ[���Rk�����S  H��#]#w���A�       @|u���Q[�w���tj����v+n7���b�~��Ȉv�ܩ�/�8�ם������\�	����Z�_��#y��p8,�H��Jk��E�
���H��=���i����~��Ə�*���mٳ�QP���om�h��e�=�,�Ԭ�=+���   ��SO�E����       ������E�7���͛��eb��۷���Њ�SAcc�����hѢ�_wee�FGG�����?_ZЩC��H���H��Jj�Xy!=�)&����n�����Gc��tRpl8a��L�����H����ɮx+tϭ]e}�[�Vy�Γ�p  �q{�J�ȝ�=u�       {��zP!�+b���^���\!��Am۶�
�KJJ�j^y�+F���;;;[������ 8�yC�����pЯ�ؐy��}���s�yw�����/�u�E��씯�MIo�����چv?y|�=3Gyg�S����_�^�[v�2  �.��ԗ�;q{�"���k��       ���;;��̷"��Hw�ƍB�ٿ�:::R2l?���jǎqy�WTThhhh��q����],B�����1w`	rzY�{���5z��|n����3���jm�d�֨x�;U��J��;  �T���G�F����%��       �X�z��
��"���]�Rf&﹤���>�ڵK���)�s��k[�paL����D����׊�*�1��"�C�
�d����;��|�v�~JC{�����)8���h�&6[�d��o`oVW�m���Y��v��V_���ߣ�d#�  ' nO?����"w        f&86�����_TT�����Bz�x<ڶm�rrr��=��)����WVVlC����S�/��қC���!�
���YR-�w 	y�k`�O5��cr�������/�2k3�����������E?U�>��z���|�G�kdd��h���ke\�FGGgt����Y[��_WF~�JֽG�ݤ�s��=+���  @�"nO_����/"w        �\��uh�5�\���4`��W^y�j�
����Ƭ���ׯ����`�t�&r?QQЩ�r��4��x����)w I��Zߊڷ�T�ͯ���L�nVe�S�TWW�����*++������lk���˴��W���ޮ��N+~?]�Q������|��w���v��׾K6Oo  ��v��ȝ�D�        ����k�<��������ب��Vk�k�����СC�������cS�'�u~�Q5�-W��>�<.�s
����?��,3/����R�����|�z�?SZ�l��,YbE�uuuI��L�7��l'2�ݛ�����r�������������e��t�-�|�ǔw�: ��F܎c�j�N܎c��       8=}/�P~gG���/��؉�400��;wZ1�����$�W_}UW]uUL��������vO�_�=�꼐:������"pO;��,p�����R�K�OA��]��ľj�*�}��Z�t����5��U�k֬�6���5�8���k��ɿ$'p����Z[��Uq��T���� �D܎�͵ȝ�'#r       `���Ո}�C7nR������ۭ�qYY�0Qww���ڴ`���^��Z���C���P��N�f���7!��	4��c�~�5ڴ�??++K�W����+WZ�S��fSmm��]y�
�B�T�={�X[{{���g��Uk;���jަ{Ty�Ǖ=�, ������+�;q;&C�       �������7"��_�ޚ�Բk�.9�N	�{�׬��n����V����&�?;ߥ-n�\������ȑS(�w ��k����������>�L5?��s�n�:kZ{ff��/��%K��nP���Ӫ>|ؚ�>��{H]O|��>��w��6���ּS  `n"nǩ${�N܎S!r       `j��|'��+��BHf(�C��)���622b�t���1�N3����D===�F��֩ݪR�G��i�����C�O|I}�w+r�.��	�_|��;�<�t*�T^^n�5�Y����k�Ν����!��kk�_�^57��JλN  `� n�t��ݼ2�!�"w�vL�;        �݃x�g�,X�E�	s�	��o߮��b+n������ �X���������W��O��O;s�Q�����^H�@��{�����ۯ)����Nf�ԥ�^jMk����ϜR��x��utth˖-ڶm�FGG����ï�Зޭ������l�-�  ���t���I�����t�       ����+�sG�ߴi�0��AmݺUv����p��n�5�~Ŋ1�Ό������rM�_bw�:ˣ_|��p0�����4B���gV�́��?ԭ�_A��|{�a�y¿�K�q�FUU��4頦�F��z�n��&k��������>�G��~��_��D�u��;  ɇ�g*Y"w�v�)"w        &��ÿE�3CE/��Ba�ڻw����TXH�<S�k�l�2+L�������]
keV�:|KoA��{!pGR3��=�ʩ^.[�F !�:�u=�娫�����UW]e����/�7�u�袋����]�<�uʚ@ 0��6�ԡ��W�ߦ�w|Y�K7  $�v��lG���)"w        ��nݥ��{#��N�D�{�=���������=F<�����|��]gAA��5e�D��z�c�/����c�B���E�
y\�t7*
��}X9�g'�T�pX��Lm?��|�GNyq��}_�j���\�RH���Z}��7ܠ���FFF&����K�����l�-�{��=o�  ��!nG��V�N܎X!r       @��h��60�r�1����R�����o�>���[�b,��1߫���	��~�8t8P�x
���d��R�;�҉q���7pTY��F^T�?���WOyY�n�:]w�u��v̞��"��=���W_�^xAO?����'Y�e0lL���ZU�|R���oNo �, nG�%:r'nG��       Қiz��$b����-[&��PH����5e��$�Qt:3��ڴp�]�i�N܍e�V���f�{Fa���ܑt��y��_�L|��?�#{v�2
�5[ý:��>���~x�˚���.�����!ydgg[��7m�t<t��K�0��:�����Z������  ���ȝ��B�       HW��m���D�7��c5���~������T���B|��w,���<edd(Lؿ�$��|�7��
�����;��y���4E������Ȟ�;��)��4��G�W`�]�f�n��f��$����+��R7n�3�<���zJcccQ/�s���_nRɺwk�]�������  ���o�܉�oD�       �t4���Q�_t�EBr���֞={�i�&nGb���j``���ǂYHRXX(��9a�=�U��tX�Of��9��XВ�ܑ4���=�ǟ{^Ƅ�&�ϩY)�ݑ����>���ݧ὿;�e-Z��n�I+V���_s�5�������V�>���~����k���jn�kͿ��	{ �N�ۑ(�܉ۑ(D�       ��˹���+++U[[+$'�׫�[�*'''f�5NOcc�֯_��+((�܍�9N�o��ʞS �6w$���j�2n?~Y�W��feW-��
���Կ���9~��)/ZRRb��� �����)o���Lt��O�ݻwG�\���џ|F��=�%�~��  ��v$Z�#w�v$�;        ]�[w��l�ؿn�:!����^���5�����Y��22b����n�+���Ԓ��2�l�N݁�D��"pO�u!ߘ<ݍ�t��
��d�Rfq|V��ǯ���wkh��S^��phӦM����fH����u��=�����z9ס�����U�m����&  03��-��܉�1[��       �`p�o��?������dE�fp���1��~�Z[[�t�Ҙ\�l��###�g=���]Ŋ��ǥ8�� �;fU�����i�o�]��<9r�bz����L-LW���[�b�n��v͟�Sj`����<���~ZO<����df�Ƒ|R#���Y��2
+  Nq;f�L#w�v�6"w       @���k���Br��﷦����Zq;���Çc���Q:��=hw�<w��[�ۃ~�)oo�r�WȖ�=��cV��<r����`�������o����vk%R�9-˵�^��.�H����u�����s����i�GQ�9W  Lq;�řF���HD�       �T��hӎ���W���Jfp�����p8TVV&$���^�\.+L���&�//��A�U8T��=3GH]��	��u�z�����H��I��gK3��}i���5vt;�st�wX+̐^�͛�O}�Sڲe�{�1y�ވ��;u�Q���Bu�~~F�I  �q;���F���H6D�       �T4��)�9;٪U��ٵk�.9�N	�+���M+W����effZ�Y�p��찊2����S3И�=��#�Ɵ(}��
��bru!�[޾#ʞw�}�������*���2fj��߮6�ˬ���ˬ_�?��uږ���_}A�#{��*���  L���j��;q;��;      �t�v�����z$A�Á�!��ɞ)[F��9�rdX��;��7���gZ�+V���ѣ:p��5,��}nhii�Y�n���ih��2��P��U�x
z\�(�R�;�7pT�)b�3p�ˑSpZOXf�{��P���W��X�d���nk�7`TTT�ӟ��~������W0�:th��z�/�iٟ�L�K.  �����T�;q;��;      �T���z!�������-�:�̢yrTX�4��ȁ"���թ��PH���a���+*..��v�r�\*((������G��j�N�7pyG��F���
���?������=+W���S�׀�z�F�?7�e�v����zm޼��3p"�0��e˖顇R�e�c���_��>��/�]  �-��+ފ�m�a�sB�N܎���      @���s��7Ц�����6oO�l��*�QV�"k�&���j�W'cz{b�!�/����M��M�pؚ���3�=��
C�Sq�{�i�;HY�H��g�
~��<��295+esL��6�9�����80�eJJJt�=����^�T�.]�x@�����gϞ����WM߼C�����7��H  ��c�ّWb}<��c�!r      0��CA�7�v~+f��m���4�o-�,�TNU��%B���|��f0%c߾}���VQQ�0�utt�,p��̴6��?aqVHy6���lœi�3s�;¼�4/4M���	���m�^hF�]������N9E�D���G�S� �aV����z�������
�N�F��?�?���ꬻ�#[F�  HG�혫�E�W�����혃��      �E��n�����=RغM�e�V+���3i<��H��l6�5����٩�{������=E��
�@@�ɇ���5888qg8�r�Q����3J����wf%���L��؈����/4k&�w��5}�N�I-��ꫯ�7�`�F8��y�f���顇���h�e�^xD��#Z����#��� ����Z�v�Y&r���&nǜe"���˴��'       Hf!�[���
��g�>���
�)�f��*
��հ%b_ee�
�����ۭ��&nG��V�^[[��3����}\M�Km���ZP�wĝ9MP�VR��mvʞ�w<"����t䇟�&iGcV#�y睺�����ի���~V���7��'�������u��z:b  �.D܎9.h0�%f�9       �93=�ݺK���u�m{��Q�µ�1gV����8�����
����D�, H]�k�E����UPP�XM^H�s���2w�U`�W���ܶ��E95+���Wu�'���r��ź���x�b�PQQ������w��8�{����wo�ٟ����x�           �\8���y{��������؈
�n�n"�̂�C�-Z$�Vcc�Z[[URR"�63�}&�����vUU��v����&\���.�G
��9�	�qcN���I&&U��[����2uuu���?���R�dN��O|B?�я�eK�i������Lg�wʭ[-           �tKcmo��D��Lwڢ�%��+���z��,b���W������ʈ�����|>����N��L�n>o޼y>�Lq7�y��viD�'��B8�ζ�6R�;����ޞ&�	mv�@X+����U%��z��#.�|�r�������Cw�?�*++���<��S����i�TV            �ĤEVC��B~�\���`��r�'�hKd�n�٬����׫m۶Y�ryy��>L���߯���i�y�Yq�ɢ�F��K#��Oa���=E�#.|�-�/꼳s��O�gw?��ϝo�uÆ��S^x��Y�n�>��+3�'6���͛����G}4bч�G��Қ�w�:           ��pؚ�>��c¡�\M����R9r�7���ݺ+b�6iZ��ݻwkhh�
��������@��,kkk'�Laaa��e�AU|�^���8�#�ý
�5[V>w<n?�}�{����u��a]q���۬�|@�lڴIyyyz�G'���������[�J            ���}H��#�k��FoW�ٗɞ�%�O8���7#�O�bj��kjjRYY�����e���B!�s3Jǔ�5]\4�r��7��D���2�{��{���V����.��o�`���*�^{��ٰ~�zk��w��]keۉ#}jx�*����]�D            ���v�\�Y���^4�7�lƋ��M�7b�����c���ܹSEEEV�8��I�y�^���+''gZו��k���W�;�Q�U��R�;b���2�$���^��]��h���{�.��r�ݻ7�H��k����ӷ��m���	�����+��^PV�"           �3@�����z������	���>uUU�0=f�֭[e��U\\,���cm'F�>�Ϛ�_QQqZ�e�v����	������
���>d�{�"pG������f��:��{ϙ��)g�u�,X`�yѢEjii0[֬Y�{�W���w"&��So5��5Z���(�'           �T�>�W�@jL��<����r�����3�}zv�ޭ��kj;�����dB555g|]yyy�{�-�,��<�{�������;~g��v��ݺ*[�#�����g�˥��>�ŜQ�D�f�{(4���:��k�⯞�=+O    0�T��*8�<%��kD#���O+�_��6
/ؠ�w^���y������_˵�5%�M��_��mRFq���m����5v���-�9*y��k��u|�y�qo��Z�g��?���id�v%Zv��_���u
:�|���z�    �Y��pv���4vt�
�],Ğ��1����Jarmmmڷo�5���S1eyy��35Y9]f�{4y����A��S��lBj!p�̍?9x{��?��h��Vݼ`X�Y9Q��Efb�ɖ/_n�:y��Hk׮�]wݥ�}�{�??��2������-��O���    sI�ŗ���T��o��{���Y�r<ٳ���￢y��2a͇�W׏Q�?�eBC�h2����k���>a����~A���z\o�`�Z�?�\e������x<����/Tխw����,\�}wݢ���T��O��O>%[F���u��z�35=�)�|�&    �tg�����H���]�,a�x�y�Lp��ɱ&E#���u�V[q;03���,UWW���������i@�c��p( �#SH-�1�P�5�=�2ܽ���Uy�Q�WUUi�ҥQ���F+W�Ԯ]���^�6l��ؘ~��Gs����gUwۃ    �\��5Z������W+0<��9��G�����]
����ſӬ�ٴ����[�Z���������+D�QR��_�������/�l��6��Ur7�K���~��N�7?6�C���}     �-0خ�gT���}P��UL�1_���}����D�PH۷o�>���	�����_p�1],b�DS��W����3�{��	��;���(�J���B���[�'{6����u���iӦM�O<q��W_PV�"U��7�    r,R�P�>���]Z��[�?�e��W]?~DޣG4J7�Cŗ\6�e~��}�1+��$l6-��5��
*�T�^��'�~;Y��U�'���2��h-�ޱM      M���t7*U��
��*��R��`g�>����ۧ��N�������Alܸ�lx<��]�d܋3C�73����3�h��'�	�ogt��ڨ��J�����v�����t����:����͛g�H���0����zh۶�7z���ϔS�BE��    `�J��&n�{��+%�}�˘)�%��C�?~D����Ny���b��^�/='L�|�J߱Y�����MŻoґ/�����q���˯�}�7.NT��k	�    HcW��c#Je��f��L8�W`�?b?��[LԾw�^kb;q;�b����mذ�|"���d�{�=1ܑz�q��N��;��d�����O�gffj��V�n�l6�������݊��/u�	�Z�d�	��l1��;�ӊ�<8�y����i���TVY�     3�U1/~�]Y5��eϯ�l��}̪�/�Z�³���YY����:��/��v��k5�5ӻ     HM���Ju��>���3s���u[�POVTT�t�v��u�V+T60���A���뢋.�z���>�OYYY3�-3�l�`p��\{PqG����qf�_<�g�g�Л������L�n�����k���ak��	�+**���l+V��믿n=Y��<v?�����TOOτc����i��˖1�    ��|}�hm�;�w��^.l��ݶ-��u8����0�����o_W(�SxN6�Ǔ��     �*
�?إ���١��%�����?f


��L��c�k�6�q*.�K��ź��+OyY�E�n�.���=?3,Ź?��S�*����_�����3�z���N9��L�^WW7�i.Nt�ɸ��ˊ��͛g�[�r����c� f�Y]y���[����p�ոMm?��~�k    �9�3O	��PH�/>�d�Y^���nT��     �l1���%>4S�	�c#0�u:�jmm�����<�����v饗Z��t�{~6�yr������D����)0ܣ��{�)�C%��O�]]]m�����xoo�u�3�}���jjj0������ַ�����O]��.V���    ��y;������?���*�U�c���Ö'     ̆��_�"0�&��f���"0:u��6bsY�v�ܩ��2��cJ�1ԅ^xڏ��J��>?'[6WHa�]�b�w�z�q�����O9_�|N��D���vs:�3�p8�m`�Ef��ϗ�����֮]����JO?�tı���U���3�     �gB�?���N3���cj������W�x��4�m�      fC:�
�u*��B����u:�]۲e�rssU^^.`*&l_�t����x���{��*~��qZB�/�f��~]��4���Bk�z,�.\��{L������0[n��F��B����j��;��o_��1�S�    @2rܯ�]���v��r���>�i*�o{�_zN�_h-���q�ئ������    �Ya�h�F�NL[E�>s�Iw3�4��޽[CCC3���066f�<\q����|:z ��MLu�+V�PHH=�8-���	��߈�]�7�ėq�<9WWW��6�*�뮻NO>��8`����ͼ��{���}N�����6����?����F    0W���Z�k0��}o����03���R�ekj     @"�}nk�y:1�1sAoz�---:t�����bJ=Μ	�M�~�%�(;;{��+���������S�;�-0���`����(rz�y"����t��L�p�֭ӎ;����g��&şs�93Z�����"}���7��kU�:�{��Y�.  H>W]q�֜]�������!��7;�Ե��ź����ˍ�wͶ�^�~��u�
 R�ͦ�wܭ��}V      ��d
w*��9&[(`�������Q+,,��v`*N�S�{�*++cv�'7i31i��S<��߀䑢�bn�	��lO�M�wo��sJ�������ɘN��^RRb�|z��r^xa��z�dk֬�N%���N����h�?�.{6+7 H6v[H]=���.Qf������!9��Bjs8�r��^Q:��A��з�gLG���n ��ʛoW���I�!�     ��	|J7��W���
��w35{�ְ֭U3����k_p�1��P(vg٘��t���4;SH�H�����Uȟ�_�S�,���)�Iii��b-^�^�5���R8ٱ/����dlB��=���M7�d-�ho�����uH�?�k-���  �����3�"w���vY�`�lA��9���:����[Z�ĩ
�{N�*oy�:��      &�W�11s�P0��TJ�k�.kwQQ����A��1�i�&����l,����������R$�@\���]	������(���n�����'���֔����'Y���Y��a�瘕Q��sz�}�C���Gk牺���n�#,�X   ��R�~<nGzI�ȝ�@����#�����p ��X     �c�H9��cf��o����r�vL�D�###��⋏���N@n�s�潿�4��
$B`�O����t��%�q�y�����ۓ����{�9���O�srrr�m�޽r��Z�v�***�Â�y�f=���Cj}��Z��Wesd
  $�T�܉��\
D���  eͯV�U�R���      ��&�����].��o�nP5q;03�w��՚?�R�����웣i�Lo�N���c����^Aıy��Y��ż���>�kVV��577[��Y�|�.\( ֮��:�޽�Z�y"��=�~�_4���)  ���r�N���܉��U�^w     �06�Ci�>���c�R�n�p�����|*))0����LW^yeBo7��m�,L	C�'�lB��)�P��M��zI�5����i6JKK/o�񆚚�f|=����Ϟ�566Z�����JFF�>�����x�������({�b ��4#�C�C�'n�1s0r'n�B^���ae��;�eϻPkϗk�k     �7�c��!C��o���=�}߾}���Z���\�1 �����.�il>]�E��{���%N�M��ٻ�6�;�_mɖ�x��N��'�@	e��BH�e�G����u���޵w׻�w�u��c��$�e�4@BBvBv��$������M��m�~_Y����N޼����y���T�-q��m��X^��︼h���j�Bz��)�۷O�۔�5''���ذa


0w��1y��3i�$,_���{�=8������ADDD�+�B��SL��R#��p;�E$D��C��|5��K���}� """""""Қ�l���V����Hf���سg�lײ�+�>����ֆ%K�(Yñ�f�Q�M�����"+���$�S�X
�[�w%���َ�f�KQQ�Vm:~���غu��+�d{�XI��tbѢE0�t����[n��ݻ�NNO-۟E�o"{�5 ""��
!w��i0$Ƚ�Յ����ԯ}�����'����5��s """""""Ғ��ޘl��7k�h͈y���!y�^%�f��l�!Inq�ԩJ�}��Yxx����b���䜯��I�(%�@[��,E�1oJ�p���K@\��ǦM���/��j˖-ʛ��ŋ��Hȵ�j�*<������ﾆ�������7n""�d��!w��)�rg����(�܄Ɨ�CѪ;�<W��.��~T�� Jeƒ<�N�f+(���q�v��X3IHY��������Ȋy\2_�D
��ڵn�YYY Lgg�R$w�ʕHf�z�աP(�q�ƻyX�=%Y���E�ۉ�ϓ�;�qݿ�߹+))Qu�P�t,�{�=ttt �22ί.�����,X����%�\���~UUU��{N�A�;����ADDD�-C���p$cȝ�vJ�3f��}�+&��S�B�-��5�_|�'q�?F��Q�r,_\?�[�I��d���������� �=��v����争%�*��8q'O�T
�fff�h �@@�����b� ����T�=bָ0�i)I"�l��ׄ��(��?ܞ���á�}:tgΜ�X��lJ;p� <�Ν���B�K�Y�?���E=���7��t�.��"""J5�rg��F"�B��S*w�
��&�Ws6����p)�SA��s�0��߂�K.�\sv
o^�����Te**B�);DDDDDD�����O�]��<��p���Xknn���ۑ����ۉ"����v�nnn.����eׅ�Qۀ�����H]�S?�P !OkB���E]ݿ�
H^4

4�O�`�ٳ�BV@���(�����1c���A�ɓ'cѢEرcG���ZԿ��(��7@DDD�/B��n�QH��;��,��O�w�ш�Uw�����T�殸��:YJ=u�?W�]����=�����V���NB̙�0�S�q�J����+R�{۶m0�L�e�(}���)9�ŋ#��Y�=�;������h���&P��)��h�WZ+���QTֿ��t �#�6Y!�e˖��K�����8z����6m�4eժU�∾��?�E����DDD�
��{M+r�%~���n�щ��C�\X,����t����^|��m�C�JW��.���	%���)+�7|,�s�էоc+(�4o|�SU�O��\�ċ�{Շ���7ADDDDDDD�sVF"��߇˒]R�@y�	ˎ�洴� �������`�Z�b�
��_Y\̀�,����~�7�%��Q�t�G�z�DhoH�]��>\9��@^ܵںe�ΝhmMLu��2ʿ_:co��
1g��8Q,�����˱aÆ^ǃ�M��(��ADDD�� ?��tuw��	�_�/�V(5HȽ���@b�}~��y�(�:�����(���!ϵ��"���h}�-$B����
��3O�y���aԭ�_L�ƿ�uz�=�a���������4e0�`�)A��қ��	 uX���X]��̙38r�rssn�AIqR�ۍ�.�G|c���f��v[�*��͓��z!}J�S/AO+"� aJ�^d���/**�$�]WW�cǎ!�������cӦM���P�+I�U]�x�_=�y��z��O?T���XDDDDDD��uk�
���5w%,�.��H(����.��ߡ�_S��%g�UȜ1��@DDDDDDD�[������y0Z� uXǕ�<��
�mmmغu+���p;�`���1{�l%��JL� ɬ^�8Vww����B�#>��K�#1�ۍ!/�H��J%	qgee�~�P��>")Zy,�3y��w����%KT]9E�OV�J�7�x���M��>~�w@DDDDDD�Ѿ�=xO��}�EC�����`-,���^��)s�<dΚ׹-o����C�
�;����6��K��4���eiŜ]�-!���V8	�sN1F"�P�㭭��ޯ���{�=�@kAA�#����R,Z���nWoQ�d3cܻ��ǔ&F��U� �#ԕ�n�w"���6Zu
��ۧ������L��Ν;�J�.��7tA������u��՟��#_���%@$���Q��oy��޼�����R�mw�}n�3O�R_����-��R�ը���hJL�"""""""�#l�S�ދtd�;aWR�����E���:��ܬ�}~��hllԤ@+��ϧ,��ꪫ�*�J̀��c ��5VpOO|T邠[�7��!?��K �������VSKK:�t"�ۥ<x]]]�;w.W�N'����U�[Ѱ�_�EQb��}�_�fː�������ׂ��@���\]-�6o�>_�Y���*�>��!�5Z�(�����ADDDDDDD�k���"��B���L���I]�ܲ~���&�罹����W�W��`��0:::p饗"##�Ǹ���ci$` +��%>�tA�31���(�:��q-ڲ"h����K:�X,J;y�$��ك�ӧ����_�\s6n܈`0��x��?F�5r;"""""�	4�вi�V^?���I�^r��ߢ��R�ћa�Ή�\׺�	�@����
���;�G��?Cx�I"""""""�Q3`�0�;�N̙���+�ϒ;8���1	Ѻ�nU
�vvvb۶mJ���Ei(����5kJK����fA��n���F�����@�IGR���Ց��{зz�����j;}�4\.ҝ�hDnn.���q��TTT`ڴi �7n/^��[��:�k8�֝�#w�jQb�֭�+�.��ܥY������+��)}�oߊ��{��{��Z��J���DDDDDDDDZ��t�b��$X�(����I}���1�766�*�
��`�|���`d!D~~>V�\�t�fz����(��CK���p'E�����<�	���"//O�����ݻ�'�i���l��a�ee�ܹs� <��u�]�t�#}���}�?p'"""""J�ַ7�_[kiِ��]{#���&�m��~�ʩȺxq\�n�3|5gA��G0���׹e��^xFf@DDDDDDD�Ǆ9��	��l�S`rd��1P����'N�m:t�ΝS2VD����J��+�L���������;::q΃�����HT�}��t�{�z3����V��w��e;��Յ�`o���R�`�]���0s�L<x��q���pWmCf�% """"""�EB!4������y��fC�M����ߪ�=�~O�纞YJ?�/=��/���Co��1m&��\��nDDDDDDDD�hu ��b�OnRx��ə[�4�v��J�}��b�R���vL8F[[-Z��׊���dR��bܛ:���
-���>��	!o"!�WD�=.̟�ky0��M�lw�7ܫWYYY��w�}W	�/^�v���V�X�9а�!܉����(i�]w��US��	�:vmG������uk1�3_�Xt^|�ݪ܍V+
o�5�sMh~�5$��K.Ǽ����]p� �O>�*�TB���(����:�쾿f���������4g�)�������1XlȜ�@���f/�p�����6|>6oެT�����`Z[[1e�,Y��.33j�p�w��CV���
��wB�ݒ����wV���1��i��I��K�r�?�7�]�v!`���TΧ�0w�\�S�����x��ߣ���d��X���W�J��k%�\��P���rwb,��V�m�f�\v��J��9o:��V���ܼ��mx�I�%�9;�٣۾4k�%(�퓨�����z�Q�ӏ)-�q=Ƚ�Z8&W��djN.���Ad�L�p�����~w�$"""""JF��|�7�E*1�pV^��&�fW�݉����n<�H$���n7rrr@4�N$K�r�J腚�A�jJ&��z�A��{�b���i~�H������jns!d%бc�@��l6�Iuo�ǃy�桠� �^�Z�W\�^x��q��7o�=
W�������ҝ�����}	���]Ǐ����Z�6���(Z}�j��5w�}�빧�Τ���������عzhnB�K�v__w}�����>����&����у���>���,k�C��""""""J2*�!�"�шT`0�Y�&�J&D�5�(�	����\.��~X�֘���JiRR�*Ք^$�-y�e˖x=�+5~tv�.2�����{�b�]���.��~��'�sE��~ǵX����X,����ɓػw/�M����rP�����/��p8��x�ˀ;銽b���%�g܇>H��7��&��[\��n���QW���OD��eq�۾�=tU�� �Ɍ������У��~��[?�L
�p�8����`���1��ᜀ��A��?1�NDDDDD�,Fd^���{h�A23�,J�ݜ߮����I��%s��TVV�:��܌�;w"77W	�����-R�����j.��
�}�.
��h����:�&�~��u����E�٬�
9Vo>��=n�8ee�ѣG1a�L�>��d�ٳgc�����wߊ�3��(�""""""�0eec�/Ǿ5�#��J�}G4����<0书�L���p=�Ԩ��O�d���T��h�R�?���x�F��w��M@�â[�Dͣ�Q�1[������z��wQ0�������HFF�΋.�ёJ��ɋ����S�.�� �mۦ�v�� ���ގ���+�v���ʂ!�9�xĪ���Ҋ�yВ�lUJQzb�]�B�0�)�}�TW�ER9r�P42t�7�6��� s��U�.���~wѴ�)L��� """""�ki&~�[8�������y<wQ���Q�ΥRy��k�:W*t7��2t�h�)3S�wQ��Cq�E�'?��	q�DJ^����1�3�P1�6)#��v��d9��/O�{���Ț0�����>��x'��L��JѾH8y�?fg��7Z��ē�{,�����={�(���$�`�x��j����u���즚b�kZ<@����F���p�1��
���ZQ��o�w\��`0���*����<�~�mddd`�J�}J=���WC����x�g0���]͏�����(]~l5�=�3t?�����ٝ�v�9o���:�/D��p>0�����u��un���*���@��z���7�u�
�ɕC�k+���k�G�k/�(i��V�#a2����HY�0���O ���`4Ya��`0�.�X�0Y2��&[�+Bc�'"""""	k��2r�9�!O�~/�	��i�]�|�rL��نH���������o(�n��H����K.��n����ݖ$��}ոM�ƛ^����Ī�%�8�!���똬���l��ω'���@ꑭH�{ｧ�Z�mY�&�Z,����;���\'�>��-��t�-��c8��J�]�֭�+�.
o������O������z"a툞w��DP��#����������wJ	�6�h��l�"�8Y�H`=�pH��W��lμ���YqL�d�r'"]Z�v�t��!"�Sw?)�����ݲ�L3�Y��f��HwL�,dM���s�:w��?�߃%��	��L��s��KO����1ѐZ[[1g��WF$O�����#f�ڀ�&�6�F�3�u,����>LAfO�_�]�Us�y��a�6��صk�~�Rѝ+S��ŋ�܅Tqg��������(g�Ucpo|�YL��oÔ����A�����;�����"���q�+�݇>�^��q�'߇�ɢ��/|�qC���`���@��] JfR�Kv�LŐ��b�o��z��=�3a��/�a����Dt�/<�=�ȅ.DD����jE�݆i+n�q�-���D�aP��[���k8_�)D�h͜U {�4��y��9�~wQ[[��ʡw+$�iooGii�R�zS�z�hkk�wL��Z3*������ �/�u,ԥ}���}������+����RޔH[Ru_����v�1o�<��۴iӔ眬��y��(���F������t�Z:~L�7�q���Qt�'�<ל���k>��⇣x�]0�Lq��Z���s��~�SJ�]��]������\\��� �}%�s�Ɗ@I�*���N��<���d�^��TmW{�T"J=�M��^�Oi�6�]��}~r��dYp�D��f��a+�����-g�2Ͱ�+��`"L�C��˚��7~��8�ԗ��}^>]u�U0�9V�7yy�.���۬:}�<m��&,Kg��T$�C$���Ɖ�����~A�j2jos��1P��c8n�8�:u
{��U���$՛d1��͛{�~���U܉����Hm�~�S�֯M��Z�0�?~6�y�q�V'׺�q�Eњ��p���W�ꎸN��s�^@��B�����:;�>�m[�F$�W��o���4��p��7���+��5 "���6���ᥩFK�߇B!N����DD#';�il�7gF��u��N�4DIH�1lE��&E=m�t4!�n"����8�a�)�%���sw�Jf�3W�/���:^S�1+:O>uvvb�ҥ����&925�o�UQ-���}]5�2@�}r�
y��ގ�3����~�UWgΜ%���ɖ%�"���r%�N�g����mϟp'"""""�y��%�mB���c7Yձ{�RM<c��!��Y����{�D\��{�հ�M���Ɨ�W����s���]��|5g���ȿ��!ϕ��O܏���H}���������~/�I\܉��v""�tz<x���f�cE^��eD��D�&G���%�m!�Վ��!����X�|��H��d����dS&�FiV#S�9����u��^�[[[��~�����grHfM�k48	��9�$�v)��W](Z3Z��ƀ�N�����Gv�ad���yp:����ɓ'c�HRbIEwy�z뭷�����s�*xJ3g�T�)�!=��}e��""""""J���a��g���3�wњ����y
�o��?W�]�q����J�"R�Y�A?�D�1����#�x�6��_��X[�t!�n��?N�4��
���B^�I�@*��\���U�����tu��J��ff��Y��"Jb�	��\�Qz˞uu����*�S�L�Tl��+W�ŧ��@��kii�w,��:Z'e��7�u*��
�������<���ڃjp�䑓���ImڴIy�.\��/5cMY����^��'�#��%�DDDDDD���_��֡����g~�D��Aϳ�"w�5qݿ��at��	ҷ���йo7��y�9;�_�����h4)-1�`�����h�w�w"�Q*��	�_t�EJA"""����ە"nR�5�Nn���º�\�:�
��""KY3������w����w�	J���`�ƿ+��I�Z��&�G�u��	�n��L��=�Nu(�#�Ck���o��p8T��-�����@�';;[���{�)���-R;s���pG$���D��;ADDDDDD�lmAˆW��ǆ<W	�_�a4��A�+���ă��)����b��,�s��������@��b�+wS�w�Я�+ˌ��X��n'"	�ISiR�]�Y�=��{O���hc3n�d��K��8���DD������`�*ٷ���;郼/�{��Т�4�_~~>L&�j�'Ep���DUGw�)_���F�;f�w
y;5�KWƗ����P�~N�:Jn��|����*x����ؐ�{,m{_a�=E�A��n�|wu",�Á��!��e���\���ʊE�-F{���DDDDD4�\���pE��<�n0���O�u[����/��h�����7a-)�\��J�^y5Z6m ��l�a8���'�Ȍ%�!W�t���DDꓠ�����n�����F����˧}�dY��6�EDD��2r�5�J��=>��֦�l���@�Kޛ+++�x�b�Ȕ���z{���1w<u�'���w=`�]��~�����>�l�ڗ��ӧO�R��fSڡC��A	[�G�����r�:޷�O�+�nA����&�<���z�`�9s��Xr��DDDDD46Z�l������<WBŶ�	�՜���9�\�ċ����_B��D"������o�>��K���D�Xm��0�Y��8@�}�cED�rX�]dwd	j���(_���|�����;�N�<�٬��E�N�*��+U���.ܦ��p�@��&sx��ײ�v�cDz�������yS]]�<�����l#\e���� ""J�q?3�"��
?Rj�>��uW�\	9�ݮ�gG������:������7�6'(�1�Ca�Vlh���:&�,2��Yy���J-2�&�pұܷo�M����
PbL�:�_�=�Z_}lŕ��	��k����,¾Q G�v6+�[wT��n͛ K~�f+�����(�"4��ʿ��5Q��������5w�}��g�QOuk����"�����r�-G��Y�9"R��b�������Aty��Ί]0�h�8��r{z�`zqq�Ҥ8�|��ͽ`�~�X,H��yY��m�{	�����F���*���6L�>]��Ϟ=�,����s.���9�9��(�r}�O��n�&��pO/х��]vمŜ4rjWo�>Q��桚v�ʳ�5Vp��u(�'g��#��dkT���ԀR�\2P��Ѐ�G����\  mI�}�����w}��$#��|'�o<��_&,��v���0��[{�T�vQb�֯ń��i�	��[�Ĺ_��P��q�\�]sC\��=sm�oQO��V4�q=�o�o�D�ݟF�?~D��������C�0|x`�n�
�D��X�=��<�H&L��|�f�&�S����@$�"A`�Õ��|���������(���+�N�<�����ߩk�?
��l�2DD44k�Dd�σ�zo���琝id�J}��7oޠ�O��|���#j��(�g�B���@kF����w�������އ����W�z�8w�(=H�]�v۸q�2��d�单�'�X:�nF����ƞ��}���u4
���}?�������h
�%S�_�9GD4V""	���$�=�t!$}�l�ySj��բm�&���CC�k--S�g���V��_c��k\�<ٯ���{�!��Kf:�<��������hj ��b�#�����9�h�d=��H��	�ۓ��mM�8QٱXڔ)S0y�d���hI`D�T����\(���/�z�Z��s�n�so�gQ2�ɤ�^�F[�ߛ�X�+�[PP�4	#�%Uߏ?�3g�(V��R;����d�r�g��Ңϭ��Qh. "������ҧ�~Fe%�;����6�O�h�"�z
U_�!�8�%�n�h>�mrh_!���:#�����9ȡ� N�̸\.Pz��Żﾫl-�p�Be���#������1p���h���/!;m�"�zo�Q�[�!�bL�|Qb�vD���#	�_�#%�Y09�H���������d1[QZR�1��K�׺�q�Eњ;�܋$�)x���3 ��s���{[YD1�Պ��?�����H��L0(+Ϗ�J`ʀ�N��8tȐ���/=<�p{R���3f�P�I�&)-//oط#au�0���_G��P{$I�ʵ'svR�=�W	�Hl7o�9-]�TiQ]]]8}�4N�:�cǎ�����SR+--U
�I5��B�ߝk�܊\ic7"�Dɻ��<�/��WUU1���d��K^}��,���YJM��ݛ��Y���Rh��оJ<%&Gu&��BCk�����Y����^ԡ���q~��֭[��Y*���V��L]w����XW�!;�`f�yL�����(�u��wc�� �s���{�O��T����Q"�������@]r�Q�p��}���@Џں��)%5ox�F,Co����z�<9_d-X��)�㺟��o���@j(���(��S���ϻ??�@D�g������z(��; h4�z;�^H�v��ǖl$2k֬M��Ы��}��%i=���R-�-��7H��%�.��z~��@��˂i�_�rLB�x?x��:���%y�6m�����B�������lE6��#"JG�LdLZϩ]��Kw�k�]���#�b��]z��b�.黨���p{��fUh�y��2�09�@�����$��{�YB���2`�f�A����"����ۍŋ+��itd�̾wIX{N�F��k@�%U�'w(�ۓ��{�ӊ�ɋX��Hcmcn�bȝFc,��Q�S�R*���e�~p�s&3
?�5���������~\��`Z6m@׉�p\4e�s-�ȿ��hx� ��3����)�Ŗ���ta��P��d��sG�s��)���+��	}H�z�̙J� k<;T�ga�8)�l�*�v�uX�Uȣ!x���K����л�J�_���)ǣ����ު������9�}��1�\�D  ��IDATNcN^/�N���G�*�����g�X[�@%Q��_~W����&��0�Mɯ���g�FII	H;jWo�������t��d�#��C����L8����(��Y����\.H?���&[���+2���@##�X<��0��`�u�#Y�]�<�����h��$ܾ���Q��H$C�=�!wJU��<��O}N�KC�[��.�<�K��Yȿ���n�_W��w6�hP���-&����:���p'R�*�\����V���:{f)�v� �VnO��.?����c���3gN�*�=IEP	oK�=چ�jN�E��=���H�]��%4�7�.�TTT(�nP����aϞ=J�}׮]�x��Ŝ�/�2[YY��a�.��Z��Y�;���(!�݅�O��R@����*ܓ�d�$Ծh�"�����T/&+}����~����yj�f����:	h�mp���f��;�f�v	M477��G�M���FَpҤIʠ��e`PZz��J�HЇΣ[����B�6������``ȝ�HU�n�bȝ��0%M�=�!wJE�SUh߹ً/�\�����.�c��m��Z���44���Q�ſ�9g� ]欹�^r�H]�p]�8��ߛ�N�~H��	��5%?K	�ˮ�_|1���<W�Q��ڥɯS%�.׎�{�����X��I��=�2��W	�ͽc�����&���Ç�݋�mۦT{'J	�ɜ�ɓ'��?�jǚ�9�$�s��(Yr��={%�������o!}J.�XT擮��!��:*�:����v������C��=���w���D��䄚`4j[�]��!N���� �lU�q�FeK�)���``~~>{�
���������G����v>�nd���H�n�bȝ�q>�~()?�1�N�ȵnm\wQ��.dL����p=�4���v)�b٧����{?���� "�x�m00�L0��0- "}��'�������iӔ�ҤpR��wT0�����7��^%�#M�ѯ=-�D�F�=����$����Wi��^Z�_K�\~>ѯZ�\��:;;�%s�x�0�|�x�X,�;w����>�P�֭[����+���>���)�����u��N�g�DD���+��p����G�*�)9�c"};Yd*�9JY̫v�v!��v�; L�Z3�2a0q�LO�P�����<�4�hS��{�P.雼�@��e@K'��oh�����KޚC����ނ�O��'�#�ՎT�Tr?���%@B�]������G1�N�I�p{C�j�^}���]����<���[`0�7������;�x�>�J�} ��y�M)RŔ(Utv4�j�(C/+C�Dz!��nW���g̘�+��˖-S§��x��1Iئ��]	�kI�$�-�=[�X"�����H�W�zޥg��|>�+��mJ���-Ŝ�N�27(_{.Z(++êU��&��ݥI�w����0a��D^S�7��3;N�҈����t5�<�e�zn�9{���S�NŒ%K@�%�̨������KQ{[0�W/:Vo��u$L@���>Ԯ�N�Wt�͛7+�X�1R�K7p߿�cRU���02*惴�=�`gRU��o�q�K����FF	�L�p{C�K*�ۣr�T"��_zş�o�s�����p��j���ȿ���O6���@Dj��������V��Dz ��'nWEEE.��r|�CRv��E���@�T\�p���񓰺�n�Т!��U�S]���@sqr=���W�׫45�d1�����g����T�����=���5�\�4�$�.E�v�ڥ�cO�&���ɓq��A��_g����sp'"Қ�lE��O�����븄pkkk�l��sK��+W�O>OJ�Xm�u��h)�����<���ϧhR"*��3�_��*O---- �Tj۷oW�$�=F�g�N���8�
v4t�����|uGa��gǑ�hR)�Ő;��J��(��)�ԯ[W�=^��f�l|D�U��o��qUz'��x�m��2a2�`�8@D�헞+��R4�~��Wǜ��Vi���P��U�e��g�]��K��g5q���A���W4�.�E4�.!��Rv�u��VWW�,(�0��e���*�r��+�P��d.��w�Ŏ;.<�FC�wY\#!��[���;ND�����E����u������YP*MvR�E��x�����T�v��������{�k`�}#�f�;a��ح�0�#��[��C����M*m�%!
��@4DR�\��Ν�����\�s� i#��驖���:eB��^d�Z��3�@=Q�R1�Ő;�T�G1�N��}`��#s�\Un�����5��Ա{;:��s�BQ�47���n��s`u䃈қTng�}d


p��*����;$�,�;��Q�[�R%\�2%������ci�ݙ�<$�.�$�.��`�Hȼ�Tv�&�$�.�%_���N�r�Hkjj¦M��a�TWW�h4�5Iv���|x������4g�/Ǹ�oD���{?u��'��}Ҟ�HZ[[�h�"�Ƙ,��.j���Q�$�~�2��d�"��Ā��D��Vp�֢����mM7n�
z\�v��1���5k��ʠw���1�{Ӡ�x����a��"�w+׋�d*��hhm�H�p{C������(����{12g�AH�UG�>| 4z��k1y��T��߁h�j�xS��D���J{��yYJ��j�Q:�p���������_��.�&S��[����G�����h�]�TfV���'�o�g�Ò�PS	�K��{�@�Pdq��.M�C���<��{�����ǪU��v��q���kJ�]�j��r��\�ɓ'�r��:Xe��(�>��~w�k<xK�.iK���yf��Š�%<'N������������v�2�5黛2�pB�pבHht9C������}I�]V�t�)����NY!x��9����)S4َ%U��]��ٓ��$H}J<����)���;��h`��퇐z��M��+	��|��pJ�ۣrW�9;S�k��|E��]'��ṧQ�n-�-͠�i��zL��?�h]���[�UuD#��ꋘ�����[9%Bs�X�&X�fXl�`4�*0Q���'�'n����W�X��~��1��H�Y�%T3�P�̙Hu�hȚ��Ǟ<�>7�9#UX���������u"M�?Ѱ{Ϫ�2(������o���7*�8��9i�pZ��w����i-{�J8�����^�>��*���>Y�(}��+W����ɓ5��%��wg,�7���Q��ɑ���c=⣮#�����R���]�����%lMн��D�!��e�J�������χ��J��u^+�k�Ww\�cB�����N�1~��(�t
�G]�d�����۵�<�H=C�4|�3Z��������)��ʷ0�o���ף��߲���:�����(���Qݎk�Z�F$@���_�����%���l�"Qz����MR����S����NOdonnV�HC�r�Ƒ�@�b����.MD+�����!�Z�pN���e�L*���/�H;q�^y�%�޷pQ,��^RR�ӧOc]�%s/�Di�����c��?���aY'!�9s��#})��fٲe�G'�����6�E��ٳ��oy'3�E"����P�p׋��HX��tN�*��܅��J����v�n�[�� �Zd�J:]2 %�8-ZsK�t%UO����ՒZ���A���5�C��7����F3�X$"��\+�!l����-����~��\�pw�l�N���Ɩ <NLWѭw���d��P��N��ouO��^A$�׍xI8}4w%$�� ���Ä��-���v]�`4�[a�����9�t$��'n��#J��n����EBd�@��3FFPTF�&%�.i��78O��o�w�߯\2-�J�׈���p8��3����!�������{�ꫯ⥗^BSS�#ב�,��'�{��8�FD�|�.�5�o��^���ك�3g�*����̛7EE\��L��*;i���V�k�$�kw�t���~�`4����'��u"־ڞ="��Wq�[�=Z	AVrɛ�Ta�w �w�B��Ö-[����b�a^^��]$@����:���/HS�x*�t�bm:�DD��Б� Je�g] �+���u~��˔�=��������_��Gjj�NW��D��#���h�Z���z��I�6��R�}\N` ��W�"���+O���QZZ��n�	�^{m�yE	RH�]��[�]~��@�4	DS���=ٹY�����4	�G�{C��k�N)!Yp!siR�]ȵ�z�j�Z�
;v����G�ݻD����
p��� ""�I��Ư����븧���ȑ#�5�;ӏ�����ʔ⡔|���/�[�$�Fe�^_;w�Ax�-HĒa%��B��ŀ�ND���={�t������&[��*wY)7�j9� �J�����W��,Y�TvOW��$�@��w�tw�-�[�=��|�w""""��������Jǣ�+�RZ��EدM��xw���Hv��_����k�Z����K1�? YD�A��k����h}�-�A�B񚻕���H}�5Ga1a�[`���lI��H"���;�p� �̙�[n��/�UKBmmmJ�}�s�����J�]
m����.�ti�ܓ�H�)	f���]LΑ�O��nW�qKXY�SiK�.U���^x�l޼9�=�\Ǜ���4ED�Wރ���Uى�'Y�6c���3^�WY(�bŊ���)�d!�ܵPWW�\=I�wK�	��d˘a�7~�׉DTp��WM�'�.�d����c6ɪ:"����o�>�R���󕁫t#�X���x�
��f���_51��D��
S'd�����]���������ݮ���o�G�s��_�:��U���`/��#]X����*$��5w���Wp��}����Uh��g���j��<�6��գ0?���9�� ���kwO0�ދ��$оf�%dԓTh�@�ƒy��9���J�ԗ\s�*��\���Pv����z�j��{d�PZ��>}:�������^����+�{�J_�d4��?h�<3w�#"J�ɂҏ~��B������Ae�%�'�o���K5�Nꐾ�|��b�\gΜ�w|����u{B���-c;�Dc�w�HDw���}8U�ܒ���1:p�s J�YQO��}@ZUUv�ލ�3gb���I~\�=���"Ц��e��ŀ;�Hp:k��������Mh��Ȼ�a�=�3O�C����}�sHw��?Ā;��"�0j�Df�f�V{>Lf�(}����^d��k�ŪU�P\\���d�熆����
�Tj�P�4��) �^32�,�库���09��r)ת��

.�-��<��o��ׯ�o���"����`�9DD	Sx�gP��O૯�u|׮]�6m����I�h���J���[ee�B�j�E��Y�'��ߜ	�DUo/���z�>�a뿍�H�d`���PD�*�*^���}�$Jم@�����ѣG1i�$L�<�n��{��RG��z�l�L������h��0��$@��ב
\��+������@�S��[P��_�U��XZ�و��cpTN����$BA��e�`0��,��_y"x��v�̱,_�w�qJK{�T!�b��YB��G�����c8�F%:�'M
�I�K榇���9춶6�I5S	�K`^��2����~���'���/+U��n7H�d1�	_�5�0����`�b��Ɖ_�������ۧ�&D�I�\��+W�%?�YH�E�?�U�}æw���#���e�#�o��T��Zf�A��Tp�K�XD	�ƒ\�2!�['N�P��ϟ�T5�
�`g3h�"� B]Ћ���p�	DDDD��$�z��b��FGjnK꯫E�/#�����5���zl��u��sH�ȹ�ʴ�#A퓿�E��>�h��]ht�F~^�2��p��h�tQ���;�p;���`�}��%�.��=Oܷ'E{$l#�4�3%R�,��p����.e��xv�k�����ߗk4Z%��;��M7݄g�}/��"����鄻�DD�X���D��?����^�%�>s�����y�~�W\�,��g�ە	�"}\��ޓ\'�<�pd�"�م��o1Ջ!�T������WkM��'���P�ǎSep�h��5�q�F��hѢ��������]��;n���7�D�{;`���$�5��:��Ą�}	�[�rA��|����E*��Bp=�{�g�3O���̂V�B0�Zkx�����s?��F8S��̴�j5�lɄ͑"J�q������o^�d	���^��J�k	744(� �!�a	Kɮ�D#!�&L��,�hii����`䚮��Q��AwY�q����o�s�=�Tt����� �~0�ED�p�}�	�G�m�Ò�ٺu++���|n�����l��gΚ5K�\f_��������W6���_@"F�� b�]/4���v�<���f]:�&MRZ]]<���z�&��T
�7oV�w��O6m�ɀ�:�>�UM����TA?�����+
>r3J�y �)�UQK�s�WB��ĵn-�?�70���}��=;@��=}R��44 ��)�9�y]'�Ck�.���r=��՜9�!��,'���Ȯ�>��Q:��'��������ߏ����$�.!�������2�"a	�Z;�)l%�9K��Occ� �RX�g�]
�I�ۑ��}�݇�|�#x�g���Y�҇I�3��&"J��9F��kѶ��^ǫ���������3٭f�ԩJΉR˔)S4݅@�#}��ҿ=h��Lkb
I�v���Pb�]?����Ƭ��fE�/�%%%J�7�={�(A�T	Sz�vv�ء^IEwxMf�]M,a�[���B^7�&��k��K���x��<�q��@�ݟB�U+e�;�M�+D�?}��w�R����z^���x��6����f�	���P��A�s=�4�n�#(��g9�@4BM�pw4��@�p8��d���R�o$�~�Q���3f��P�BQ2�'�xl�Ǳی���U�_T��h�ddd(�����D Uݥ8�@�<)�&��hH^��"|��W��=�v��	J%G��\DD��	��O�|�P���-[�`��ժ��R���V2N�b�����P\\���K�]>�����ȼ��H�<m����H��3:���p(曾��c�b���+V���K ��2` +�v���|>̛7O�MFVp��"�'��@���DDDD�^yw����Q|ǽ(��vX����;S�N��ŏp��k^ @+�?��.E��Y1���G��=%X��t�;_WB�Z���#��尕M���o������5h~�e��� ����hFC]��ʸ�Ś[F!�(�I��q��ۥ:�Tl�ꪫzUZ�*��y���N��J�ܵ���|�"l*�����ށ��$�3�.8�2y�d|�;��޽{����ԩS��e5�/<ID�,2*�����W���W�}x��Yt*}�K/��JS���䳦VB�N�8��n��	Cb
��
`0��&��Q��x�3	��z�S3�>�vo�W\q��~����j3پ�h�� ��cǎ���3g�����L��3�cwU��Н���DDDDԏ��i���A�O����� wŇ�}��O��"	�>�������P��C�7�#�I����kP��o���50����Zq��A�#�%���'��h~���+�܄�}�Ƚ��ϣ�T�\�(��]DB!$J�c�a��h���N�=���e�b1�h�"3{�(��5�.s�7�tn��ve�.J�BR�}��o���,a_�Y�p(���s]F�:::��{gg��G��R�]��׈����?�)6mڄGy$f�LJ}f������-۞���\��v�¤I�����t�YiѢEI[���&%{f�p�E]��}K���j�c��H�z{6����a�]7��Pf��cVpW�E5GH_�K�.Uޜe����RV��y^H�����ĉ1e�$�H( �D���,v"""""����`SF&,E%0efjz�ao��z�:ڑN$�\��/��w��ċ���;[�H05?õo߂��5��p��Y��z_���������ӻ����uv �:��ā{V�0�
���k�H��>N�؍�,l6��s�����<�R�^��2���|F�`%��jjj����t:��;��t����4yH�]
_DC�������y <���j,Y��֭�/���)}(���P��(-��Y(��G����{�~�ƍq�-���KY�Z^^�ŋ�R�,0�3gN�l�ZdѦ|����ބe�g�(��<,6E1�N�$W�Q,X���ȑ#�
#��А�JqD=ɵ'���yܰa�2x+U��{�y��k�p���������ǍЩ*�脽^x�D��:~Ti4<�A2�H��������X���w��;m�����̽&s�(��1�^YY�x �gϾpL��IB�>�"�v	�J�A�t����4Y�!;t�]d�Z�����N����������cǎ��`��dr�)��t'�����ch��^Ǜ���J�� �����W�X�dJ���V���ѣ���O�>�����J\qaK��So�놶�n����J���ӧO��4$���T����$�pK�Y	*]��X\�>��ܪ�`��[,GQ����A�������̴�n??N�5�V۸�v+%�䥷p��n��~\s�5�1�o�J�҆zM�y��.�C�V�4i�b�J� d�~Dgg'�?���<�y"&YP��o[�l���k477����F�������x{߳g***PTT�T'Y$�\z饚�)1��,0��xW\�Tz<�^�B��ٸY7|�bv��hu��'����J���F�M�oH7�b�Ѯ(��i2��w�^e MV�������7oV�Ņ&��hЙ!e��0��DDDDDDDDz��q��Nd9m�ZϏk;��#�Y���Q��[�}�ҥx���]��$�+Uۥz�`�R����s!Dzc�ە����C]]݀;�|�T�mmmEaa���eٲe�����SOᥗ^�9""�Q��Lń���O}��qy�}��7q뭷�t(\�R�[�Qꓜ�Y�4�<%}�s���;�Ǘ_.��dNϓ��u\���a����w�Q������%�Lz!@��FD�!������k��gݵ��sv���9g]���]�.vE,�B(�{�|�N"�� If&S������If"�w��y��C�����������CLL��nr���n�e%=�P�^i��wߩ�#�����mmmu��Շ��!�~g"""""""�c��U�ȡ��E����HF�-D�B)�.ݐo���}��=����T������+�^	���v�\tzz���)Aw���Tɔ۫�������L�Pdٲe�={6~��߫j�DDD4p	�U��C]�j�����z�j\x�4�����A�F<dѣ\�y�a���q)`|��!��d��_���1���C��W�hf��<��|��{���9s��,t���/B�D}�A_�v�ڥ�&M����X�=^_բX��3���k��5{�-��p8:Pp8�V=tz,�	��(A}m��&5$/����ag�4�@*�v���;�<��N�B����T��xd~#11�ۉ� au9n��թ �,qG*���婿����9�=�>��C���W��DDD4 -2�������:��$�+y�	& t�K̜9��:z%%%*3�ǐœr�y,��{m�F��=_�����"wp^�k�f�aYYi�)�z3��3f��y�f5���$)0�@�,�8x� �n݊q�Ʃ,O�}��+�<Bg�����EBDDDDDDD
�s��ވ֖N�Ե���¬V����j��E���̱f�@*�v�����;1q�Ğ}�Y���5� �z���.�����2)�&��}�⑾:.K5V� _111��t�?>N?�t��w�Î;@DDD�g��@��y/,s�mÆ�V*��+�.�s�3�8aa,B̤���)S`�X<��%@_VV��_o���w�� �b�L�F�3��WF��rw���ŷ'+�K�כd .++K��ؾ}�Z9����D'"�:�݌n�IKFF��<��3]�w[܄
�Y��ȱ�!A�aw"""""""
��հZtj<٠��d�~\�d��=Z�D�B!�.�c�-��ŋ{��$�^PP��}��2�!U��gQ�H�+��^QQ�F�
��>Yd"RSSU�IwO=�V�X����5�GDDD}�����A�����y���Ώ�1<.�Ǝ���dP�b����*������@B���&��D�DD��^_�[<���ц����ބ��F�������{7��<y����ݫ�h˪xV���"�=䪬�ā��y}Vcc���:�4x����e:�j
��Hh�<� """"""��`2������8p;vt�C���x6yO(�ۥ2���߯:�v��)�s�9>�>-![�LD'�����Jii�
���ޚ��TI�eQ��.��2U��7��v��"""Ꟍ[��]?9�凜����'�|���B���z��t��٠�"a���\�3�#?OB�r�ػh�\����������)>�O��?���}Z�w~��wC�k{�@�k���j���Þ={Ti�F4Td�KN6V�Z�V�N�:u��I9	rG<��CM:��8���ftt4��ю�i���TTU�����~Z�fk,��	j̜�W(��%s뭷���oiiA~~~�s�d2�`�T�&"ϑ�Tb���Tlw�w(����r�YA��������g�y��^~�e5�HDDD'G�����=O����̛��Y�f��ҩE�I�9��V��"!�L��K��677;����^�/���]�1 :�C�F���F7�˞l�&�2��nպ�>\m�m�65``4��,���㯾�J��J����&e��;:k��5�=-�
�w%":���4� 
D��됄�V, 
Tql[NDD4��hi,Eei-��DD�#�����*8m�w�'�� l'
t�n��9��~;�=�\��̻���l}��I���Ύ�D�%NF����j�I��͵��̿ww|�j���y�����O����ۈ���䄏>�?xG���m�=E�9��kr^.��N=�T� �H��$�(ݴ�СC�cPo����μf���u�1f�N��ዀ{�õ�������*���W||<�Ν�N"6nܨ�ݕ-���D���N��IE��=�illt��wϑ��Z���f3�):�DD'r}U>���|#ϟ(�H����#�ڨ��|�Ѕu��"݅���������;a�Ʉ�ݵq��(�{�}��ɸ��{UP]Ȝۑ#G�[�]B=)))C�i�(T�1G��d�IYY���'�������|azz:�{�9��oÊ+��hQ J��~��G�Ʒ]nۼy3�V+Ə��#�d��P���5��ݻբ���s�Ç��߰ar"���<����C�� ��C�F�
��ǐ6hr��jf�yH��d@A��H�	���9�RD�%��ڵK�.'M������~O_�6V��Q)h)ُ`f�Ne�m":)fG�TaȝJw�}T����+j��G��)�H�}f}����3$.VS�1	��ӛAD�!����%��+���ŋUWXQUU�����߷7	�'''�ngq�� �R�]��������r�7߿��枔���n�-[����7�A]]��������/�3oCK�k'���׫��Æy�ڴ,:�Eks���;r���'�+�)�0��ޤ*�G�9>|I�7������{��E��N��n�𷧪:H�WV��y>3f�P����d#2�A:�&�f�J�q�Ʃ�*�TVV�ݯ���1���G/���R�FSL��NC�Hz�ۅ�k�
�k4��& n'""��n�-�-z$�(�s�=55>���}DGG�
�KeȾDEE����hhI7�Q�F������n�HEN	.I5w�VV~��ߩ��;w��>,
����Ǧ����<Y�{?��s\|�����$s&��iӦ�27������CFF�Iݿ��EK�})�˗?�1_3J�H����D��:(h���N���]�v��	{*�n2���d�ON4dRc���jpAV��� �EEEسg�ZI����t��қ,���@��5X`�JAke>��)f4V*#��aȝ��p{7r�)R�3�N���v"""�jn���s;��`�K����[^�`�9���6���@��B%�9.�ܳt�*�*�K��/��B��Kǆ��<�����?���^{��nDDDt�%yF��O��ǥ��hw�MB�|�	�͛���8�=��v�N���=D'K��DDD�0�(�}��Q��ǒ���/������:���b��]��p%r@��ޅk�&��~���*� ���.H�7���݋���'8h��kO�e��ʕ+���)�������dh||�
L	��VU����ב)�Uʈh`r'v�p{7����1�NDD�9�Si[k�'��c�;��� ��AP�@��v�����h�"�;�qL�3�������'>>^�u�{��?�"��)]��ȕtd8�������O�������k��'Nį~���vn """�>�B���?�{a��m�裏�`��A_/�{�t^�p;�@H.�j���9O�p{cc��~��������{a���
ɣ�b�A����ހΎ6xK�!�� ��2�%�.<���D =z��:��T�䆃�4��5(����KU��� �jC�3������&����B=�@1�N��d���r'�p;�g�Ftt��И�@uz��*dL<���`����C=��1	����*)H�̽I��ߋL�����U�N�� �{���믿��O?YYY�4i~��_��?�9rrr@DDD}���������߻�&��+V�P���������;�<f�hP$��{�n�z�����8Uvv������/���a	��k�I�� ��C�Vo���ޢ�LFu��7���S��})==]m���ضm�j�(�뉆�nKEww-H�Q) �0'�A[U!m�;&%	��������C��O�n�Ɛ;��ۉ��<Oo0�h�@��@���������w�lD�߂5�>r�H<��#HHHP_K�i_��{�&]_���؉�( I8N�[Rͽ�����\��c���j��Ts���g�}�?�<>��cQ߆���h-�C���]nkjjR!�K.�DuK9R����g�uV@w%�&����\�;�g_w�������u���ۈ,���j�><D�ŀ{��
�-�U^�˅��d�hUx_�֎s��Um�6mڤB�<i����DF0��=���S�p�3J8��'��ADD���;����ۻ1�N���v"""�(/Ƀ�&�y�0�����Dx�5�~�Ea���*�*����U|��OJJ�*�CD�M����Ts�M*�ʜ�/���/�\�����5
������vDDD�J��c�]���_]���/]n���|�B�;Yt:q�ĞE�D�TVV�:���]w����u�h�ڵ��)ѧ]���(O��tGaC�Tp�*�����jd��'I�@�w���={�
�oܸQ��A"_�hw,)�@�c�'����҃d��L��cAD�I��PL��C�4�n'""���Btv�èw�`�%<D��1�.a�[n�^x��Z�JH��];z!����TUT����V�c�tl��g�ι@��^{�5̜9S��x!ȟ~��>����B��hA�}�!��h8������Vr����dױ���Z�-i�ԩ ���aQQ��p�t���1�_��`��� ����E�vwQ��O�B�S�%�.����lƌ3� �Tt���C�W���Wws2��f����P���*"	��G���r����p{7��i�0�NDD���娬�G�����a�h���#
T�n���裏b��c�2'����B�I%���DU������d����+��¥�,��ꫯ�1��K/�رc��s�ᩧ�R����ȕ�b��>ƞ�f��`���r�������T�R�Uνea�|$�6y>����?����֭[���:�\tߐ<7}x4�aQ (�C����
�]*:\�Hn�5���ǐ��DV�gee��O۷oGqq1���Vc�h`I�2�a#�P���u$:KD�s�
�W""r�!w�%O�ۻ1�N��p;�w4�W��� ��t�a�t���I��1�.U"����T���Pj��7��KKK�����B"Z�������NR��Xr��_|�E,^�			��/�_���ذa���ȕ>"V�ܳ�<��\nooo�'�|��s�L۴i�T�V"_�r�k�.u�w����t�p�[�w�CC�ܴ���N4���*��hݯ�ill�X�]Z'#P�<y��rrrT�	�k�$%/pp��
���t���6�L���
��&�Ɋ�Q��6��|�!w�o�ۻ1�N��p;�w�֔���"��s�vX"��h��`�O�4	�<�jC/�������B��o"
tz�7����y���h4������.T����o���^zI}�2Ƥaܣk��9h)��r���?��3�t�M���H����=��߯�>p� �~�m\y�عs'��X���?�PT���OS�h�:�D�U��Ύ6xK�m
\ެ<V�\ڧY,U>X�3FmG���ݻ�*�y��ശ���$����hFĘ�Q��t4�w%w�%�#τF��>D�;��7y3�ލ!w�6�ۉ������0*a��w��u�j�����U0��gϞ���KU�V�yyyn��d^I��k�(":�m۶�J�W]u��\�t{x���1eܸq������?��*�GDDDΤh��_��g根x�������/���V��y�6����/���X������&����ڡxz0F�Ak�L1d
m���т�&�܍��q8�[�3�i]�gÛv�=���d�Q���R5 !�8z��'꯾���eL���`F���h8�-������VX����x�@D��r����c&�'�"�ލ!w��ۉ��<OB^Ņ{��hE�̿i�0����`���_�x1���j�yss��,!��L&��>Qh+++���?��.�&Lp�M
˭^�EEE*�w��� ���>�
f�3ct*�>�9?���#;\n�^@V^^��h��y��ڥr{ee��۷wf"����hk�PЇEAo��'0�b��k�� :�w�w���z�>�T�(..F����s��EMM�l٢�f��h`���8�{�a���R��殭�~��:��K��!iWDD�M��+3�N��p{7����n'""��6������A���V�"
T�n�j�R����̻:t.��94)����D�M:;���*%!v���J�r����U�-)S��_��=�**8�@DDԛ������T!������g�ʕ*||�M7q�)yԎ;�?�	---noO��0R��9m�h.܃NG|Ik0��"Oa�=�H��ۊ�\_VR=B��zӎ��F(����f�RU96nܨ��DDD��?�R�;��\1'���jG���:�JZ���I0DpE%�����"�ޭ;�.�ض2�N��p;��57ף(�0h��ނp�hu�I��-�.�}y�L�4I}-!���|U�X�{&$$��IDD��1c���*�~�W8�1��C��/��"���Z��;�.�"""r&թ��d5r�u٫��G
�������oWR��/��믿�s���|.��_!��՗�A��>{~����h�ؚ<��㋀{b���X�]*�ˀ��+�
��>c�U�cӦM��m�̒��c�`�J-Y�k��EK�~4��:�^S�p��B��>D�gr���p{7	�_���r��`��������*QVr ���k��f�v�ه�	9"
L�n����O ##C}]RR��ޤ»TmgQ$":�� U?/^��d�A�������\s�Z0�_�
�?�8���"""r��Fb�C���7�r�?��G�=��3X�|9Ǝ��������?��W_��]�3`��?!�����â�'���� �z_dS)�0�b�*������I�ѣQU����(��555]�&??T�ݤe\VV���ܽ{7�����;�L��boa#�@�AV2J5wcT�
��V�KYo?(�1�0'��:�d�m"�_��@�C��C�4P�y^}]��p�M��m0�"a�W��D��-�.�`O>�$����<Б#GP]]�r?�ժ�#š��NFmm�
�ϟ?�'Ov�M��/��2.\���D��F�y[�n9�Ly�+*�Q���n���Ѐ�����7o��8�@�QYY�?�����s{�><#�~����.�#Gk#:���Mƨd�\�<��P��&�1����䵇0�Cn�jd�
�˅�'�����с�	&�m���j��f�I�(//w��%l� ��5���>��B(-��V��u�����0Za�N9���AQ"
�S�S��C��_�y^cC5�sm:�a4E�jK�x*Q sn>|x��������SO!))Iu�ywE��v��ܮղ��O{{;�y�TTT���s:�"ko��.��"�P�?�)�{�9�_�DDD�K�{hʢ�`������F����.r��b�
<x7�t���At"۷o����7�H�s�d޿��̾H�������ltv�y�yJ�xCd����$� ^�ˁ1�Q����e�M.��M�'H�[�QH��ȑ#�VTT���l���y��9>���m�,���%yl�6�uh�-Q����oew�V��0���V�l"�@Ð;��wcȝN��DDD�Wh� �����H���lD�m]_�B���j�p;Q �+����RRR���O#&&Fͫ8p �ͮ�O�krrr2��J΋֬Y��/��r�L���d~��?ƹ瞋�'⡇R�gW�Z"""r��L���� m��n�s�N��u�ҥ5j�ܑ��7�|S�w�+b*���@�=oC{��`N�梜>�@iMV�Ↄ�[�zAZSP_���(���R��S�2@)�w�&WR�C���2�2NV��FPhs����Fq:��iԉi��ig{:�k�hn@GKm����g5�F�����C�7Ag�:��w}�A�g�Z"
����s��C�t"��X�A��"�1ş��4�W�����2�b	O�F���D�*���ÆÓO>���x�
�����;J�]�DD��w�^U��k�ADDD�~	�K ���	g�q��^U\������7���~������OUU��2{�l,Z��EKɉ,<|�p�ȑ>�?���Up�dI^���֊#���s�(	(��[x�A:��ۜԅ�Dmm���~���j�*���1�~��h�ܹhll��͛�>��
=2�_RR��6n��04	���c�pNbQ�bȝ�	�p{7�ܩ/���#MU��X��;���B��Ip�:�	z#ۂ�`�K�'�xB�K%ܾ�~���:�G�ժ|��7"���9�?��O*䞘�س_Bw�6mR!w��|�rU��> �2�e`�cp请�|����G�KW�\��-Y����H�&���K���[hiiq{�9�o~1g]=��0���hi@�
#K�̔0�_!{��`�=iu���g���0&���}p�i���WVVbĈ{�ݮ����#WV�3f�P�����ޏ]�O�O��K��l��Q�bȝ�H��n�So��<��U�]_�Xst8~G��C}m9��v�3ZN�ƙ���_�T��	&�?���ˑ0ÁT��X�A��,bDD�"�إ���ŋ��,����V���>n���oŊ """WZ���
k���C�lw�k�*��<��ϟ�����+����r���j�C_,�1���aN;��2Ŧ���GK��tB���Z#�M��pE�&+:����L8��nY�-��fυ�bccQXX:9�  ++K�n߾]��a�����߉m�� ""
d���p{7�ܩ��DDD��ц�%oO=���j�`4Z��-a4E�������_4���c��g?��
�����]��2�����B�DD�$ǡ�^z	�]v&M����k���,7o�-[�Bx��.���Ƚ����3p�נ��}xY���j���~�뮻�i�7�ھn�:����}Vm1g�×�/����?����F��0{@ő��?BU�'��C���݀{�"]�\콺L�III{i�ƀ{�ɿ˔)S��999���Gd$'t���Ç]�c���8DDD��!�����n���DDD�s��)��}W���-�5L&ۡ�[��AD�%��홙�x��T�]:�J����9d �x����]*��<E�Co��6���1}����r̕9����^z)n��f�z��@DDD�eLń�7��K?B��?�y?y���/~�ٳgc��0�L��%��_}�Uս�/:�î�/�θޣ��1�`��@sɾ~�16]=/"_a�=D�b�&�4��}�#2��WTTx4������fcƌQ��:��Sfۛ�"+�JKK]�GM�DDD��!����n��.�ۉ��J��Yשv�`zԨc���Ո�9Z�CobWK�@�� �������W�\���s	�K^	�sΆ�|M��~��Z|s���w��c�����q�%�`�ҥ���G}"""rO*o_��/Aޟ��������Z���?�ƍ�p�B�y�꽗�GSSV�X�U�V�\ۺc�x>2��Ƙ4�<	�#��Z]t��#�E"_b�=D���ʅ���,6d��b������ho�
9�{�Iw�o���j+**Bvv�T��Y����=���""�`{h	�p{7��C��DDD����_M[
�*�jq�675�����2Jf0D������D�v)��O�Nݕ�{��v�
�3�BDCiݺuhnnƼy�G2�(U�%|w뭷��HP�����u�"���¡�ކ�-��y?�����Ś5k�x�bu]@�M2[_�5�z�-����y?�ъ�����o�_�>'CT2��ho�9�}�]�5��A�kL��(�V�B���^}��mq.��]YY��x�����Tˎޕ-h`d`U6�wڱc�F��(p>|�e����s.����C�!���r�y�ކ$���kuN��a���p���t+�(0[�=66O>��z�R��]�=22iii��_�*�`�0�Nw�K�O�=Z*�Ο?��s�*r�v�ZQߌѩȼ*7��_��jK��������3�`ڴi��6&�ճ��}��7���	}62����L��1.��l8�Z���!2�kK�P`�=�I�uo�[R�p��z��d����˅tBB�j�F�#��3g�T�C6oެ�Y,P`����S/�FǷ""
N��`�wc�=�1�NDD�͎vj��H�s���������h� "�l�vy�P�9-	�J��w�&	������ȟ�ܹ---�ꪫz:��1Y:���G���q�}���;�'""��>k1l�.D�k���/���~RHvÆ���T�K�s��?	�K��ݻw�~��($/�.�K�×�H�)~$���·�I����S:L6�0��Ty7��'`[N�K����J�u����hyc'ϲZ��1c������6�,���|�����:}!����Yw�����P��{��p{7�܃��DDD�u���-1�8���ٮ�57��b9ڥR�5������Z��U���P���m6���.te�^��R��XR*11DD�(77/��2������Rh��O?�\�Gy�>��	�\DDDt4�<|�u�"~�2�\;�\�_}�fϞ�9s� <<�$�����c�֭��1v]�ƞs#Ү�%��*Z���ah)�s�o�Jf�vr��0��
�΀Ύ6�>΁v�J�2)UܥB����fU�B~.y��d��g���|�oߎ��
���������烈�(�I��f�܃F(�ۻ1�|n'""�c&	��0l�(h�BLkZ[����h�N��uhk�E[em��m����z�ȟ[�]��J�]
BI�������b���A^^^y�\{�=!w9Fˢ�իWc֬Y*������0MDDD��.��g���˿"�_?F�q��ԇ~���R�T�EFF��^aa!>��|��7',�kN��� ۄ9���8���Vw4wi�N���\'�@1��$������ag�С5HOOw�_RR�р�HMMe��d�b�����0�S¡C�\�GO�
Z����(D0�B1�ލ!���p;��i�B�o��wU3��:�Z��_[�]�����#��KU���8�{|��W�*�˱zϞ=�`�Yg��'�x>� ���@DDD'&Ej�f/GT�(|�q�~�t::��KK�
��Y�ӦMS�庂|K��r��g��6'
��mqH����]����5����	��hl� ���WB>狀���ؔ]�p���Q�ʤ�DDD����l�1cƨM���&��e����TQ�V��Şs���B	C�-����r|�yW�	Ě�&th5'���v��p�X�|9�����ޮ�Qz��K�v�ۉ(����/��*�K�]��täI���c��J���� ""����ư�~��soB��?A���{Y<�v�Z�[��ƍSA�	&�k)������o��矫°'"��y"��{�5��/u�f�I��>2�G���'OyC;���:���z��K���T�c�$�ܶmȷ��lG�Avv�
����&ߓ
���3�9DDD��!���p��r\�y�渷�lp���
"z�n����1o�<�m������Ɽ�q|<+�Q`:|�0^y����?t��~�zX,dff��G�O~���DDDt|��)�|�}��G�돢v�ǽ�d����lr�1c��U�f��<���D-&ذa���Nx�ވ�9�"������~��v�3L��8iu�5G���֫��y6oY�Mv�_\\���4���7���HTWW�|O�=e���Rd�~���VCC��U���ިV��"����r<�=����vq8�"j�n�@���_��&mjjr�=66V܉���^{�5\}��=�Ϥ��g�}�*��?��w~��_z��Q0��c~�Rܥ�{}�~��}뭷��类*ӧOWU�u:����֭[U����ܓ:��-������1Ƴ��B	�}X����	�*���_*UTVV"&&ƣ�'����BC'**
�f�Bcc#�l٢������Tow9��hs�u ""
e����Ɛ{�`�����wz����܉�R0��G��{�G�<�M��~2����"�`��~������+{�sv_�b/^��H�W_}DDD40��a��z��C���@��\Cz�NR�ْ�j����ԩS1q�Du�B}��S��%�ڿ��;477���i�ማ�I�>C����w�.,
���^_1]����}.�(���<p���P����%'Hg�}v�j6�P�.9�ڳg��~�)��""�Pǐ�c���r������t8ZLd��q��DC-�퉉�x��GU�[��XQ�|]`�ۑ��
"�`"���.\���c�?��O�x�*�.��U�V����.|�dvmM�;Q��s���t��x\C
�~���j���Ĕ)SԖ���Ӆ%Ե��!;;۶mS������^�=�snC�wA�׳D��G'�F�����*�ذc%�_��{UU�
=[,�>ވ#��f�3�`4�����7mڄ��Zu�D�!�ݝh%\x7����(	��Ty/F���П���Mڮ��TbT+��'"!�+�� W<{�����WW�\pMDD�k2,A*a�ɏw:�����h�����p�`z�����GMM����n��l6lXϱ��(��ر�����9���W^y7�t��n��g��� ""����ND�-C��F�g���/����b����j�^�Zm�כ0aN9��;6�\�-ܽ{�:?��R��?�3�#~��κ}�-��`��Y9�퀻�g�DKK��Zq���B�9ң�%o���QZ?����g�q��<''���`���d �7s�h�']"""���с�*�@����UՅ """"g���ގ�N4��&�`�K����WsS8r���~OOOg������͛�9s���kooǛo��+��?�0��>�����������<��+�@��U([�<��{�����~)J�q�F����$�3F��%�'�t�I]]rssU��rN�ћ5u.��g����wRt�H5���j�ѳ�n��s�N����T��ݞ$?S�?J�?rB$�T߿�j��ݲ����L��{K��i� """"""""��$���ா�������|!��bɒ%��z:t�P��'�V+��D2֮]�B�ӦM��WYY�/���g��O~�<���hnny�F��m��jk)=���F��W�Z~�_?���HmR�]��ƪ�{FF��n�����+�J�]ɥ8p@}t��:)-"ƞ����S��uV;���p'E��t;����@Z=�7��<��)�,�|��(�tO�j2`�o�>���� ��5����<�ߎf˖-.�dK��@DDDDDDDD,z�DU���>��T���
-�D^���s�=���WU������nR�I�X���B�'�|�:W�n{��UϦN��{�?��Ͻ^����(��G���5��B�W/�|���V]��U^^��o��F}-�pqqqHMMEJJ
����ޡ U��9JAPɞ�M���.<K�8DM�bϾ��� "�b��z�#b�p��9�l��:�N��_�X�O��y��u��a��ւ���[�VUU�m۶�F#'��C�He����[
�9DDDDDDDDD����m�g�Q/�n��ᮻ�R!M��
��d�kĈ�`LD������o���:����o�UA��ӧc�x뭷@DDD�cI��ԫ~��+�F]�jT}���~�֊#�y�/9<�6o��t�,n��;Y��͆��Hu>`�X�G��fsO>�w(^����ڪ��Au}�������=kjjT�����u�6|*"�.@�i`6D4tp�R�]�3�S��86l*�#��~�fQ\\�B�6z�h��:�UY�r�3k�,466��ɉ�ئM�\*h�F$\p7����������Y�1���FI����
*��`�KG����*�QXX����w���Ṙ�(���k���%K��ʮB�l��>n����� ��$"""��hu�M������oC��Q��}4�����A?��e4Z��f!j�e��z)�Q��.��0�N��h`��E� ڑ�WC�\���&��???_U��t�F	G�����lM�KV�͘1���غu�Z��*�}���������K`�IQ0�t�h���zt��}B�tf���Q���e.���S�ZR=��������T�iQȓj����*�.]�sL�����<���G�
,��T&�-i�#h��@]���۳u9k�tx�G��Jk0#l�4���B���>�Lh\�L�p''����Q��rc&�w�/Af�p!�~�&w\<�z�ш��,59�}�vTTT�v6��o�q�ޮ3 �҇ADDDDDDDD����Z���"����� ��.��M����UW]��.$�)���������" 	��t�M0��ّ���{�]v~�a�I�w"""�=�F��Hm���u{ס~�Wh��ܵmA[m�.F3�e��1a][���6�Lr'"�ǀ;9��H:�M�^���yؾ�SL:e����*�Ҟ̓d�t�رزeK�@*�7�<y��<''G�V"##APC>�?n��]'j�ADDDDDDDDl���~�x�@� ���=�������~O�2�/VM�z켓�[H�����'s�o��6���J�~ ���U�3�<7�x#^x����Y툜2Om�Z�
Tн��4ف��\4�샣��Bs�h�����<N�%خ�kP�Pŀ;��G��$ஷ'�˽m�t�����6`ذaL�ժO���
lcƌQ۾}�p��5 .��B�Tm���]��z;3}G'�ZZ{��6����hyV�.�ۃ!��*˜��ۥ;q���p�Q���\�޽�V���ٳ���ްi�&u�\�`��}��� """�c�JQ[䩗:�o�.:v��Z+����VS���BU���}�c.�	{��)0�`�N��:Ƙa0'f�`�d�(�0�N.��H�����~Ś�1�y�
�v���R�;11F�@j�_rr2���PYY	
|�F�R���A���0���uh���Eyy���ؙKX�����������VZA%�cǣ��@��-�ooAkS9**��q�è=��B�#�T_�``�FC"�n���F��P�=�ܣ��%%%����`��`Pś�+��5k� >>'NT_˼�+�d�u|=t�*�GDDD���������y���:8Z��t4���֤���h���9:k$t�0h&Q�	�(��F�pj�������5�L��p��--��533�+�;z�hl޼٩�6Y!�,^ضmL&�WH�y��w.��D/e��@DDDDDDDD�:ێ���ZDh͈ЛP�R���u[{?~^��}O����9��F)0S�]\~��4i���PZZڳ_����<DD����)L'��7���W_���=����sGDDD�Lջ6"���(����C[u1:{�v�Ǥ+�f�K�5c��~�|!�R��Ӥ�����}��������Y���ب1tvv�j�"XI�����eҥ��DDDDDDDDD���z?*�6����ddd�q�` �d����������j��[JJ
,�����8���˖-��HG�u��aƌ���k��/������B��F��>"m5%^,�ņ��qFC�S�]��߯*axCDD�X�Ǡ�#�v �
�[�nU�w�7&���ؽ{��~cT
/�DDDDDDDDD��ӤCks�����uU{�T_"�1�#�n6����
�P������M����W�����o�?���!U�w�؁��4,Z�H��J�n"""""
]�S��x�ז:U�����p�oq�E3����Ԡ��qqq^y\�___���Sp2����R�c�����nG���g͚5n�>S�zZ��;�Gj
��""o�*�R�]�d^��ۑ�&""�?Y0����.P_�t:|���X�d	��^�y�N�\"""""
-�S�4z#taQh�����iu�g����5@x,����R����T����/Y�?e��yNN����@%a}��ޛu���9�Z��M�6M�/���PZZڳ�`0 ==]�?���_����?~��Z��o��6~��஻�³�>"""""
M��q�	�	�w�������Oܲ�9���ڊC�a�ȑ^y\iy6a��欹��ƌ������MP�� PH˾M�6�ޠ�"��߫�DDDDDDDDDDD48��Ѹ���p8p��ឮ��LKKS!w""�w�}��񈍍U_WUUa��͘>}:fϞ�/��DDDDDzp�����[�ho�����O�_}�.Ξv�����BuAk�۽�2 y�)���{[[(4Ȣ	ي���{�n���y�S��� ��U�����r[��[�9DDDDDDDDDDD48b�����¶���ܖ�����p�������_�ҥKռ�����1˖-Ss����)�GDDDDD�ÿ���Q)>��#��v_&�թ�c�����N�Z�m�ٌq��a�Ν*DL�#11QmR`۶m0�L0��G2�SVV���������ADDDDDDDDDDD�w�b��ɨ��u
V�l��*�DD�%%%���O1o�<��N�Ûo���o�w�y'�x�	Qha��NHk�@���*�<��+���_��7�iSS:����=�T�?~���͐{艊�¬Y���ب��I�Q��
!���y��~�F������������'::7�p���+�ۻIؔ���}��wHOO�ĉ����z�ʕ�3g���s"""""
��I1D%�,����`۶o0y�$��


��cx���ǎ���lp��#��3f���7nT{w�5i���_�]xa�r	��X"""""""""""�[o����8x� ���{�����`0�������Crr�Zh$����	�l�2Չ���DDDDDp���5���F{}%|��<��߀��F�
�8����i���ڒy���333�w�^P�2��>}�
��ر���P���/Q__�_��_�G��ɼ�Yg����J����쏍��b8DD�N
����;�����jնb�
,]���v�|�IQh`��N�12U>�jnʺ���9ܸ�B�����*x>n�8�>~BB��`�@=+��6yL�<Y}.�iG��߾};����ޖ~���
"""""""""""���0,_�mmm(**��o6����""�Çc�ڵ�9s��Z��W�\���?_u�^�n�����(�1�N'Mc0A���2�<�ވ�1��n�G�q�4����Xii)�������T�yϞ=��7ј1c�&��}���������B|��no�9�ZĜu5�����������h�,Y����@GG�ڧ�h0l�0���3�n=b������e^v�ĉjҖ-[��� """""
n�S�"��.U�;�}�x��X���n��r+� -�W��d�?�w�fȝz>\m@ߵkl6�z�R��_�}�I��a��DDDDDDDDDDD4x��;w.jjjP[[۳?))IUp'""ߑ�ѷ�z��z+L&�Zd����o���_�����7ܩ_4:=�Ih�8�Ǵ�~%������9N�1�r��O=�T�t:�>���(5�)!��v߄�)0$''����۶m��`P�,�%��O?�T��]h�ȸ��ЇE������������G�������6ݤ�Rll,���������'�`���k��Y�]tV�^���lQ�b�������28ښ}��N��~�λ�馦�&���
��f��1y�d�on���N#223g�T��͛7���V�u�?OgJKK�ޖ4��`�����������h�/^���T��磭�M퓮�������̻�7����k���2e�Z�t�=��8Qc���O��1&�Ź>{H}Dr�.���ة���t[EE�p�� ���b�\8۞����Ff̘���l٢�R�?����۷��m��r� """"""""""��KLL�Q__���ʞ�III��;�+V��n��bQ����k�����û�"""""
N�Ӏ�,6�v�7���1-ç��r�R\������.hcbb��<�b�)����{����D�ȠwVV�jg�c�����*�'�g�l۶��m��d���F�ޒ%K��ρz����#**
DD4����g�}����s�Nr_�v���$"""""
�Ӏ����T��N��3������_��ˣ`2�z�wvv"''�'OFXX�ן�V��رcU`Y*m���#�y]
y�J�����rۺu��ަћ0�GoBo�uqp\��gҤI8묳P\\����O��}�5���N�t�?~<F����9�1c����o�[Q�a��Lc0�����>��s��Ko�K/p����C�Ԟ2e�S�ݛ���T���ۭ�� :d�M:���ݮ�EUU>��sU�ݝ�~��g�������������hm6��V��5��J�d|~�ҥj~G��vKHH��h�)8�b�
�q��-���?����S���iP��7T�����Ԛ�P5�f���+�l�N�� ��ݻU��N��#!�SO=U]4WWW��D�����"�ڵK�>�裏�\$��;o����������{��f��\���U�����5��������Z�
^x��Z�cWTT��[o�����g!1"""""
L���h40�Gsa�Z5�+Ƙa�n��k�`�3�n���W!��'v==�o��шSN9���8x� /��$%%�f��?��?�����1�:��#""""""""""򔰰0\{�jl���V�9���T��-Q�}��7j^>99Y��"b�_=fΜ���DDDDD<p�A�-����VS��ǵ;_�@̮]�8a��mRI=;;�ƍ��@�\HKE�={����wU�)0�������QPP��v��S1�A�㡚�����������S/^���H����싋�S܉��I����{˗/�V�Ess��g�>࣬?�o_���0B�
**�ZP܊���j��k��{;���U[�*�։Z�*V�����;�����{,T�$w������.�w�<&����}V�݅^�7�|�:�
   `h 5�~��(T��I�`t_0&M9V��~�RS�T\\�����֮]�����SR���o?+��i�&�ܱC�@@7�|��7�#��S���]N�        @�0��Ι3�:����i}ͬԛ��+ @������ŋu�AY�/Z��
��x�z��G   `h ����pʗ=Z]U��D����C/�_��{]��Degg�{�ŭ��]RR�cں�eFF������*`�`0�[o���0�JL��o<+oV�        @���K�sG���[�xĈ��  ��K/��ɓ'+55պ�~��5w�\=���   ���7�iړ��@Setw�p(�kt��_���[�򏫨��Zԣ��n�6�iӦ����js���b˼����������4��r�-Z�b����&����Pb�T       ��3n�8͘1�*H�z�Ƅ#�y ��aι���:�3��W�^�C=Tg�}���.   ���_y��lQ��=�;v8�x��tǓ��O=�z3����F,B�ͽ���Zڲ���
�G��1�cǎ��]�ti�C�����ӟ��U�V����W�yT)�        �_�w���j]]���9�SPP  ��c��N�>]�G�����5g�=��S��    /��_�|9c�Y�B�p(��v��;�:��������)11����"ִs�7,���v[�꼼<�_�^MMMBt���[?{Ө�դI���{�Y������C7�|�����ˣq_Y����        ��ĉ� �ƍ��b��' ����3���+��V�6Es---:�st�7
   ��F�����ɛU��ڍ1ٷ��u��?�g��a��4s�71͋�X0!����
�oڴ�z������l�������{��
���ިo~�&ܾe˖~��ti�P�~'	        �?����ٹ�)&2�� ������:������}��Z�`�N��   �c@����hVO{c����&*r�wt�t��G[!珫��ײe�4e��En��Vq�566Zm!mmmB�HMMUQQ�233�g��׭[7`�RYY��n�I;����֘��Q挹        �Ϝ�6m�6lذ�k���1=O �/���u?o���$���r+�����V    /�0���
:vE}�O���~�ÿ���]й���j�6/t�^�bɴ��ͼ�޼y�N����`��Z������x֬Y�[n�E;����S��)c��        ô�������������p�W ��c��.Z�H�gϖ����~��G���    N�1pN��J�U�R�p(�����x�wu�ӿ�e�OWvv�'�oB�K�,�B�ny��6�b�`5��kkk����t:�߭	������m���X�g�_/^���_�`p��w��Tz��J��8       ����~�i�������}����
A ��w�yGx�U���٩��2�u�Y�կ~%    �w(��/o�(u׬WL�<J<�����4bĈO|;XM�&LPVV��ARR�Ə�1cƨ��FUUU;m ��sf�м�<��{vWf� �4i���}�����m�I	O<�.\���%�k�7�Vr�!        g޼yV��)�1���v�0 �B��^z�%�y���W_}U��F��M�6	   ��C�Ν��pZ���ձ9 �KI��N�,�CgLi��ɓ?�m�bwŊ=z�F��x��x�@��ZZZ��{}}��3��n&"�f�tJHH�&,_�|�oô�u�]Z�l�N�x��T����X<U        `��6_�����vz4�9 ����?Ԍ3TTT���.���3���~�;   |�#*�#t*���p8�z�z���T��?�O|;�hÆjnn����������Z�9���F���Zaw��L�===]999V�ݴ�s���͛7��u�u���ug����kOZ!w        0�L����u[{�9���� z̹�_|Q_|�5����_�\���竲�R    ��J�b��}����ʕ
�cv)����׿�����)sfo��������V�{bb��y!���im�pXMMMV�����>T�	V��\��{��e�̛��gk�[o��x@�@`�cҦ����&��eO       h�������k�Z��s,yyy ]�6m��ի��;������SN9E��v�    .�5�[��q�X�H8v��cgheb���W�y��^�'����i��KJJ���N��v7�j�ۄ�M}KK�g���ieOKK��S̖���c1opO�8QK�,����,fR���o�%��kU�����x��        g��~�u������ܜO��9! �����/[���y�7�xC�{�~�a�4   ��A�Q����7!����a���/Us�u�q���p����C��5�ۼ�5/~M�x�KHH����B�sx7M������vk3�_�f���߄�͖�����d��x��x4i�$}��VS��lܸQw�}�jjjvz;����sԥ        �a��|���{��9���+ ��WYY��+WZ�{�9���j�|�ɺ��   `����.��?Y�������p%��5������5gL���g������Y!�	&X������߰5��&�n^ț��n��|gA��a�(6-(>�o۶5�n���fߙ���;v�ҥ[����O?�g�y�3fެb���J{�        @�� �Y�֜1����r ��`Z�ͪ����E�t�)��o��u�   ��@�1�N�T��[�Ɗ��é�C/ҳ�^S��u�	��.|m�ߦ�{Ĉ=z��@>X��~kۑ`0����r�Ǧ�}k��|��u�4ڛ���K����P�PYⳠ����`f��������5��L�>s4��;)C         z̪��wܶX�y��� ���|�rM�2�Z񼣣C�{��|�I   �#f<���l����(i��Z]W�?�{��?e����i&�\__���R���k�1�%f3����q��Y!��\���?����8\n��C��mSc/        ]��U�c��� 0<���+�<y�5��4��w�Rw�l   `�pGLy��������C�7{�t�Ou�k�q��u��l7���KK�.���M��y�C[[[�����f�ݗ3Fc��_�        �>s�fΜ9����V��� �/�X��Ž��AIII����x�b   ��s[�|٣�pH=͊9�[ɇ\��6��?��N�-�߿ݰ��J��Q�TXX(=&�^VVf5��|>]z饺馛v8�?��5��[��'        ��QGe�»r�J�s��NY _���ڶ�E���O&�   ����3!�ܱ�T�U��U� �h�Zs���'n��Ss���f��֭���%%%JN&�<�F���
+�����I�&�N�SO=��k����J�~�        @l�����z�B!9egg 0|UUUY��Ǎg���5k��R�ƍ    �pG|p8�����5
u�)�6_������g)%%e�q---Z�d��&�1cv�������I�ׯW{{���'Zov,[�L�3���?ʓ�+        [��)$���n��=�  ��믿n�M��io7�f��r�    �7��|V�}������P����Ա#{t���p\]]����k���M�����U6lPss�g�ۼy���)*�ړJ��D       ��p���[E6�`����v �a
�L{{qq�>��C͛7O��{�:;;    ~pG\q8]��W�ir�nW�px�x��R�J-��#:m�����n\8��93a��#G���P.�K�O&�n��0>�it��ǵ*<R9'� Wr�	[�2        @ly�^q�����>7+�&$$  ô���W(Ryy����p�B   �_�w��{�xuU�S��E��_0Q�y�ҭo>��=o���Sbb�v�zzz���񻠠@EEEr���/��#��^{�5=��-J9���o}=�Tw�&�r�        Ė	*�¡�m��� >n͚5����J�/^�9s�p   ��[�'�S��q�Y���&��[i^�-���Gt`z�fu��vC��-[�X����l�G����F��a�(�y���_S`�i�9������ �/Y��       �ؙ5k���뭏�~��� �V��lk�����
��7Nk׮   ��D����/w�T�A=퍊7��T%��W_�e�>�c&fj�����X��n�M�ڼX1b�������USSc-5�����x�;zr�?U�1]Y��^~�w�c���%�n�.       ��Q�Fi���Z�b���9 ������:�裭��|�M����    >pG|3!��1V�{O[��7�X:�Z�c�b=��'4k�RM�2e�cMغ������ӕ��o-����w���i�7��`��;yz�����c����>�cf��U����pqw
       @������fkU]���9� ���A-Y�D�z�֯_�.�@w�q����    ���D��B��t{h�T�J{�Ի=��}���3�5}�JKKw:�����̛�yyy�ff�c��	f	Rj7?[;L����^�Z)���*+9s���Pw�z��J��U        ��i�5��YYY�
 v����A$��e��n>~��W    �pǠ��(���S�n�՜�F�P�`�b���Y>e��N����f���-[�-55�Z:�l�MY���-�f������Y-vTTT���^�fo�2���r�2v�B��
4Uț1B         :9��|J{{�l��ܵ ����ҢU�Vi���z��w5s�L�   @�"��Aŝ�%�۫��u����c%q���ݞ�������f������۽�v���̒hiii��͵ތ%��I[C�݄�����-]�T��{�j3�Sڱ?W�?�_�)�T%�/I�D�>        L{�9W`���: �����
����j�����[K    ��������_8Q�Uk�l�����I����Z���B���a3���;c��MMM�fGRRR���yq����ᨧ���y444Xo0������f޿��Z�	��~��p���_w�F�o���        ���dk�5k�X��� �cÆ��fs�ݴ�y�z��    �pǠd�VȽf�B]m�)9rx��:���*����o\�f̘!�ӹ�뙰��f��7���+==�
țK�׫�([��M����Qmmm��bWlٲE���/��LW��S�6}o$�����L��۔�) �Ý���i������p�:֬T�w4ys��49}>œH(�`C��6�S��N���W��I{�~Q��K��V�����RE�}�zZ��=��\�_4Z	c����*Ծ�Ϗ{�s�*Թa������\m��]�^�KjkU,�G�ț��`]�:ׯ��1$M�[�����x��C�����-�I� |6�oѝ��xa�;V~�p �� N�WI{�+Of��[Զ|i�݇8���t���յi���  n|���ۭB��) �/��{ｧ�;Nk׮�1�C�   �C�1h9\���+аE��o�R�?C=:C�լ��O-�xo��o�rss��~WW������HHH���,�i�M��`0��6577[a~�qx7N������zKK6֫-�@��}e{��zt��n�|9c ���r����Q������De����9��N�_c���v��[��YmK�W�CV�?(
E�ܩi��_+k�I�`�m�U��G����R��C��+���ߨ�����H0���n�����`�<m?�}�2g��pe���Z��o��ݷ5�L8t�=����n���o�Qєv���*a��m_�\�F�x�Z��WT��W0B���E)�g�~z�ռ��>�������N�;J?�(œPk���z�*�՚�4�rz�������ͭ�俵���?�����h�eWk���B�[��Rk��:f�  ��;�#����v ��X�d��>�h+�nί���L    �wn��YEr������4������+�n{Z��5%���O���Wvv�����촶�L�	�'%%Y�yAn.�����
����	��fd7��=h�3�}����ު-��R����۫D銍���oғ��� �T��	'f��sf��[��q�<�N�O�z����k.�Z���{�&����6��L��W4J+.9+�m�gZ������0�q�G#.�J�����;������8r��3��G�������"ś��_����dM��3y������7}r���	���jZ�Ҁ�'+[S��rhf�D��N�������럨ᅧ ��RR5���_T��?�~@���4�?���f�s߸�ҳ���[�����H^��ד�|RK�9�
� ����L�<Y�V��J� v�9W�r�J��^Z�x�=�P�   @����+���ərz�]�N�`��Wɓ��z�U]�zo��Jk]�	����$���پ)�zn���qfyN�������Z_�z���f\3�=Zˁvww[�sf�zi������ܖ�Y�t�U�
�0�H%��G��v�a�\�D9���O�:n�vr�:op��?%q�d���g���K���Q٧	�on����R�EW����+��������}�jx�Y�/|J�9����Y����<���Ғ�R��]�ě����OQ�?��<�Y*����oe~�~y��|�����:`�Q��G%��i��њp��jz�%���������w�Ej|�e5��p@nߛ_�Q��`��w�|�7�>$j��>-e���۷2�yJ~�[}x��  ��	"�s^�=Qz� :�}�]+�^^^�9s�h���   ?�c�0w�$j7���I��ӟ��)�*�c�<إ�+ޔ��WT�iѤ�"M�2�
��*<7[k��7.��
��K��n>�Y���n��݄���@ڼy�>X�L[]���?�x�f�S<���7ջj�+a�$9\�����O:]�[� �9�S�4�O�iٹ'�c���_Ωg�sv��a>�s'�9δ�p߉��dcx���:?��d�(c�,�=���	-F#��=�4��>{�	�g3[�d@����O8E��~�LM��?���/�u�;���:o��YǟbM��,�EJ=�5���b!���}�I=� �F�{M}  &�v������io 쎍7���QVa[qq1-�   @!��!��tɗW"WK�[��5�9<~�L�)�n���6W�Փ�Uv�\��;J%%%V{0u�cԬ�i���Z�b�6�u�*��p�T%M����D�)�EBAu׬�?|�/�! ��W4J��`�9��S4�������R�g�[M�̄���5�
�FxB��=��� ��0�Tر�k��p�V	%���I�2U���P˿���$�N�7n܄;�2l�Wb͓�����M+�|���\$ �m [Ɣ�<�q1���1p `�0Aĉ'jժUVs{JJ�_+ SX�t�Rq����c�B�   ��1$�Ss�LHQw���;4$8��Z��ȕ��Z�e����Pi�j�y�5:/ÚY^XX����x��ޮu��ic�fUw{U�LE�'(ḁr핡$N��6���) �*��.�-�9��M�*���U��=����D7nwx<1	�;|>[�6�7�sNՈˮ��1����
.�b��N�J]		v���ˊD�b�3!Q�t���s�:V-������vz�=n�}c_�>�p�  @lkk�������` �{L����Wuu�N8�͟?_    �wYN�_	h�P��JC�ˣ�Q�Z�QۻU������x�}�E����T^�S�����UNN��fK���Җ-[T]߬�P��]�Nʗ/�`���g���@������%ɝ�! 0Z���R�;P�l-�%�vp�ЖX:Q%?�]�C��-V��<fv�}�hu�m�PfB�m�����Q<0!�	�W�2S!&nq��݁�   &����d}��6�{ ī��z���k�ȑ��鱊�***    ��chs8��!WB���	h(s�d+y���z��-ܣe�e
�ڠ��V�lU��K)��R�!%�JNN����Tk)O�qBB���`0h5�wvvZ���fkki�P{�C��ڕ�vg�z���(�g��rO̶����6��6��M�&^ @�_�Q޹ɝ�	��Rq�-�>��A��8~�|�#�]�E��0��x�$����o���o)n�>g͟w�6�����o�Q�t�ⅿh�F\y��~�3�?fbLŽ�  `(1�/JKK�z�j�|>���� �3|��p7m�3f���?.    �G�Â˟"���
6V(�R�a��/g��m�����`�z���lV��U�-m�7*Խ��{]r�t��vY�<���zzz��ӗ�`�����˗"Wr��T��͒���0�Y 4Y�W$Rw�%N j����K4��{���uk���/kܯ�4�C���%ܱk�N���f�G�U,��X���\��d&�x�{�����Q��ECY�?��������xQp�����4[�$�ݭ5�����6  `(�w�}�����25���t ���-[�Y�f����Z%��;   �c�p8]�fɝ���M
:�ޟ��'OF���Eʮs%���� �j~����*8��L�!Wb�nߖ7/_��\E��R�����sJ�{9��tO(/���0ov��]1��k�q��b��H0��͛T��GT�����R�s%%+��sz��u[��[���-�~1q�^r�m�p'�X�$�jkU$�>v8r�����8�^���+����`��}i8�=�;�D��S�w��p�dA  ��f����
�w @0+��_��Z!ĬbV<omm   ��"��a��K�Z��-�V�{$��(1�9\ny3Fȝ�- ��`]��n���N�W���_���4�n�����=��K'�9���
�+���*���t�pg�����=���+��q} \p���z�"���:3I�l;3��%���y;^x��?�`��f�N�^Ӕw�Eʞs���1���A��Jر�;nҖ[~'   �>31wڴi��������o��� �˗/���}���ӫ��*    �E�Ó�!OZ�\��
ԗ)��l�?OJ�<#��;  ���Q*�ͭ�ڷ��ilЇ���5+5��F)c�l5��{L�t˿߶���^ָ��h�o������    ��c����X�E�� �ӊ+t�'���Jx w    ��İ������PG���r�\�$y����   �r�4��{�NM�}�H0��_�p؇۷*��2�������4a�
.����ܹ���?��   `�L�>]---��� ����K�ׯ׸q���t*   @�pz�Ӕ���`k�����Cv���7s���Y  �Uc�K%M��K�����u�;�GR�?H�{��{��7(��3����s���S��WZ�    0L����M			�z� �?-_�\���Z�f�JJJ�K    �C����'5W����V/���%OZ���~"  �]Up�e�9��]�N�ӏ��{�O�?�R���*aυ�:Uq�-�M{���s/R�=�*PS%    �OIII*..��u��(� ���+W��OԦM�4m�4�   @�p>Ŵp�rF[a�`S�z������=���  ��H�g����w�:kVj�w�&l/��ST���)PU)칪�Q��Wț���X��^p�����    �Ӿ������t ��:;;UVV�Q�FiƌZ�`�    �w`'���r���ݮ@c�B�-lw%e�k��n�A  �ϓ���7�%���d�P{�V_s���n��ϹPe7�R�s��nU�{�F�����oQ��N    �_�O����V�|>y��/ �W�֘1c��x�ǜ��n   ��@��$��K�n��ѽ�Y�������  �'L{��w�j��&Ѻo]��u�oy�pW���[c�ξ@[n���:]�~�^^|����D\t��~�S   @�2e���ꔕ�%  ʪU�4k�,�_�^�'O֒%K    6�6���/o��]��i�&�>��`�;%[��|� @���+u��v�:�wެ���pԽe���J=�;#S9'�U������~�-�߬�]��{oU��^    ��233����H$��� 0P�	U.�K��w    �����O�6o�[�����)	C���;9K��|9\  ����P���w�:�o����A�Y��w�
�_��G�j��c�U?�g^�Ey�
�k��_x��~�   ��2����r:�JJJ  ɴ��CƎ+    �C��M�Oެ"y���R�`k�"�a�s��nݩ��d���   �S��)*��ov�:��J������!g�/=�������sl�z��^Y�s�Zܿ�[��ϿT�ݮ��   ���4i���ڔ��l�� H�W�֡����.y<�A   �>��r���dZ-�=mV�{��]\�\	ir���^�
 ��ȝ��@eE������[�S�4��{��'ؾN�'��_�B��zw&�_��}��l�/��2����o���_����JLR���j�M����<���A  JKK���-  ږ-[��ݭ͛7k������    �����;%��N���Z��Hxx�l�;�ۻ���py �P�s�Y*��ƨ�7k�iB/�S���U��Q�t�?��Z�[,|��T��ɕ�����ÎVBI�:׭��iq/���ݟ�_p�e�4-�-�0|�|��~��z�X:Q��'	  n>�O���*//Wj*�4 ��
��i�&��~M�<��;   #܁��&țU,o�H��7~����&���)WR���Yr�S� �`	t[�S����ؼ3?��;n��aE�iqΞs�������|���o(����t�ڿ?����	�joS�����}�}�gƭ��uB��y�/q�U���hqON�~����z�����\�y�_Z�hʝ;��؞� ��4a��E���Z  Ѱ~�zk���   ���@2���Y��	Xa��ٺۅ�r8r�Sz�r'eX�  �nox�Y[!r��b�t���\�h��=.WR���uO=��*y�q�Wv�:�W�މ���T��K�p��kV.(���il�\8P��7k��~nk|���[�/Z܁����'��b;�$�hܝ^�rN:���`]�Z�K   >M�8Q�� �jݺu��e��c]F"   �.�@�8�^y���
�w4}v��}�X�v_�\IV���� �����m���9/������	�T���49<�������[�0�.Q��S�^��25��2����X�߯���W���G�#Ոˮ��➒���-��N �����s�j%���X����+P��Rѐ9�$�32m��yt�"=A ��4i�$uvv*77W  DKmm�ZZZTYY���B���   @tpb�
���Z[$ح��f�;[�lU$v���+!��-1]��   �U�^SW�F��G�96����R��~��+q�$��܎�E�T��BCQ��_Tb�D�W�D������N7;Wu����F���Uq�-�Ͻ	0�����?h��ik|�EW��w��A&>�?�s�y��s��*��FEC��y��>��<��  @|r:�***Ruu���� @4�_�^YYY*--%�   � w ��<�\)�w���F�PG�B�-
���f��{�hO�>���  V"�>�7��7�j�ĳO���{o���;�^{�Q���n��ϻd��c��_Z(|���P��eJ��W�c���ʚ}��|T���l�W�W8�ϱ��4�{-��T��C*��[��Ž}��;��*��&)<��̈́���5���יP @3������E�  �6mڤ�S����D���    Dw �8���ǍHO�
����>�tj��hw����X���  �<��F^�u9l��͛{�*��
��ϧ�ΰ56XW��E/i(���	V��.��|�{��r�J~n���+��#ӆ_~����l�/��JU����xM%=M�֤���'�9�7�Xi��7�1�u���5��;  ��1cƨ����v @L���Y�����	   @�p���;9S2�L�{Ha+�ޮP�G��H�GC���g��%�wK����L   ���T�k/)����0v�R�=@��-��ɚu��i���<:_������3���]Y���^���.$�S��c*������slҔ�J�>C��-�j�eW�7��ϱ���~���O �s_`'�n��Ł�;\ne�r���&����  �k��������� @4��׫��U===V�=<�+�   �$�� b��]�i�����"��t:�{٩H�K�ld�������M��w���D��4  ����܍���4��;�<{{���<���"�ǣ���5�LZ\s���il��~�~k�;
.���{?2S�������/WU��K����7_Uw��
G�96����R��~@�%������[���
ww  �/l7����D �7oVQQ�F�i5�������	���͂�<s����ӥ����}~t�J�	 �������3�Vs�(9�e}䌄u�����[��Kr�.�\	fK��#Ez
���?��翗��P�R�V7��fs�}rx|����  �Ɨ_P��J���>�f�6����ii�����.Q��3l�m~�uu�m�P�4yo9�~[c+�|�Z����ߧ�ˮ����sl�1��_4J]�7	����q�Wl[���*퀃���0��ý����d#3�+�������9�ܳ쯜b& ��VPP�@  ��� ��0���kU��]�-�B���?]���&oxU��9�`hz��T㳷Z����S��HHc�V
�p�"��
��z7�Sv8Ĵ�F�=�u�>��5��kVP�4�G>jX4㬛w�>�/g��������n>7��shwy>�>~  0 �cy��h��W�9���N8U���ߏôÛ�#v�,x@CU�>��g~o���)�`}��yB9����X�˥��_��7�P��`P��Ac�k[�3�=��;0���_�ֺ��K���Ty���{��[P�����5�u�;�X�J   ~%%%Y��ͩL @�P{(�Z�   D�
��G��޻ �  �R��_5ⲫl�M��5�Գl��ijTË�j�2M�v�/�@��Ja�U�{�Gw6��s�:O�o��B�-B�0��#�x�|#��y�lm����=�
 ���X��*���}�M;N)������1�9�V�ިyd�N� `�0M�]]]JNN  �RYY����   � �  �AǛ���C��oD�<��r�c�R�9;L�q�tmޤ�w����slҔ�J���ڗ/��gΜ%OV����O<�pw��*WJ��q��?�L�����]I��=�lZ��Q�'���ޭQ��~�c}�#��/Tw%��bxI�k���:�_o3�ؠ`m��8k5�p7�$�~�;��9�[CC��I ��6f�uvv*77W  �J8VUU�F��Wf   ��p  ���<u_�;J�q����x�����L��N���=s�6���~۷iǶ��P�N˰5.P_'�9X��w_p�e�z�EB!��>�F}�Vȴ/��pǰ�1s���n|�m��w�\�Z�����z���ȓ�w-��S���WOKs��;㈙�V�0�|��� ��VTT�P�k��� K�����V   �  ��N_�m���˃*ؾ�iU��������L�Դ>��t�6��G
wu��~M�,��m�m]�:֮�P油lm���]hxi���6�_<�ϱ����8�sjx�Y��kն�?�D��$N��Ɨ����JLR��S�5�DU�{��~��L���zT��*��K}�u���:�TU?��~�w��]�`��  񯠠�
:��@ �����R�����5k�   @tp  @|s:5���)���5umZ���Q�g��KuO>��y�9֕����'�����x��s���r�;�eM�F��?��\�_���o�����/'����?�p���@�s��*���J7^�������y|/����&$��>o菀�i��8�[c;V-�&�  ��fB�999�� qak�{qq1w    ��   ���7m�ݨ��������
�&`��wl�9�l[cC��I�����*���č��p����GmK��GW���*ܩ}�~ 쾌��Ӹ���_�B�DwU�uj}o�R���slҔ�J���ڗ/ݣ}�~�n�����  ����V��4� k���
���   ��!�  ��e�O#.���`C�*�|GL�mJ�?����ń�L�k��ջ����g�W0��غ'�B�@��Y!�����5>�%Z{�ཏ�7=m-�ƹ�	��L�}�%�<�P��]��A[w#��y����wgG�m�kk��n  @����SW�c�	� k�HD�����gUB    ��   n_s�\�"���^���0k#�n�q�6����W�Y��[��J�_�R���Z�
�%���T��_(P])�9�?�ָpw� ������y�
vGS����o�X�Դ>��t�6��G��ع[�J;�0����;������f �����k�ip �pw�s   �`E�   qɝ���C�Ԡk�Ͽ��E/��0�zL���9m�NsO;G����]ޏ';W�G̴5�4˷-�����]�Y�/-T�q'�9���(�����_	{�W8�ָ��&x޼ey��>���@}�3O(���JIU��T��û�����0�n�  ,rrr�t:�1q �h���U8   ��!�  ���~ȑ���i]{�Uj|�X�B�-��I�zV�c��ʘ9���r�������h���i+�n� f�7E��x(J�w[�z� :2��\��F͂m܍���v+�n=w9�x[c�6�S˻�  ���L%$�[!
 �h����VIIIQkk�    <�   �)�9�L��F)�֪�7��/wY���a�	8^�F��������Ԩxa�J�܍ܹ�v=��p(��sl5�'F��q��f�ȿ�-��N��J-���Z) y�i}��df)��3T�;{¬䐼���ƶ��P ��?�$&�5���˗*i��}�M�>C	�ƫs��]�G�ig����[�p�}|$"  08ddd��� �xa����*,,ԪU�   `�p  �v.���p��O<�_O�� ��{�%g[M�ɓ�ek\��U��)B�m
�T�s�:�}�"���M˿�V�5J()�s�i���VW�F۷�v���u��V�=��ȫ���_�v�V=�~�Ap7��z����&[c.��j&����O8���_��KM��S�団�_OF�5��/ެ�Jͣ�5�F���=�\m��G�t��:vD�A��}�� @�p ě��577+77��;   %�  ���W}m�p�V��t����G+��9p��T���7T���;g��G}��}t8����7���m��=��q,�!{ \t������IuO?�Q_���,ޗ�q�v�j~�Ua7��w�{�����:um�(`����Θ�7i�T[w�ǣX��ǂ��ߓӟ����������B�@��m��w�u�mG�?���{  ���t:��������C  Muuu=z�    Dw   |�+9E��3ǘ�n��n��j�xX��~Kw�!7ӆ��O���F�N�P�1�m�i�oyw�пܩi*��u��Lco��?���o�oZ�	�#�U[c^|��|`��������s�}���S̜��瞴u�yg���G�` �`b����+  �	��?^    ���;   >!y�r�X:m�!�	�Z���Be}��>�z�
�~�L5��B�cM۪��	�� �: R8X��$aǪ�ߧ�EN��ϱG�TBI�:׭v��/}�����O	��Q��A[w#w�<[wWJ��f�d�6�j~�5 ��#??_�HD�C  ē����Dl   �h��7   >���no\z�0x������af��g�k��L�v����;3Kع`C��z��ߪá���?�^�/�㬉Qv��i��o
����οԵi�����96��#�U���6~渜�N�ӟ`k�Տ��֪4   ~���n �%pw�\   �  �I�D��^Eݕ����sl�Q�ʛ��@M�NǤL���q��c5��E�/X[#|���nW���غo�9�l����45
�����l����NEB=0�D"�y�!��}���9�,m��W�9,��y�����	  .��ɴ� �	��{_k   ��!   ��z�![aT��m���i�c������y�a`���-��Z�JNv�c�J5����:�ϱ�8��z��o��1s�������P{��p_ G5��?���9ܞ>ǚ7���;m]O�2UI������E/Y��  �����(����  D[cc�B��W�J#�HD    w   `�0��W^#��eT���]����JIU��l�3PY��-�	�o�����
;g���܍�y�����	
���P�U_�=����jm��'XW��W���cf�9֛W���g��v�}��Į&�  0(�����  �Ƅ�M��<V���   ��"�   V���ה~�Q}���,VڌC���׶�^��gXM�v�P��ZX�?*�r���>�K_����j|�yunX��1%}�5�ʬY'���ǅ�˜9�v�r��C���* �W͂m܍ܹ�vpw&$*{�i�n�
տ�  �����@�;  n���)55��;  ���w�mUw�ǿ�-�W�I�
��M�+��g � �2
<--�I-��lV�%J�R��d��{ٲ����B��H�$ޯ�}ٖ�9���^����b��;   0���Y8w��ة���srx;����B����&�<��
�=HiUa��<�+0��B!5=xoؕ��8����8�>��I��6�:_}ɚh�V9�5�p���VV!os�n/9�kBW8���  ��T�MKK  ��Tp/((PCC�    Dw   `i�9+h�**�m�j�`�oSs&ov��W_�@C��{�8�[}ʎ>ad��eر��˕��?d�쭶Q��;�����*��r��6���>�f�! #�Yͥ��GU}��C�u�����Tw�_�u�����Bj~�	v  $**� �Yww����    ��   #H��S���Ty��C�u�\*9�5�w�׷�.��?W@��{�����:����W�6����8�9����7���X�{P�3.���!ۖ>ߨ��fk5#s�f���a��7�Y�B   1��=) ��b�f�    �G�   a���Q��s���P�O��u��T�.9�Ȱ��kkQ�+/
�'��R崳���C):����j`��p��7�*��V���� �|j�����hȶ�������z�5�k�|$\��` @"���  ���322    ��   #L��e���}�n��m3�M�*���%����ܰ�����
�}��@�:�����<lȶ��U�<]������9��yI����������+�n�;�
�;��Tz�1a��wu���g  ���t��&����3����>33Si��~  �	��������QQ�e��k9�Z   $�   �df�܍��Z���N	o�PH͏?$ 5�WXw���S��֛�/h�z{o�f�! ����kl��ZX4d[s�YUT����
�����<  ����6�B9���S� �zzzl�	9�
���g3x   �;�   ������_�U���#��zζ?k�wߔg�
���w����ʙ�ݐm��G������̼4��z��� ������㪜v��m.�J?FE���-O<,  ����� @<���   �� �   �@��>�>��U�z(��,M���a��<o��x�8g�&����VM?G=�|�����Õ5i˰�z��p�]��1�Ȅp7�N?Oi�a�5�j��/  ���R
�g q,
���	   @�p   F(0'�n�UV����ݥ�����ڟ�Bi��C�M���&y�hN�jν8��To�!}K��ӏ����C�M��{\&� ��RSS	� �����    Dw   `�2�2S�4{�"6f�S�*���g!�OMݧQ]V{Wq�F2���43�.��{�}n�=� ���dd�Y\�}4�d�j�t:	� ������p���H��OH   @� �   �`-O<���&�������T=�"932��Y���To�� lH��'4��k������^ ��9k��>do|S��l  �3�Fx1���-     ��_"   `kyz�j/�����<V�'X��P ���X���o�!�_���ަ�gW�qS��W2�eM�"���z{#�ۑ�̹:��:�fU\��sRD�k�7W   ���Tp Ļ��>   �>�   ����T��Ϫ�У6y,�e�f��H���ppff)5� ����V%����Tٱ'�҅�w�@o��K�n_?���#���O���ig+s�z{Էt�Z����������k~������,T�g  $>*� ���   ���D   �gf�p�*�>���Z[�jW��Zu�5
b[%�h�)fm�!ۅ�>�:;����-V�[�)�=��*;�de��,��&��@�v$�q��A�'����)9���~Gk}��VȽq�,�|&����{�y8k¤M��  �CZZ�  �w   }�p����<M�RF�|� O�@�ҽ�6�3����~]�5+�Q;v��h���nΣ�4а.�v�5��<m���U��ZX��K~V[oc�*Y�P6���=N���:����P��[@�(:��o���/gz�ʎ>�ں��
������OVJt͏?�1W^����j}�q ��@� ��^� Ŀc?�C�?�dU�� $�����SR��XWܞM
�;CA��s�����   �(R��������!��+|[�G�ݶ���+��a�=Q�g���7ߣ�����w���Y�_T��e�7A��	�ovíV��p��:�ގ�S~ⴰ���pk�6ԫ��j�7G��vah-O>����rnd���_�X+H  ���r� @�#�$�,_�� O���Z��&�  ��2ƌW��S����h���qr&oV��UքIC�s��*��z�r��N��Tn��Y���U�)Q4?��F]�S9R�D�[�0�k��~���-MJ+-�������*;�Tu���L��@ �����<_l���s�� aǋ�+��Bj�{�����Ji�U*=�X+����������a�Sy�Y����_�*(T���*{��mO���+�K�$���[��c�6k/��jοL��1x.��5:+��
��j��$����u�xʏ7��<&� �L� A �_k   ɂ�;  �0(?����:9Rc�Ɲ	]�-٤W���xSq�t���w���wJ��fu���
�9�vߦG��eB�M�<�Q�4�>fJ8Qb�T#�x�%���Ҩ��Pj~��]��kܵ�˙���6�	�6Ι% ل�����LOW���*����A3�nc�U�����  �#%I� $��'��!    �E�   ��w��
'����á�Z���{nU"03�����Z�y\X��{nSŉ��*)S"Z��?(8��z������:c��Y���Մ��%���n����HJ��+�^Y�D7P�V����ʳf�2j����4��Ŭ�  �G0  �n``@(>   `��  �ب*��#��y7=�@B@;^yQ��F��U�ݧ�_����)�_�ϭ��ܨq��A�ƽ����1��s�Q�i3�H�ߗɣ��:���˖�q��Q�S�*�=��:_{Yq/R����3]~��_�O��k  #w @"0�	�   ����  $!�˥�mwFgf��v�I�}I�΄�L��z�Ea�i�7Wذ���S�wVɡG)Q������&]��b�~������>\�(��FY�m�x�x���
�}��Y��p�U|�aJTw��_z^����Q3�R9RR�jo���I   ���~ ���    Dw  �r��+Y���|�Õ�_�Da��g_(9C���Y�����
i�U�(c��l��❙��'gɳjy���B�P������wWq��F0�W�THV�ܴ��s�s�tU�w�\E�J4�w�"g����A]o�W{�V��y
  $� �D�t�B/   �  b�T�����U\�D�Y�Z��n��g�ju����w�}ȶM�>`��14S�zѹ�h���(w���}n-��u��Z���km����A�������c�L�N����)�A-�ťj��c��������jz�~�{�*�����D���S��{�IӼ9a�͊�o�"  �|� AJ���   �4�  b�u���<m��y�@�Z�~��ɺ��0d���ަ����g�g_L?V㮽^eǜ�xc�f�f�"c��r�[��������19S�}�nQ��6�˽�3eo9y؎��Ѯ�W\���^0��^�=�����8*����)Gș��x�Y�R�9Ś\�H�_z�Z"{��7�nݭ7Z�m  @�	r� $��Tb6   @,��   �L(�T�5Z������������J�l"�~�m�=���9b�B!���jz{{B>��_u�:_���\q��*���������Қ'g�0@H�o��&����mҷd��{0&����?4��_*��B�f���-�{\�������SZ������J�@<���#-��B���*;v��O:M�Պ]o��%�̐��S	g�\c�_l9�9\��61+m�<��  @r��;  8�N   �>�   1fG_�r�&\��!�dǛ��gU7^����mnԊk�H�J�K���
�v��p|}{��o��[�y\�x&D���s���d��<8��cz��o�K�R���˳z��Sۿ�k�o~��W\��(�����ɱ��\��{U{��o��GK~r����/J�ˏ�������O����^� �/�*GݝS��[T���*=��cJnްO߲��$Js}1���@i���g�}뾮�_ג�δ&f ��D� ��   �A�  `x���c�5iKeo���i��nO���}K������?/��ܨDcB�&8���k1�F��4����Uw�-��i7�JJ5P�N�/�K��faәﱩBk6gf��~����ʭ���9��"�?g����ʽ�3��X�xbB��/=��)G(s�X=u���u.�u�����^]c�_�G�)��Ĉ���R�A�+s�D932"6�9g�P�9��~����,J�(�X3秎��dmfu��-�R��-�*-WJNnT���&��|����#Y��yU���ʰ�������  �[0  ���0    ���;  �0�[����]]o�jm^���F��/a��G���A��>܇!G�V\}��	��>��b&��~���a�ܽj��c  #K(�W� ����L�   b��;         �a��� @�KOOW�    Dw          ê��G��J� ��F�   ��         �����Դ���������  ޥټ�9N�}6�?%EL  @2!�         � )iiJM��ۄ)�)�ڛj�>�/�� ��p:��:8����=.    ��"          ������v+??_  �+'Ar    &�         V�z;w @�s8   }�         �`0h� �W�z��^   �>�         �2����/�4��X[o�Ooo�  �W�z�����{�?�fE[��M   @2!�         � ��޴���ü�Sa�OOO�  �W&����o�ӀW�    {�         v}}}  ^eff���   @�p         0�lW�  �L�P($    �G�         �����  �;   ;�         ���f9 ������`0(    �G�         ��kjj"� �[yyy���   ��#�         `ص�����)%%E  ě��l�   @�p         0�<�:::TRR"  �IZZ��N�    �w          Î�;  ^���f�    �A� 0�z�sՑ]*     �DV�۬,o�  ������S  �pw��   � ����{j�N3     ���|���e�� l� �x���e�4    6�         ����  ޘ
��`P    b��;         �����(��I� Wrss���'    �A�         @\������  ��\�����v�    6�         �������WZZ�  ������"    b��;         ��000���&�5J  ă��\�|>   ��          ���Q[[w @�0w��-    �C�         @\0r�p8
� �p��;   {�         čU�Vp č��<���
   @�p         7�/_.  ���Rvv����    v�         ����jooWAA�  N���֪"    b��;         ���v����B� 0�L����	   @lp         7L��Tp7sC��  .f�Uoo�    �V\��.eM�B�[l���1J�͓33KA��]]�6�ɽh��>S��O�,%'W��쭶UJV�<kV����o�b%�Լ|�ǰ��_>�uk����?�/���O����Z�$�/�W�g˾�6�\�S~���c�H���L�|m��6��7���
        ��f���� ��Tp��K�
  ���[Ζ�(s��J�/PJv�(��]}���Uz������#챷\E%�wv�������K�E��ө���|{�UX,W���{K���P�?,����*��FϚ�j�7wX����P�#���nr�ʑ�(��З���6+��9�;�mi��^������T~��*�1'ߡ=u�����xd���߃߳���V���k���2��[��G]�S5͛�U����^��Y���h�/o�ܿ�<����i�5�+80��:�(��Fs"�u�݄��\�[U�8ͺ '�Q��9!7Ι��{oO��5        ē+V��tZaw  �Czz�������#  b���O������	��crb��>��G�X��d�VV��7ݡ�v����ϑ{��Zr�yV�P<˨���S�[N����1����V��%1?��&���4�t����s��&�x��**��B!u������;�~�a�v3,w��:�g�R�>��gf/p�����Vχ�*�w�&����W�v:�
�i�UZ|�iq[Q���5�w7Y���c��#����L�f�2l3�E�?�	��J;Z��UT�Q]���i���d���_       ��3��n�. `8Z�l �gZ��ϻD���PJV���9�����i�m7�aάĩl�&�����*ٯO�[k������S�Y�Z�(��F[?��w
%k�$m=���C�Y�\H>�R���Γ3Y��aVT�y�������G���+�R�;���#��ث��r��M`N�[=����z�uBN䓱Yj`��_��L����g����o��+�X����\ϭBr)���
�����]s��P�C�        �˄�4f� 0������ @,d����n�Cٛo�I�i���½��+.���Y�����p�W�c�p�-���í���f�o��������h���`������L.x��7'O����0v��Zt���w�Gt��ܫN?O���&b���/�f�,��e	r��zz؁��3f�ၻ��$V~�)V��pT�q��g�.��L*���df�7���B~߰,Q       �Hb�k׮ոq㨜 &����'  ��T!��G��v��ﶧ������v��MJDY�mn�Ñ���������;�'�&�,�
��)�����~�M!y�ﾧ2F�S2��agmy���|�
z�#6n���x$���Tv�I
�{����T"���Ga�M��Tƨ��Y�x���]�n�*)S����_�TH�r���Fr��^�	        ����hŊ�{� @����(//O�푭B	 ��ert[���R��#>�	�n9�1�*x��[�&�=l�7��x���~��j��n�ҒL�6##W���6�����#6fL���1���r�����#��B���m�/.����PKh�_i����{�p�gȑ��H`����I��U�        D��ŋ @���t��� �hqffi���D%�������'g)ѸJ��*�ec�v���cF�K���HQz�qjy�Qu��ZDƋz�ݙ���n�]W�ïc��N�o�"Gb͠u����0�"*�8�6CJ�@�e%�=J���H`f7��8M�sf	        DGGG�UQQ!  b��C��� -�/�JY&E}?���ÎN���v3����U�;&�9L�=ok�F���~�ώ=("cE=e\}�J��X03�F]p�V��g[f�M��h�(;�d�        DQww����TYYI� S%%%���  ђ9a��O:-f���_����B� b���W5��l���&n��%7y���]%e�:�|�R�����;�Y�R b���[T���q��@4do��ҫj4P�N         �z{{�z�j��N
  RRR�
�  Z�\q�)Q�O����JU�r���;��՗U��)
�> ��Ug�'gF�bɜ��ϹH˯�D b����/ש�ҫ4R�Lގ�;        Q�p�B9 +���r:���|  ���F?�'���>�|5=8[�>� �β�_���WzM�F����Fd���S�T~�4��#�պ�n���5;uw�,oc�j/���J˕��*         z�����ޮ��< %%%
�B� @4���ri&�Lg�	����� v|������5��ߪ�#%�S��U\�q�p�:c�R��m�z����V8=��B��d{G�K�3.Ԋ�/�1��yC��+�n�9v��v�5��w�Z����c2'���\Ż�<��g�V�vT�qJ�/P�(;�eԎ	����X         z����z�jm��VEw  ����T� Q���d��F�����~�.��w�S�����̙jzh��� ��ש�����ޑ���cN��������5��9��W�[+��;ڵ��3��k����J-(T��;^���v�����*�p73}*��n�_߲�Zt�)�[��m&ɿ�]Z'v;ʎ:Ѫ��m�`W��YA�p������������]�L��������֖H�w��V�=�gR       0�zzz�|�rm���� Q������\uvv
 �h�9�2��ۃZv��j����os�������B�v�J�T~�)jx�nv�-^`+���̲p���fk"G�j/�yBܿ�kkQ��H�w��V����
Q	�WM?�v��@O��y��Mߺ��0�7M�?����.�˥�.����L          ���ӂ� b�������z @�eo����=�v�����o�ۍP ����ZY�P����������
r��"pO�/P��3l�[��?}'��s{�=�}9{Ɇ�cOV����Q          Oss�֭[���j�B! -���ֵ��U �h��y����=���'���W��W*�m/��{̴�J�s���- �W�W�6C)9����*�M�<��6���Pũg)5/?�q���:s�V]w� ;��(        @|����ҥK5j�( N�S%%%���'3  ���	�T��!�����Ff�����.R��T�����f�Ej~l�B>�0r��,����<U�r��~�wߪ���m=�j�3K53/�5v������-M����׾�K�&�����c        �G���Z�l���� ��1����Tuww �H�9�2[U��������n������WŽ�J�G��ys��+�������@_���63�OD�z��
놿�]M��V�S���3mWq��~�V��ka�23�
�90���*��/_��I[��޳r�         ]0��]]]���  �P^^n}�Q� a��7S�A������*�ݷl��^|V���G������#
���Է�^N2>s�K�'W�0"pO��U崳m����V¬Lmf4=x��Ͻ��>*N���Y����&�L��<��.k�Z�ۯk��N���T|�a��_�D��        �:::�b�
m��6V� �H+++�V
�: �����گ޾�3u��Űۯ��*��[��5Z%����F&�14!���[�680��g�T��|���Z�*.�q(���C��e�z{g��m�O���[U�M�>\��,������F&S����{�ߝ1�-V��*ţ�W^T��ϩh�)l|�����k�        @"0wS�}��'x ����|eff���[  DR��q*>�Ƕ����F[�/SŽ���Tt����S3��x,U�G��߱������=O��ǉ����66(��������f�mȶM�> ��υ���{JV�*N=�v���w(�����թƹ�������W1���s��#Ӫ?\kMv(;���o&\,��L�b��]q�&��.��z��|Zq��z�U        $���>-Z��p;  *�����^�W  D�	�;RRl����/��������7�^�ڱ*��c��B���{KK:S������m
��~֭�W��|Ҫ�>��k�����Z��_�#"wS�UTl�O��[M޻Q����{vN�}L�wSe~���$�L!�O˯23�W��*{�v��^�������M��T�_x�)*��8i�r�yBb&�t��%���/֒!         ɦ��I�W�Vmm-Aw @DUVV*
���	 �Hɨ��Î��o��7H�o�"+_��[�jλD��>�Q�Drh{����}UN;[���
�{�����VA��O?R�k��.u���U<��G�X����tϧ�q�=V�Ϊ~�p7�+O�a��	���6j��ҶU�}�E����4���_$���_���5x�my�Qk3����`��G         ɬ��],�رc	� "���@YYY�j!  D�	�;R�E4��/Uۿ���}����*��`���O���T|�aV�#���^���+�V�r/�LK~r���)���S(�&�+N�n���ÄqM�|S��s�*��a��{n��g�m7	H��K�        ����V�}�{� �S���x<  RҫjTr�Ѷ�����M���^���U�M�݆��/Sۿ�S�I�\e�ۤ��3=]��ϱݯၻ7���U���٪>�[���p}��+          ��Tmojj�ʕ+5f��� "⫀���  �bUoOu���Y�Bm�ozu����٪�5a��o߄�� I�p/?�t�����cJ�7>p�"�~�-Vy;U�S�T1�t��y�          $���}��?~<w �&+,,TVV�
� @$�WV����m�[w�M
�������ʿU�ρ���̼T�/>'qM6:�n��W�~��~̒��M�`��7=t���:�V��3f�q�=
��          1���iѢE:�� ������>���G  �S}�O�p٬޾f�Z�?�cX{�*�� [Uܳ��Z�{�o��`�mt����iJ+���'��W�}w(��fݢrS�=+;�>������{�          $�߯��F�X�Bcǎ��; `�9�NUVVZ�{�^ 	i�U*=�D���n��BĎê������0��˭~Tq0�6*��LKSՙ3m�k|h�|m��$G���Ϫ�nG�Y3��1�{          ����U���&L�@� ����ʔ������� "����|�ujy���ڿ]oUd�U�}�mT��>�|�e�pڨ�{�qS�V^i�Op�Aý����������O�U��U\��������         ���ڴh�"9B� ��RSSc}t��  �J�Uv�I������|���U��՗U��~���\pw ��v�ݑ�Rՙ���Q�#���ܨh����_u�y��U͸PM��(��         @�3����f-_�ܪ�n� ���eUp7�^�  ��Gtfd���m�W�+Z���*�s_[U�s��A���H]o�& .��eǞ���[}��/�gݪh���VU�4}��vk���'����         �Z[[��'�hҤI� ����N�S���@  �*)S�q���Ww�ߢR��+�/>U�k�Q�	��0���	�V��z{�Y���7ϛ+oS����֢���W��sl��>�"5_4/          "�ܗ,Y"�ۭ��t�A ���Z�c__�  ����]���I�OD�z�W���*��>����`'����{[ 0l�ˎ>A�5��v��T?��B�ݷ���i���WV�����        ��HIQJvN����
�˙�f��M���h�������J� ���"���Z�۽<w��S�9�6��g��"��u�+��He�ۯ�^��
z<�6�����`�}l��9�R-x�x�p;�n��W�}���F����f5=�*O�a�_���#{2        F���1��7">�y���/j寮���m���=N�w�r��Q��.����jzhvD����sUs�O���������_���0�577룏>�n��&��a ��ѣ���z;� _I+)��~�q��z����Jy�7j������u7)o�]��U��U���E�8�O��Q^����~�����by֬�S}�J�ʶ���֢�y�+ʻ��?���ﶧrw�Y=�# W���8a�K;J�F�����Y�To���0��r�I�y|-O=*        �x`��(>�0+`�`������E��2[�&Z_��r����u�x��9��)?֘+�����]�Ф���g�OQ(�7�����ޮ��F�Z�J�F�R��9 ����TYYi}���/ �6gz�
�=H�K��I����l��Ŀ�R���Z_�ׇ���F�����c�^�Y��b͛�v�>9r_�|�Jj^��O:�v���o�I����|���U�w��V��/�"�����W`�}����a�+N9���-O?��ukKޖ&kfS�g��W9�l�         ��xZe�����eM���p�7�~L��%���۲��F��6S��E��T�mjj����3��; `H555r:��5��� b%w�_'MP��%��eԎ�:��M�u]��Ň���2�o����U���Vv�T�����jz�~ŚU��f��L��~wW,������_g{D�V��,[��冘�uw�]á�ΛU~�)���go9Yy?�Y��3�        ���i�OZi��o/�P��J˾g��&�p�B|��r�\
ڭ�	 1�5!����&J@,m���y�U��u߻��vLZN�*N�n�[�=�*��V��	]o����������b�Z���	���p��IUvԭ�Ⱦ�
��u��[�?!Ϫ���{�csmW�/;��         ��|����	�wy<�����O?�N;�D� ���˕��e}n� K��R!��︫�kjm��wv����.k��'{�A�G���FA�W F��s/VF�[}�/�Ⱦ�
��h?{�����/N�z|��ʙ�v��=��#%Ū>        0�����zU+~u� |���F}���e�]��T� ��رc�����L�3&����Zq�dҒP�^6s���Sw��Kχ��ה������wS����p����U3�R�]�j�0d�=k�͕VYek���_Q�����oS�Z�y\eǜv���"�l��u]扏�i�hr��5�       ������Q]mmmjhhК5kT]]-��/  �)77W�����n�[ `�;��R��U������?Aӣh��Ϻ�V��(�� ��0r�����W#��Nr�X9ꊓOW���l�mn�V-��!Ӝ�?����M��*4Ιe+�n��w �R��U��A*��`�l��\E%r��+��lJ        �%S����Y����=�X�� �eܸq�G3	���	 �M�����	�l�i����j���z��e�7!�>y��! ��LKS��3Tv�V��D��ϧ�?j"2֐��	mP�k/+�Y �U˕1f|�}� H��Tk�ɨ�.���L����,        0�����h�"uttXUzM�  #==�Z�àz;  R2���Um/>��
�����>�ⰻd�'��eU�}��E���9���J��_sfEl�!�Y�7�5`��o)��W��|�Upb.��P�n�Wy;�d�Y�F        `�������So����L�B� �1c���tZ�{���O� ���T?�^������Eǫ/�
�;R]�;A}K
@t9RR4��{*�n4ϛ����oȀ{z�([�|�x�^����
��I��і�SF�%+w�z?�P         >����O>��{�-��E� ���T+�n��P&� @$��U�Ч��S�o�R0(9�a�1�J�@�O9By?L��¾����#:����[��X�xҿr���fgF��� ������ݟ��v��՗��        񢽽]���������p h���֤'�� ����e�'�>���MJ���OJN� D_�!G(��-��B�;�#:��w�'%g�≿������\��F���5iK%3sB����        ��T孯�׻ﾫ]w�UN�SAS� 0"����q�Ͻ^��~�  ���J_gd���`��v�܁��;A�d��Q��D|�!�δt[�_ē����>��L�/g�mUz�1Jv-O>��e�       �({Җrfd*��ߤq̊��	���_cc�jkk���k����`5j��ӿ̼��� �I�͔��/w�&��HIU�I�}�t��ʍ�1F��l%�J FB!%oscT�2���+%+;��6�Ƃ����s�}5\>��סdַx�V���      �x7P�v����������ԣ�4~�A���0���7m&���Р7�xC�l�U�`�r8?~��y �*�@"h��2���8f�q��G�q4~�>(��b����u݆��M��\���k�"{�M������8E%���F�-��;����{m�]�%�'i�e��z���e��)�}/%3oS��<M&�       H }K�����3y���W~��M����>=����p������˭p#�F yL����,����n@�X�F]Ａ�]���}�ǟ�����NY��}K���O��gr�v�[��L�p���V�}� 6Nۿ�p��(L1���K��x��O��:��;xR*-{���)�dM��V{�g�r�춗.��U�'j�gDm9       ����\o�=w���9a���-٨q3ǎW����4o���d����z��75a����c����a��{"���`^׭/��5iK�l��F��**U���뽯��9�-����$œ�������N���g�P��3��?�x���V�>�B������9d�}`�j럔኷oh��;�jOE`�d�8O$3�~֭��-
 �C���ݪ@��ȭ�@��+G�B��B��t��H�#�%�+CΌ��-[�Y��[�u? $;s>����+��|y�����J���:ߗ�ϓ����Ε)�[f�Rs�ϡC�<��
�k|��e�+��ʠo`���疁�i`�#���\iΓ�s�\�r��|�	 H<��<��W^���zˎ9I��������S�jo�W��[m�?#`����iժUZ�r�ƌCw Ajkk�����c/| �����w�V��E߹Ϭ�����c�ʑ���M>Ƽ�Ćy֭���U\���j4�)��U�+�@�~->�6�c����Z��������+"<�;��˗�`�}�0g��J-(���C�͙��������,����[Fg�Dχ�����#�	 b-��N����7R�
w�}����N�R���*�PZa���d��ϕ���nV��,3�p39H>�;x�������[�gV�\y�J+��3-K �,���:���l����z�!��Ε>��=_�+vO�-���F�Y� $�@�[����ңN��}eG���7]g{e[��g鏏[�}��P��O�p���SGG�^y��~��Tq�￪�
�4@3 I��fk�瓪8����Wr�1��e��ϖ��e��'����=C��0��Xj�O������
�9�V��ǣ��� 6LH��S�I����㔵��q_��d�+���������-��4���U<�5=4[íh�C�a����-&�l��<{ol�sD�c*���Z�v�> Ě�2�m]����Vh32c��m���u��/Wz�8�f
 Q($�;�4вJ~wd&V�1�Nk�4.VJv�2J��UP>x�C ��̪�+�I@։.����6вR)�J/-Wq�5� ���b�p7�
�=�v�����|oѓ�ysċ�kת��H˗/׸q�� #��ޞ��eN�Togr�d������j]���'�5^�{+��f��5�.,�˗~��WG��%�zd\�Sr�T�����-]��J� b�L,���6k3��Ԝ���p�|�*-S�λ����^Sk{���OҚ��Sȷ���!���e{Њ���E����i��t�� D���I�/> ��`�@�J�����PЪ�i�ԜbeTN�X$ ���|\Ձ��g�z�$ɽ7lcj �@¦� !dC!��M�ͻ��f�Y�R @B�0���ӂ1.w[�����w�16.2hd�43���04��hd�ѽ3�yN:0�[v��~���Il�4a��fu�O��8�b�|��zs FS��Q���m��D�:�S�V�Mv��l
Aw H|72�jRB�D�!����C��:_}I��7*{��C�3��'p��o3��o���5REGG�mq��5m�4Z� �y�^͘1c�y�� �K��ׅ��^-��l\��5���`�!י�D��^8��}�����w������z��cOT��Y�ټA���g���h'W	�.Sp�ў�1+x���S��k���ᄶ7�E'�W��>u��˻�����S��)��SS�_|�j}�-����`��	m�_���   ��P{�zk�*���5��]�V�F���r�� �*�Ӯ��k����0MKq����iܦ�����	 RU,ԧ���l�5������o�߯�߿, �m.�O��|)��=jy�/�������;��{1a�I���C./:�eM�lC�a��ǟ<�uuw�~p��۷���X7n��GZ� s��:����Lr�ӊf ��ѿ%��i�m}���q���wۖa�>L�p��{��c
M�J���]��ۆmEH'h}���K������F�y�b�%_Jx���� ���kӷ�$�w����&�m��'�L��h}�I���	�q�W�Հ{�׾��6-}L   #�4���\�P[��~&`�lVN��J& RJ,�'4ٰM�Z}��`}�ƿ+P1]���(s�r����Y�Xt����{Խ�e���+g�B�<�z� p�����'T|����Q����)���ݪ�������"��[v�'��ڟ�~*���]�`&����RMWW����m��	�{<E"��� Hl7w��io0��YY*��ď�N��o~aXrtM-Ӥ��h����������Ѡ���ِ��b����t�0xfC嗿��6c>r�j������ćD��un«���
 ���]�r巴豿���D��ț�H�aP�4��{��]����d7��F����J+<��6����}�   ��6o��"#��~8�h�6�;�]�P.�G 0ڢ�>�lU��V��X_�&�F��%r�X���3�qf�������P�nu��ڱғ[, ����h֯n���Tߎ�Gt_���>�Ā�
��}�j~�s��%�k&0�}���k�˟Gd�d`(���UZZ����k�ܹ� ͚5K^��� R���<���T���Gt_������C*�ħ��L\����m��;r�l~ ���Af^��+���:�Ξ7�m\�*���Qiq7&|��	oW�mR4* �ӿ�Fm�/W��6f���0��{��j���k櫾��=5�#|�P���&�Mۊgջe�   �)�Vk��x�l٥H_�r�'��/ -�1�{�+����j�]-�����c�'�@ 0Zb�1�k�K�1�C�&�U���;q�|�� 82��|M����k��}���
��+Ʃ���l��;):�t{ہ���v�j��ٳg� d8  3��婪��~m���Q0 {���m����}JG��p���a�#����Ǟ��IS����w��������'��iq���_�w�ȶ����D��c����U �ˬ��H��[X4,�;赂ko�!�{v���lq�?�8�pr����r�   ���i�zw�����!�]�k�ߔ7�x�9���lR���V�T��k�ʝv���%��fV������n��hT=;^Uvd��c&
 pdJ��L��i�;mƶ.�Wr]���k��"~����;_{E@*۾}�JJJ�v�Z-\�ж��� �aΜ9r�\�k������+_I�B-�Gt?�+_�e���gr]�9�k����xy��V�+����2M�ƿ�W:f�ۘ�	_��6�).���ۛy@��p�p{[B�7��à�&�nR�y%� #��^���$�M�k����  H�=���J��um^��'��� ��pW����?~L�U.��Խ�%�N?^��b�H���ԽqE����Fg��Y-�$)!w �-�o�a������C����ʉG������x�ݪ���C�*>����*�P7���
�������m#��/����555i���6iZ�C��  魬�L��h|_���O 0���י�����V�v�ms��܍�ew�F����&NQ_�������������� "$.�۳���Ѥ��{Bۍ��'���kF�Ž��+0�*�m��i��p���ߠ�F�uWk�onI�F��=ɱ�u�v^�3�x  Il��Vs{���Ե�%�O?Q.�O �l���ܞ���b�H�{~Yy3�#OV�  �bᠺ7����}b�����㗯h�  S��k�;nX�k����������Lha�i�����xU�����u�9���9�Y���O�
H;v�И1c�b�
�r�)r��6	 HO��}޼y�η��3��PsӰ�-��c�[������t\���ݪ�������gJ�W�t���>v�܁��W�5CWw�4�_.K����_���M�f>�����δ��T  �P��u��)��>��Ox����l���  ��"ݭ�ٱJ6ٓf����پR�ӏ����$������mEO7�pH=��=o�{� ��������H_�ҍmr߱Ry����. `t�]v���C��+ν@�n��7���������ai FBoo�l�}ѢE*((P0  =M�2Ey9%  ��IDATy{�'�fE��8D�����J��#�\W~����˫���\wΧ����=���5��E{{����4�Kh�19�N4Ov���ۛ��a�ۯ�F 0Z
�����q*8�Ą�����ho  IaC��W�U��B���ߢ����䈩w�J�B�JW�`�z�W)w�R��d�}S���X4�*���� FV�}wp7v�������x��&N���C@:پ}�mqꩧ�O|B�G�HD ��4s�۫ޘ�v ps\7P��7����Z�����/Z����/��G�7k�g��r-�Cmoo~�O�ݺY 0Z�4)U[�'~�{	oӽ~�Z�~B   �гs�=����7��+�7�X 0���6+�٤tj�W��& ��'��*�E���Y��I��� ~-�W��i���Ϲ���{��x?�5�j�y��4��ܹ�ۗ.]��'p�44{�ly�{"/flgE NӶ�Yۺ_y�u����{�'/�~B͍�熉iq�������+�.�-���!0�*������t� `4�.�,=1��Hh�d���6�������紷 ����)�V�L`v�z�_W��Sh&0���=�ۤL�W�^���r�� �&Uo��/2A��F��Jy��b ~�PH������e�\W��i{I�B-�����Dŧ�9��4,�����ͮ]�4v�X=�����Km@2 �JJJTU�vP���C �8�c����V��Wr�Y��?n�����yOnހm�F���ؕ�1<jo���]�iqw������؟ճ�M�hR�����Z������v�jq����1�i(  n�hT}5�I�}]�oܦ@�T�p�ݵ����HD}��P��%���W�9�/֭L�S�f��I�[ ���p�v��'���M{\�-7������~�!ۛ�߆����Ѩ�mۦ��,�^�ZGu�mq�Q� )�?�\�`���===
�fp����P嗿i��3���:O5�]mϛc<ON��������I���O^8`��;��� ��!�������&-�ǟ��cNHx����/�"   )��[	�*���n���J.�O p�M
�7(�[w+P>M��B������߰Y�&�߭��j�L `���;_{E�K�=亊�.z;�~��n���S�� �t��Ԥ��v=��S�={��~����  �mڴi����w���S �T��Z��x�6����O�Ƅ��QrH��+Ի5��m���n&�O�|�������ٸ^ 0چpO��ʯ��}�����   �],���m�D�hX��ە5v� �H��mR�2�-w�R���o�jW�D���(�(�hq���pߝܳ�NW���r��ʞ6�� ���! �mٲEz���u�g����&w @j���Ռo���U9 ���q�@���*�B͍ʝ�@�.9l��-���o�0�톻Ž���;.��b1�\�  9�n��nq/<�*8������%��   9�Mնi3S�7nU�|�\n� `��ݭ
w5+S�:���;;_ 0T�pH�Mە���>���R��J ����胚���������Ͻ@.��#�����r鮻�[���z饗4o�<�7�%c�T� ^,�۽g�t8V__� ��Z�z���Ɣr]E��.��2�v�v�<������nO�{I頷�ww �	��j��5?�z6�! HC�k�[�+/�V���nިf�8 �$�oޡLf�V��Z�K* Cl��R1���Zٕ� ClۥX����ɡ�`tE����؟Tq�E�\7�;�J��� �`ǎ*++�C=�K/�T^�W��� �j���4f̘}���ۙ� ���m�������J�����Oj�o���ö������ �톫ŽⓟR{��� ��#
��A->������l8Z�O<EKoo���ho  I�iW��S�.�RC���Ţ��k��B���=a��r	 �"�\�L�nU��[�@�  ��,g?P�ݝ�3�����- S�Ar�x<z��u�'گ#>� �IVV��Ν��|oo/�� `?�ޡ���!�I�|>y��Yv��\��ݤq�|q�[�M{��K���v-}T�o� ��#��l��{�jZOđ��W^�̈́��ݲI͏?,  �d�f~�w6+�˗% HT��.���h8/�-( $*�V��MNj�%ϸ� ���5�Խ~�r�����_�����	�$�w�Vyy��}�Y͙3G��ŊF�4@��?�|�4;::�`?��s���?��Aݾk�k�8�e[�o�A���	mw�-�f��"�����! H%Gp�;�������HZ܋N��!�����紷 ��	u4�b
u6��`H�3V�y��E��Aceg���H3ނBM��J�/9V}۷������w:3�}S��ɠn[��2�	InܸQ�/�#�<�/�P^��v` HUUU;v��mmmv 	ON�&~��*8�D��T����g�\Ԛ
��s�w��FN�iq��#��n��?wY�۵<�[r ����z{y�����n�-�_��շc����   �!�W��KNaZ�	��pW��"��$ 
'�ў6�"a�<��6% $�˥���I�'�l��L���3>`[������S��n���?ߧIW\)wV�;�.�ֿ֪>& uww���&�2w���_�QG%��M� FQVV��Ν��|0Too� �HM��_����_�̘��z�͖�c��?ޮp{�����؟4�_��N�~'昵��?	#���G�Ž�S'�����k �fx>92-���iq/:��A�6���_^�X$"  �d�t��bs�pR@���{�'�| ��T,��� $��[:�iK�t��[X& H�S���p��i�����߱�����_�̞'wVV�����X�xw����G�����?���2Uuu�ƌ�'�xBӦMS^^�S�bz� R����ޚio�#�;n_�}Y��jⷯԄ/S��Q����zr�~O~�a�I�~e��O͏>h�����vNq[*������.\]k_ ��a�F���˯H�{����Y   �bB�N�(��i��Ez��il��o^� `���=9I�?>V��;���+~�};b��/��������Ɏ��v%�	�[����d��}ӦM6PiB���'��z
� Y�'OVyy��󝝝�Pj`���9d�����>���Ү:hB��%����������!�,��~덚���'�]�-������c��j��Z ���/��i�o���koJh�DZ܋�{��Z��f���Rǩ�4�%��H�O^b���}  �D��ڌ����K
 ��w�X)��&� !�ۯ�+�������o����}��4����߹C����
[dZ���+�ټA@�kooW]]��zΜ9���xU���Ϸ��^f�������ݶ�cy���vÝϊ���w�F%�i��~c�r�.��������Ja���z��_�y���Q"-��_J��j}�Iu�Y�T%V������n���Z����#Imq����۫�����"��	�>g�,�=�\�����Jkي��  Ø ��D�]�$$���2Fh@��8VF������pG�6﫚����-(��m������bjXv�&~�^�p/-p��[����X?��*++m�Ҵ���"5 `��n�/^l'����* .Ѿ>m��2��ٯ
��?�g;��ݥ)�	�s\7z���W}�{	m7�������������ʢ=��w�=c�RM���	�>B��gX�����5����^|�Cko�Mj����Z�Ι?�ۛ%pv��[�N�RA�Gϱ3�ѿ�F F^��Q�7G�$�Jl� RU,��e�é�� �8q��FX�@b�8V�+���'U�KW��ϳK�gO����3b����G��_!����&���؟8�i
޼y��͛�x@���g���&� H�in/(x�\���S�Ǎ ��)]���T��sTq�%�l4��w�T��?�Hhzh�&]q���fC��=6d��S{�Mw��u�������[��������疫k�kJe����n�7o�rfα�����	*8�=	mӿ{� �1����'Qφ7�3knB�U^��÷�����D�����W��33�N}ߠooa������F�-�j�*��턶	57�7����e􋥗+��n�& #8p��h�7�$&q�Ę�� $&u�A�@2�q��r�m_+<�$U��JN;S.�oX�{�j�y�%�tvh$�Uw�M��?���U68IKK���/���N8�y�^�)} ��)++Ӕ)S��7���h1���N��q�=s�*>u�J��!�|�{\׳�Mm��%
��h$���]7�JU_�����
��	����������>����WZ���S��+���ؚ�.��������g+:����)���)x7�[7	��p7��_��f^�X�{���Tv�'m;���}�R{}�v]Mʷ�����q	n3�[?T��_u��N�%{�;�Vy��ڮ�� @�qf�y�~ Gȁc�#�> 82Q��cE��WHc���_xޞ�{�%����&T�7��~��(�uߎmj��cj~�A�F�����~�Ho��|�,��l���� ?�D��ݴ?��Ӛ4i�ƏYD�	 0�����hѢ.3�� `$t��=m+(T�ig�����U9Q�2s\�N���=ݶ��e�㶜5ق���V,T��>i�e�ǆ�1����>����7��{����ISUyٷ�>����:_U��g�ZE����'V��c4���i���I��h�O�V�)�'�],J�V}`$�=�����eL�x"���*�ǔ���;�5oq��W~�	};w���˔�_^awdiv�3|����|࣪��������@+��P���*=��v�U3'�,o��o�� �b�kH����3�ù8n�+$��X	 �*�֪�ew�S:3�z��nN�ә��7�|S.���߯/|����
��� ��p�\Z�d���:::X5��3���ў�Z|_��	����~��4���u���ڟ�U\^��O}����O���M��0�����w��BE'���v�g�豿ٟu��O+�P��������Bǟ��|Q�ʉ	߅y�Ѿ^����?���hpgg���&%�nf
�%,f�"�w���+�ɼP�YC���e9Fz��P�0�ߞ��g$�m����S�0��-O<"`�aO���l_�j����r d&��"��1\\.�  .OrAS�����ȸ����r{+ @�2˚��|��'��}H>�φ� �c���*))�w���_���  �kqO���ؓ	}�|�9��?u����E�#&p7L�|��fO�"]
�1t��2M���T������L5\�'$�ӣ�'Qφ7�3k?�p{�.5��^���;?��{�i|�n;�H7fƔY���3��~dw6`.�Y��ON�"� AN{��H��7' @j۱c�����r�J͘1C3gΔ��Y �Ayy��M���Y!���M  d�HgǞ��~gHۻ��#z��ߤG{�^͏�I��Ì��F5���B��[�H���]��1�t�Ɔa���}b?�0M�3��A#m�uW+J�ն��V輅���L6K� ݙُ��c�Z������ܾ,E��gb�pFg	" ���w޸��3VH���q���  @*3a�6h���z衇�/|A�����H��������E�pYkk��Ѩ  �d��ިq!��#�������KJ'��~���zM�ޏ��v��Z��Df��ٿ�C��R9Aߎ��r?I��j~�au��F�sh��UoW��(m��j�=�Jn�2Ѯ�U���Ҟ�eC�-O�%�c�+ 0\Y�Rg���� $�ȕ�x+$ȝ弱҉  @�����֭[m��}�ݧ�.�ȶ���	� ��x�t�R��k����V0  �δ���W����܃Ə[v^�3����oR���+{�Le��o���Uu�wn7Z�}jX�'�kG�������w=d�#����J�����֬Ү�	_��2M��+�s2�Y*�����u�� Ó� ���� $�ic��Ġ*�#�	���r9*$�Ŀ   =��թ���~��O���|>aL ���竰���Z�"Fgg��4 p��7_���J�S���㙲���^Q:2y�����������M����~����X$,d&�ǣ��HN��-S�܀{\����ո�~)���ϩ��G��v^���[��g3E��N�qi�N< 'g�� ����I<9E#6�@��d�2�Zg,1���X�@���X��BEz��v�  d�n P�2��͛UPP����0a�.\hC�!>�A�:u������7����&��  G1Y�-W~K�n�O.�/����Ԏ�~�tֵ�um�ɕ����B?������^�V�\�1���)��E���a���܍W��r�.P�q�I�c���黗�}:33q6|�s�w��ʍ���]��M�/=_����dѾ�����7X �τ�L�1q�Y��1������+��,'��2����Kpw���  d���|��L
���a���6�������L�ƍ���� �٘1c4gΜ.kmmU4�R  ����K���ה�iRg돾���j���{n��8U~���;~��jzh�2Y̬xf����Ao��UFqP�0�ڢ]�]=l�7"wھ�b;�vs�����K.����	̌�7.9G�~s�
���k�����?������vnO���ۄ�׻u� `/`��(�^/' �`���ᔀ�����}��-r�\� @F�Đ{WW��nݪ3f��{���?�yegg�p&M 8���-Y�$~��q`ww�2m�  Qw�����jⷯL���\w��yP�b�/���=ݚ����{˱����?T{���t&;ܿ�F�ʉ	�>����pG{Ʒ���![�j�,���B_���5���Q�?6l�k������|�e���<M���Uq�EJ7�+_��o~qؖHuf	;����XHo��&��xN �?_�8G�]���v� `(|Ec�W�A��%o�X�P� �>�f`���  �|�r�������-[�.�@>�O�`�`` f��c�9F~��e�PH��� ��v��+��Z5����;�;�����������i�ϫ��Z�~�sy��N����߻\��>%�h~����u���?g�3I,Q�����O+S��	[���:^yaX�w��F��W��EU��B�����DǦ+.S�.e�h����v0�r�O�M����������:�C�}�Q�����̫oxכv��FM�/�7��m�4 ؟	��v�U,��KJ&��M C��ʗ7�P�ve2Nu�� C�r�_4^�M;��\�|�  �)/�m�!�Đ��-[����m۶���)��b�����@���裏����0�dKK�%  oi��u�}]��+�̘}D�nm��|C�O?�L��؟յf��P|�J�O<����o
�9�4x��7�Ze=W��w^�:?��������d���(#[�ͤ������_�۰����������_���}K�g�/wvNB��n���JM�AJX�u��j_�l�g�i���ʪ��Tcf�4,�K����D�f�������v����[��+��+HS�1����Q� ����f�`Kf-�t0q�O����%Up��2V82�Ҫ����'Ho�  @��j��q���А�	�_�^�/���?����kƌ��� {̛7Oeee\���l�Q  ���k����U���T��o(P91��#�]���&���u
wd�gqFM���҅*<�$M�����S�=���N�ߟQ������Njn҆�.���o���d�ۘp���վ2�)���5�7�[T�L`2�&3\�˫l�O�c�J���4k��P�W���L(~���[�X�	U����=�P����յ�5����D��Tw��Uw���_|��uTp�qʞ6sT~�̀b�ڝ�^����g��ߣ�������J;y��;�<{����p��|�5�tv�'�ӭ����e�" 8�@�T[k��*�Hނr���k�/ ��WZ%W�F��a�ۗe���Hxr���+Q��E��tʦ  d�SC�R�����x��75�|-[�L]t����{(�Վ�0�N��ɓ'pY{{;c$  ��D�pߝj��n,=^���Q�/:Z93g���t۰z�mQ�k���_���S����iLs�9�ǍW��>��cOT��
�?��hT����ߤ#�=5��Qkw��:_U��tU}�����ȓ�g/��Cj�۳�y�O���:e��W^���'�������?v�҉�B-M���홿���G�$�d���^&����=�d�6woa��y���)�ަ�	�X�ʊ�:W�lO{yrr�����K3����0�z@�+��'O^��L�?X�˾�3�����]B%���f� Ov�|
�'gv�h�;] p�̊����ݨL��&��������Fo���r  2�	�����S36���֦;v� �=�ܣ�}�s*((���U8̪� �k�ر�3g������  xѨ:^^aO�	��\ea�b�=Y�Hg�-��&H^{��d��~y�����Ǐ��*��ƿ�a�j�����}W�������Q��9����:m�ɕ���,����O�pfx��3��AsR�08�Yڜ�Z�ND�f焢�k7�	� 0��ؙ
�7(�j�}�c��- ���)�o�fg�g��^��r� p8�²��W��ݭ�(.����  p�S�]R���w�ܩ��=tw�y�>���*(�)��%H 0���-Y�$~��wY0TG+� 0�3�Ps�=apL�<����	)��.�Uo��E���	��rw  �t��)�L��M�]�gD��ʪ�/ .�e"{���\�L�]9�6��pɮZ����`T��*�*OV�  ��8!�a���~��ir���m��A�������c��{�U�ѨZ[[3��   @�p  H���sn�S4�KO!H;�eg�4����+' N����LR�q�2�Y�"@{;  ���!w�\�~��:�(�رC�<�>�ؐ�	tFGx)o ���:����������q   ��p  H�ǧ쉋Խ�e)��HL�*k�L��s)g�"u�^�hX��6�O\( H3y2�٬H_�қKٓ���-I  �,�C��`P�֭�!�U�V���X'�t�z��h.���*&ܞ��u����ͬd    !|�  �$��rʦ��a�ҕ	�L9z߇� 0���\eOZ��m+��\RNբ�s� $���Qn|��s��������3��#  �L����ؐ����3Ϩ���~m����d*�Zű����W�moo�c    $��;  @ٶ���;��n\&�9i�<�\@2���+Rު��mJGY3�+� $�;+O9�{�ki�B���ɪ@  `?{C��+������2)���ѡM�6i֬Yz衇�s�<y2!w ��M�����˻���    Hw  �dr��;�um^�HO��IV�|� FL�����C
��(��K')k�M #�W<A�񱲷f�҉'�H9���(  �gC���26���Р��,M�4Iw�}�>��Ok�ĉ��d�ۭ�K������{{{���)    
�   I��x�;�8uo~A���x37{�l�L ���6�"!������]�@ 0�e����n�ҁ'�@y�}a��# H5/���EB�8��U���	Β�!���jr����=�ܣ/�P�ƍ���S("� ��\.}��*++;�r3~���7@��.��%B�X�ۮ�[ ��"�  0�>��f���m�(ܕ���U3�r�c&	 F�˭�)Ǩw�j����L�4�r� `4d��%�7���u�s����*w�1ryx@�y%�X.+b�����q��\:��Up�L�o޼ٶ���;��E]dà���3n_�d����?3����@�]����1�L)�|Y
��MN�j  G�O�   F���S��Գc�Bm�J5&x�3i�|���bއΩZ �/����J����.0n��*�	 F��l������uŢ�q�]�Cn�  ՘p�����S��71B�Γ�!�h4�7�xC��Ϸ�o��6]|��*--�!�`0( H'{��ǎ{��HD---L��t��S�������� G��;  �r�=ʝr��-5��8�*xr
�������Q�r�vb��۽�5�©d0�q�LZ"o�@*����q=�^U��C)��V��9
�M �"���������~���А��u�`�{���o�%�\���B��N�;�t�v�ms�@����&;�@2nO�� G��;  �(�TʓU�����i�o��VV�4eU̠]@�1A��'�g�:�ZGq�מ&�	s��� ���U�̓�_�A}[�QEysK�=qA|?7_ ����B���޷��31�nk׮=$䞛�k��	�Hu���P{ss3�v IG�=�r 	�   �ēS��Y�Q��Z}�7(٥���ʩ�'w��v ����R��*mT_�:E��F��=�v���
 R��LZ?G��J����pg��>�/������'�U8  nO?�ܝ-�C��p�6�/\�P---6�~��+++��;��f��K�.Uyy���1����p;��#ܞ�� ���;  ��r�_:I��*[w��v�����>�iD�7K��b@����7����W�)�_�`{�|��%d+� ������+�ݪ���
u�+�IN�/[���v��j@ R���E���29��z�ju�Qjhh���]x���˓���r�J<�q؄������p;��@�=�r w  �T�v�	��T)�^�`kM���Rlx�v����]i[==4�H[.�
+�+(���P�N�j�Cexx��㓿x�+�L����z��}]�o٩Pˮ�D�r۱��[��c��:��鏐��ez�}͚5��݄Co��V}�3��Ϗ�;�TbƤc�=VEEE�\��ԤH$" H&�홁�;  Q�  R�	���X$�pg��]M
u6)��m����x|��ٶv_~�<م�� d��x��+����
w����&{��u(6��(��c���XiO9�v� d
wV���ω�f+��n�I�_i�6���s=����d�/K����� =n��ܝ-�C�}}}Z�v��777�&wr7!RB� RAVV��;�}�����pxx�' �p�gr7���vr �;>�  HQ&��+kO����~��G��.H�E�R4b?�u{�un_��,@ry� 'p�����<c�\`��P�+
*f�ɷB���X�r�Oހ܁<��Y gp�ɏ���n/�����R$�?��V��2;�Ϟ����W���ϑ��!��go����xB�!����^�Z���W[[�n��f]x�*++�!�P(���U 9996ܞ�{રf⍙�C�@�n�LO�ir'� x7�  ҅�%wV�= Ì��l{ ����� 2���e�Mz�ɝ���dz�}͚5Z�`�=�m��.PEE�|>!w #���P�{�����p{SS�v IG�=�r w        ��g>B�Ζ�!���^�����B��z��?�|UVVڐ�	�F"@����kɒ%�z��n0R�;!w ��!�        ��v� ��l�r7���ի5�|{���o�y睧)S�ؠ���"X
 �����p�B;��Ϭ"���� ��;!w �;!�        ��v�!��l���@f__��Y0�r7�鮻��Yg���s����9�B!�p�9s�=̬a��M� ��p�3r w        ���;!wg3!ww�v=Y1y_�=//��?�C�!y͚5�7o�
u������Q��r��n��~���b�| ���<cZ�'L�p�uf<2���$�vg#� w        ���������24�n�׮]kC�EEEz����ѡ}�C6�����8bYYYZ�t�gfV�hiia��t��ar ��;        H;�۱!wg�䐻iL^�n�f̘���r�Z�J���:��s�5�Ӭ`(�
�s�����_�����$�v쏐; `�       @Z!܎�rw�L�oذA����4i��mۦ[n�E�����m�{8��� 0X�ƍӢE��yk��_OO��L �F�!� ؋�;        H��q8�ܝ-�C�Fuu�mT6m�����馛l�}�ر�z�r�ݶ� މ���̙3�X2���uww ��p;�	!w �A�        ���x7�ܝ-�C�&�nB�s��QWW�mr?�s4m�4p���6��1J8�#/^�����omm͈�@�#܎��!���ȩ]M 8w        ���c��;�	����ɱS����{[[�^�u͟?ߞ�뮻t�	'��N���{C��hT �Waa��.]����C�3�bZZZ �F��x"Ϥ,B� �L�       @J#܎Drw��C]R��{zz�j�*͛7�>�+V���Ig�u���|>�"���� ���R,�7�ό���L�0"�c(��sp        )�p;�jo�=��B�N��!wӴl��gϞ���RmܸQ7�t��=�\�����l�Mxմ3p��kW{0����Ь
�`$nǑ � �D�        �$��8R�w���=M�ܝ'�C�qy�������ĉ��Ң�o�Y��G4w�\��n��~�B!ڙ�)((В%K��y���Rgg� `$n�p � �C�        ���.�ܝ͆�k���qS32�n�����mXu֬Y��e˖i۶m��>`C�>�O�HĶ��|�'O�7��`f�0��0�H��1����p        )�p;�!wg;9ܝ�!wô����k6Ԛ����+W���Yg�}�=o��	��6wp�y�k|�ҥ;v�כ�.f�`���B��@� ���;        H�ۑ,�ܝ�	!w�<V�Z��ӧ���B;v��7ܠ��:KS�L������Vt�9L���������~���2���!܎d"� �@�        ���H6B��愐{4�ƍ��ѡiӦ���Kw�q��=�X�~���y{�^�5Aw®@�3�i���;����ӎ 0R�c$r��G�        �:��)�ܝ�	!w���N===�={���^z�%m߾]���m˳	��6�P(dC� ҏy�p�� i0<�z�R�im7�s )��1��@f#� U�yc�5~�      �Y���˅�!܎�F��ٜr7-�V�Ҍ3TRR���z�x�:�3l�����lִ�H{[��ڶm�~��}��X����* F�v�B� ��� FU��;�+     �t֗U �v�B��攐�it^�n�Ə�ɓ'���qmڴI����s6�ߜhsR����fr�������/�Ul��� �$��M&�n�����; d�        `Tn�h#��lN	��wﶡ�ٳg+77W[�n�o�[}����is7w���H=������O��ZZZ�y��mjj��U `$nG*x�&wB� �9���;��a�RIo�4�      NC����������v�7=�C�����^SUU�&N�h��s�=:ꨣ����OYYY����ې{$��g^�f�^����O��_�7���U7n$�`�nG*!� ���; 8ȴ֭��+�P*���W�Q      p��H5�ܝ��p�䐐�	�VWW���C3g�T ЪU��y�f�y晚;w���ަh���.�˾M�}/�������qϧk&�}�v�J �4��HE�� sp        #�p;R!wgsR��hkk�m�3f�Pii�����l�2�^�Z��UPP`õ���ÌC&ܾ��l��s��^�7餽�ݶ�g� �nG*#� ���;        �ۑ������O$��8N����o��1c�h�����|ڴi����z�z�:�c�5H���	�G�QH��n^s����u��c��@�a^�;v�Ю]�Xa�� ܎t@� �w        �t�ۑ.���#o5�rw��܍��&��:u������߯�\�֭Ӈ?�a���ٰ�	��`�	������$&ྗYY���D��:::lཧ�G 0�#�r��F�        $�v�B���Đ�is߰a�4c������o�I'�����=�ga·~���;0������y]���Z�|��pbD"UWW��`TnG:"� 鋀;        H��م�ۑ���ܳ�_-�i�ŉ!w����k'M������P��>��+W���Oׂ����M���@���b���3!����/����wYss�6oެ`0( -k��	�#m��{N,�㺙� 鄀;        H����H[�ww�/K�'rj��ַnݪ��F�枛����N=���z�Wt�gj	��{��M�ݴ�xwf��y����טil_�f;�v�޾e�p��Vm���#�m��p��B�          �Ԑ�a��������TYYi���]�t��7�&�3�8Æ�MH����P.Aw��
�������w�X��~m��Rmm��o��
	    ��;          ��C�&h[]]���:M�<Y��իWk�ƍ:餓t�q���.Aw``�a���u���k�����L�W{{�mm���    8w          x&��ݬ�r7�������ԩS���o��	�\�R���5c�{۽Awp7Awx��p�v`_�|�}=�e^O۶mSSS�     �         �]�V��SC�FGG�V�Z�1c�ؠ{ PKK���nM�0A'�|򾠻	���~��p���w��m��&ȾW$QMM�=��    ���;          !�=L�tkk����l��yw��e��:��S5e�{[��p��ۛ����3�h�����744ذ�Y!    p �          0H���0��۷oW]]���Vw�4Q�~���2t7�wc���ٖ�jd
�mƂ���mmmz������l7�C�k���K�|f�   ��p         �r�y����<�I�&����^n�����O;�4�?�^nB��d�&�nN@:2�Ǧ��� �	��X�B�V���ٻ�(�{���d_H¾��+�k+j]�G�ֺ��؞������9mmk�ݭ[W��u*j�
";B ��'���qh ���,3������d�'�L�y&���9l!GUU��[��w   �S�         @r?��Q��JKKӘ1c����n���c�=��S��SN9t�P���mX����
���n��`{AA�V�Z�|4ol����޽{U\\,�?1�  �N!�          �@Ƚ%k�޼y����5~�xedd���m�ܰ���4cƌC�P`8���<D{����Gj-�ns��}��v����'&F    :��;          t���}�������ܛ����ƍ5p�@�7�ލ~mX���E�4{��C߷P�������]�)&&�='c�)[`}ǎz��];{s��n��"��P\�E    ���;          ��M5���=���r7�ѣG�FwSRR��^+W�Ԝ9s�p��C�3�Ŵ��������بM�6�`�=�����q����b��8$�#    �@�          ��5���{�JKKݰ��ȑ#������v�z�j�Y�Ƶ�[����CBAc���@wh����"{����{jhh8l��srr\�hΞO��F   �8�          �,���ߥ�O"�ފ��jm߾��G��aÆ����պu�~�z�;V'�x�fΜy��ha���87,����� �E[m�b����9�m۶�Z��-�ؿ�***����   �8�          �E7�*.��%��&�^�ڵK{��q!�ѣG+11�������K/��B����s��4$vGGY�=��n׏d�06n��\Xs{s�|+**r�v;� Ж����`�   :��;          t��M�!�v���������C��V���T�;W֞mcĈ:餓4k�,	��-o!w���Mۀ9Z�ݞ3��k[�nm�`���=ǀ��3NL�5   @�p         �.FȽc,P\PP�Fzz�kl��{�{�����^˗/w!�ٳg�0|(�l������B�ƞo�6mr����ޜ=w��ݞ{���<��!�Ǟ3��M   �q�         �X�ݛ�K/r���J7v�ޭ��Lv8p�����x��=--M3g�tc��ч>�Ȱ���ʍ�'��[���P{EE��mۦ6�F�#544������9Eg%&&*���v   ���         @7Y�T�8��;�B酅�n���j������R\��?sWUU�w�q�Z�g̘6�j�6r��_������i˖-��=77��co[K�����xn�����܇�   @�p         �ndM�"�~Ljjj�k�.eggkȐ!��=##�PK�5�����q����_s̓�bnxGthho���X`}�֭ڱc����6�nϫ�"
;; �����ssvC�    tw          �fr����#&r?D�]C�!nX�{(�lܫV�rc����8q�&L��I�&)11��}���X���w�N�wdho��/k`߾}��������܋��ܨ��Е�9�����@��1���   @'p        �"���Zx�$yb�h��К��TTR) ��[�X�ܻ�5n8p����������,��R^^���׻a��cǺ���ɓ5t��������i��N���c`�=�vc�={��v��XohhPqq���t[Dc�����{�3�h50#UKL����:;�Y��n�� �HE�        ������q=z�b�Zeg ������B�8��.B�]���ɵw۰����[�=--��>֨����Ɗ+\��-�n����CBA����ޏM�0{��h�q�����ݻ��hM��=v/--UII����x����y���⮟R], �k�4e��iT�}]��o�������J40#��;  �p        �J�:��o��?���� ����}y;�Ʉܻ��u�߿ߍ��4H������?�[�w��݂�����1c����n�#�ax�ۑAvO;Â����{���v{Lm�B8�=��4j���Г,�n�op�3v �r�:����K!w{��`k���J @�#�        ���Rȝp;�-,�K�{���tAA���Fw�[�=��6��6pk׮u����#G�����z��{�&�暇ݏ}ё�����ծ�=7�"j�v�ڍ=����*++s�ށ�`�g������+
���C!w�� �hC�        �;�;�v�[Y�{L�.���{�5|۰6pkw���P�{||�a�[�z���n��B�ÇWVV֡z�t��wk��#/{[���yh���:Â��yyy.�^[[���Xؽ�����?�B�g���Q�՗	@�B�� ш�;        @w��;�v�G�m�US�N�0b2!�f�ߡ�v����B���>>r���`�����K�M{��ޛ.o��u�ͷ5���X544����}�C�v�n��ګ��\���v=�G��l���Ǘ(��(��Dqȝp;  Zp        �N�r'���E�:�����܆��=\MOOw�w����9�s,4VRR���͛ݞ�����Lt��4h���������f����R׬���FMMM���XþڭA�@;"]rr�;��SW����}V��]�}[���J @�!�        �ݢ)����E�ہfM�
r�Ps]]���=�Z�m��cb���SSS�V�v���݇�-�nx�؂�6�>���z||�z���u��[P���]��6:��w�9v�6B�e_����~^�=�//�Q� �iQr?n�$� �N�        zB4�������Y�ݗ�Sύ�|(4m��P����
t7���t(��<��V��m��C�y��Х�jCM���������߶���͟C�����s+4����?VZٛ��@���v;�CȰ�B�c���(�n ��        zJ$��	�a��N�4�G�P8�����m@��yk#\�{80��t�����}�9�~��755	�K����F�U�@?�!w�� ����;        @O�Đ;�v ���������֍p�m=v��uv�kc5��eo������ky��]vE�;�,
6���^}�([���@?�!wn�Z��*�� ��G�   @��*��/r�81ŧg	 "���\��E���Lyb�  '�B�.�^�ښr�4��m^�W���n���P�=��vx{Nx>��m&t{�ca{���߳��}��۰�l�1����-%%��C�����vk����ߊ����-E��f�2 �o௛    �T��^~_�F����q�E�HP`��Ah��S��!  �"!�N��h��#B�4��/�X[K� �������C󰱟͓�j~S� �srw��� ��         ��7C�ہ�`!w_�N=7b�aM; t+Y��v�f�U;#�����X) pz9�N� �p        �M�:�����أ_��!�D��:���N� �OBB��gcbb����ii�n��T# 8L�N����5���{c� �$�         �������ѯ�$	@��&w�.=K� �Mbb�RRRͳ����ty�n���	 �q��x_ @W �          Q`~S�bhr�.e�ۓ��Z4�ڧ�Rw��U��'    ݏ�;          D	����x<���+..N			�5>�OSJ�u}m�    ��          E\�{�.�m��!wk�z� dav6?Z���L�n�M|E�n�8���&   �Y�          ����lrOII ����T���|-n�   ��A�          ��kr�ߥ�5� :���+��R�Ujnpn   л�         @�rALB� �aj�����2]X_�A�    D�          ��@���^���Q_����Z�T�T�_    "w          �rrO;�]{� �R�>�|�rL�II��    D�          �L�5�     ��                "w                @D �                ��                ��;                 "p  �"ޚ��>��W+�kr�c�������            @4"�  Ћ��%j(ة��|5��SSE����By+
�-w!v_p�j�}�q��\���qiC������^����J̚��a��$ �o�����h��9��88_�����"5?���|���Y%S���u��ĺ�@��$�)6%Í��C��Ӈ)!s���r�6b��@4�ŏv,�T��1m�l*? _]�#876ֺcK_M�}F���΋1I������i��ؤ�82~�HwL���_�         t�   =��p�j��W}�v�������ܻ�kz���N�<%��a��8|���#e�l��?Iq zCci�js6�n��n�͡����
�;u����Y0�<��i���((y�t%�>NI#�)i�L7zb� =�B��In�����d�v�xҎ%GL΋^��Ĭ�̑         �0�   ]��x��w�Q�u��^���h����Kr���W۔0d�Rǝ����1a�Ҧ�⚍�+Yx�j�������r6�6�=y�Ki���*�h΂��cfi���Juc���# �
ִ^k���w�\�.�mR�۠H`����Q��öy��2�xw,�:~�����v         �5�  �QSy����R�+T�i�k�ԷQ���ck�&��NQ�qg+}��K* h/A��lpsf��U������(�Y������sw����N����<�~�Y�'��� ��W[��ɪ�o�a�&>��Q���|�(��6���?)8G���I[D�4@         @a  � S�*?�����]��/WCQ��Lݿٍ�W�<�����s.RFp����b -4U�b�K���Rp�|E���u��n�6���+��i�OW����1�%Y�; |��Tm��*�{����<�R_e���o����w��Т����Հi����         ��  ����X��=�B�_����ۿfrr���Ҕ�����$%&&*>>�]o�n7��|�������N555�FSSS���C����M��q��x��.���* ���3���Q^T͞�=�͏6'�e\\��G�illt�]��hs�͙��W[�^?l���S5h�27R'�s� �/vlY�y���}687<�ZۻKLL���ӕ����E�������J�46wڼ���{ή��?4����VUUUn�<����z�[n���[�0؝�"#xL9褏�EB         �_�  ��W_���Y%o�VU�W�����,6L���n<�]Z i��.pԕ,�T^^���2wYZZ�FAA����UYYyL��,Rɪ߸a���']��EW�л'>Q �6;�C�;Ϩ��U`k�޷-�:t衹24l��m6o��t�:���]��.KJJ�|i�������@gW��߮�g��FB��w�-�BiSO!��aj/]���<��������X���G;����.����8�͑�OW��Ҏm�,..VQQѡK�7;���[<F}�n�KT�qK5x�UnQPlR�         ��p  h�$+�E%������������E�ƍsc�ȑ1b�YȽ'Y���6±F���B�۷�����uM�e��o=�Fl�@Hr��J�~:�M�i*�S�?���n:�����c�j̘1n�;�Ew5�0S�L9�m�ʕ:��\���9-�Z,d��m2n,٧��r#1kbp��e�z�����竫Tٺ��c��M�ݱ汰�u;�5j�F��͓]�0�=l��;�=�͗��A6�2;;����w6{�C�~DC�\���ϕ'�_k        �U�%  @0�Q�?~���SSEA�����M��?^K�,q͙��S�o�b᤼�<�ڵK;w�t������r�}��4b��.�MCN�Aq2 ���,,hX��#�x��N�5-PnM�O�0�6m�'����չཱ�A��h��J�[kqh�\��u�������_���|C�3NW�i7j����Y1 D��]kT��a����[��Y^�<y�&N�����ÇG�<�͗�EJ���;t�͍t��}�v|�O[xZ�֓nħgi��k�u֧�4r�         зp  �W �����?U�����fGY���6���kJ7��j�V� �k/6�T�e˖C�B��U��M�~�9�>�e^p����)�M;U "����|Y���j,���Ϸ�Қ�gΜ�B��LNNV�[�v�[ ��+��F���B�t�EB���n����*7�t#�ן��3oѰs�Rq�|�U*]��
_��j����}��3fh���nؙ���!C��1�|�quu��mۦ�[���J�7ۣ��P/�ЍS�h�y�Ѡy���        �G�W  ����T���*x�G�?��ßo���cǺз�R&$$���Io���N>�d�%�\�x�ָi͛����{�=��䴫�3�mP��߻�:q��_�_4�<1�Yjs6�p�OT��_��Tߡϵ �q�whD[P���\;�����a��067Zp���}�����̗v��翧���9�g��� r4�U��?P���__��Ϸ3���={�kj�����2`� ͝;�cs�ƍݰ�-:���o���9�5�=�ť         �w  �oX�ȂGy�ݯ���\(�7�k�l����]3��w�"`�3ƍ/�Peee.�~�z�ر�]�͚��Ү}L�C'h���T|�bR�v+6���P��Tk;?�\X������m�u����^6_fee�1o�<��չ���ݻ�B���8~������i��_pg'F zGm���}������/������,М9s��Ad��K�.u��dǔk֬qs�ю+Kr��̗����OCN�A#?�%-         D��M   ����T���H�<䮷��-|4e�����^l-�g��?�v�{v�g�Q^^�BIݹs�Q?��([9������~��5�ܻ��* =��OI5�k��9���:���p�B͘1C���6�[=--�[��^�N��Fcc�����=6�0����~��y��9Ѓ������/ =z��ϟ?_��f��g�q�%%%.�n�����ڙ��^}X�o���G\�E%fM D���:�74�����J����9�u    @�*+kU_�������u� �=� @�e��y�W/�@���v}�5��������Zz��?�6�P�6����w�q�Ѷx������*x�q闔��S��'
@�r��g��Ϊ�^� h��Ů�=))I}�ƍ�-�~����C�=���.�u�V����(�n�fe������~�݁nV��m���}��������}ѢEn:'33S\p�{��uǕvohhh�s�_L�_�Q�}M��&	 "�G��5ړ��W�zzz�2ŋ,    t�Gy�ڵ{W�|�i�Dy< �� �  ����IE+����*
��LL�&L��iӦiԨQ�7�]��ߚ��l�����Yc�5�\�e˖i�ڵz�7\[q[챳F������OCN��<��е*7��ܧ���]�kkZ������̾���=�uSRR4k�,7


����{[��u�
�����xҥ�u�r7����5h�/�g�>��o޼yJLd�^W7n��_~�[<�ꫯ���5�W%�~�ҷ�rǓ�.���3�	 "G��MeeI��   �sz7�n��˂�%� �[� �>��s~��.�t4���.�>s�L��ޝ�u���s�����,Y↵oZ ��7�
n6��Ӟ�>��c�{@�\$ Ǯ>����U��ڵ��a�t��gk�}>�i��n?�}�mX�-���{}}}��[�}�Q��35���+e���y�%9������3�
��"��ӧ�`�����&q8;�?�3t�駻yێ+����C��r�`_}�݇_���?��" �]�n!�    �����B� ����;  �js6h�w�z��G�wРA:�4y�d׮�S�����z�!����O|���K�b�
���jlllu������5�K\p3i��8_m�����_|Po�Q���Uk.X����?���u���Z��Ν�ٳg��-����mu���+��W�i��˃�����9V ���X��羫���w׏Ǝ�l!�y睧��,�g�B�3f������_~Y�֭k5���?ܧ�?��+��!��(���wx�[P��B�    ��n!� �KHW ���*��
��X���}�l�Fʹ�4�^�Z��v��oC���W_��/�X�����/_�fCq��gU��e?�������& ��h�/����������w�q�袋4i�$�'vv�H
�7g!�Y�f�3�l۶M�ׯWMMM��~��_���ѯh����/ m�㌜�ܭ��=G��~&/^���H�7���c���[ouǕ/��R�g
j*;��o
�������3�N�' �9����Q�!�    ��QAq�v�ޭHC� �Wp  Q�H{u�K���_ff��͛�Z�{[||�kr8p�p��0�駟�B�voh�.�6�V��U�Ѹ�A�.��������>��ͯu_[t饗jڴi�v���AUkҷ��S��>л���|�o�Q����d��4��5`�"h��`��<z�;��X�ݎW.�����gĈ�LA����y�]���F�������v��y��Y<	�Dn�=��;    ��`�}G��C� ��   �X�� mZ��~���:餓4}��^il'!!�l�>�l!<�-[�L�{�^x��\������<�|p�2O�Vc�{Pq�C���&���;�E����&Lp?{��
����h�N8�-Fذa���}�|�����{_[���z�s�w��. rg *x�n��7ֵ��Oڱ�e�]��C9�t��[t�9��O��;�E8�<�������^��-�B �="?�B�    �p{!w @�#�  �J�_+牻䫯ju�ϙ3G�f�r������.L��Y���>�1�z���_���)Y�{UlxQ�����.�M ���o*��7�>o[��Y[�G?�Q-\�0b��G�6�`���k������	�c ��WV�{/h�'~��'^,�?��6O����Q���&�q�ȑ#��cgr��{�q�F���V^^^����k�CW�����<�6D �u�'�B�    ���p{!w @4���  @�ԝ��-.���,Y�ą�#ULL�v�ڥ�����0i{X��w��7�z�)8p �~ޚ2�y�.�>��G7 S@d-���M����
�}����.�Hg�yfD.�i������:���]�}ժU����_ci�v|�e�r����S�$E��7�Qn����(���rg�h�5�[c�ܹs��gg��E������������>�~ek���m�4��_�@�h���C�   ���p{!w @�"�   "^�;��'���},�g��1c�(Xc����	Ku��i�t�}����_o;�����&|�	e�p������V������^��~���k�\���}�]����/;v����J�]�V�6mR >�T��7.�9���h��%���������s�-vF�/�P�s���[l�t�Rw��?�Qk֬	�_SE�[4x�w�/��k&��:nώ�p{!w    ��Gy%�����B� �h�_�  @��7�+�7�Qѫ���5�[Ps޼y���U4���Qcc�P�}�1�@҉'������ڸqc���*
���jع�֘k�+O�c�}ū~����!CM��dee�ꫯ�q�'�[]]]������x�bM�4�5����ݯ�([[����su���/��*Y�{�h�W[��~3f��u�]�!C�}WFF�n��f�r�)��o���°��bۚ��Ҥ��R꤅����p{!w    �Ӈ��]�n!� �6� @D��ۦ�]��}ﷺ����~��1b��Qjj�V�^�3�8C�k����;�n�:=�䓪��j�S ���R��՚�駕�5Q@_䫫T��7��_juk���K/��&�0l.INNV_d��-[���aÆ�m��Wy�~G�;�֤��V|�0}���J9O���%%%���X���_x�;K�W��U=��Z�|��~�}��h����1�ܯa�}F �>}'��<�    }_�	��4� �H6  ��S��/�~�m�kZ���>�������bB;i�ܹ�:u��~�i��_�
�OM�Zm��|M����8�<}�[��2�����>#G��7ܠ���-y�ް���^+,X�ѣG��W_Ummm�������;I�?��L]"�/����'/S]�m�7{�l]��JKK�;�-n�3g�~��_)??��>o�r~�YUn^���|B�) ���˾n	��ì   ��#������CB!w�o�� ��Dw"  �).4�{T��'����N;M'��6n��y��w]�2:ǂh��r�N<�D������V�j��.Ҩ+�G#.�W�w}A�[O)��[寯��Z��;�<]|�Ţ��u�ln����-v��+��k�)'''�>Me���Η�Η_���{^�z�|�������J'�|� {�q�}��O���+�-�*_�7m��M��3J7G ���|����y^RV���&   @_��S��"��b_}_W��F�  �d}�U  D �z�
׈ؚ�C�����s͚��֭[5}�t���}	z�Ǵcǎ�~�r����w������bS2D#{.����U�҃��c��M7���p����~�(&�56[������ƍ�f��=8R��U����.�}���a�$� �C�]����~p�lu�)S�����233�X���W_��3g�׿�����Z�cg�����#�\�q��|>�jj    �NV|��:  zw  ����i��/qA����Z�p�k$�k<�rss]�/�������{��/���{.|���g��K4���+a�8����w��Z�<n͜9s���JMM�f!��no�NPVV�V�X������_��k�����������J�|�koo�{-]�T�_~�bcc�c��׾�5=��ڴiS����z����j(��ȏ�7g        �B� @��޶J;�Lު��-tt�)�hڴi�ˬmٚt-Z$[$p���V�GyD���-����@���HS>��R'���h���&{]��6_^y�:��3��)))����_>\W\q��8p �>5������Ӕ�z^)cg�dM�y����U�g}��0���Ϛ5K���"���K����򗿴\<�x��<�ܤ	�=���d        ��p  ���G�����5�ݞ���s�=�5��MMM����u��آ�/��z�ᇵ{��ۛ*���Ԥ����������B��%9a�[H���nӤI���ٺuk���$%%��/��ի�y���4����o��/�	Η��D�xm�w/lu�46G�\��>:���;�<�(���W]]]�}J�~Z������?+>��w        �N� @��{�;�}�K��0���L]p�.��_���;Ｃ�K�
]Ú�?����w���o�W_�߻Hco�������HT��+���+��5�ɓ'��fFF��~���n���3_��R,���[o�l(և����[~�!����HR�y�v>�L���V�Y�d����Z���0t��ٳ��/}I?���Þ��z����E�v�r%c�        ���z  �g�}�^�=w���=Zg�}���X{�fF�)t��p�3f��y��̀���$�)ӈK�$ ���V�~�1����n�P�6ccc����ɡ�9�Y�fi��z��W��z[lx����*Ѱ�S@$����?����p|��u���6l���^=��#ڸqc��E����gh꽯(y�        �s� �
��e��L�>�6-��Y{ӦMܻ�5�gee闿����[��s���|u}շD��տW�/nP��2h��xt�����۾};��?~�.�����˪��m�C �����/+5r�������T����̓�Ύ��O~�_]%11Q��~��~�i���k-�7��j�7Nє�?��	         G�  �k�����T��Z�gΜ9Z�`�����Lr�&]t-��~���C=�������N����[zS�?~��O�i+�Zl���wg%�?��q������Z7t�P]v�ez饗TRRv�����Mu,
B�)z��y��a�Icgi�뮻�\��f�q�������?�A~���Cou��}�M��_�>�l        �c� �ng��qC����s纁������z]�;��ݾ��/�?��
[l�{�ۮ�}�?��l=-���jߓ_��ڈ-�9i�$�s6l����h[jj�.��R�X�B�����-
�7�k�u?`�D�*\�c������ؙp��n�Ԁngg<x�y�555��__�\�)�{V�ǝ%         ��)  Э\��g׫���Z���O������z��u�)�]oȐ!����/��.�Y��g���k��?Г,��Z����|�3=z��9v��cg�����l�Y�&�>/�<`�D�������[��1�p;z������o���s566���X�|DS��Ҧ�*         �w  �}�}�v���d��X�{�̙BK�GUUUJKK����?����G?��v���b{��)69C������P��_i�?v�-ʰp{VV��y�ׯgN���D�t�M��}�ʕa�q�e� �Z�uݩ��'�n?���UPP��;w�v���w�q��O������P���_@�        �� ��a��_ݩ���lu�E�noCRR�k�=묳���B�?��O�m۶�������}^@w*�ן��[�-�>܅�lQ:���N			B���l���n��UW]���X�X�"��������?p������y2|�}̘1:�sw�W]��n�Z��~޼y���НƏ������~���!�߿D��]�ԉ�        ��pL|�<��Hi��H�/����X��� O�����d)6��]����y^��9�G��F�*��*�CU�Q����eyi���h����*\�V�/X�@'�p��6����h�رB��v��˅ܷn��b�������L9��C���k׏�Q��c����r�ۏݺu�ܢ����us�����W^���/��R���?.%CC�~R@W���Rp��Z�/�v;N�p{l���&�3��k�iԨQ�6m���d-Z��j+����5�+�T�(�      @ċ��g��g-O�����v�e	c<�$��O	��ɓ�t�.�o�����46(��t0/X�a��r�._�,SXZ,�~@?G���gH�<#F�3t�44x}�pwcg:��o�z[�VI�En�(t=_����N �
��Dy����vkќ3g�pt�6j��ܻ����q�����۷�1��r�#�*69C��/Е�w�u0��k�
��s�=8p�pl,�`ai�466j�ܹ-n�������_n�I6_>~��҆���t��ok��P��v�ĉ�t��6�322TUU��˗k�������]�
�{�K����j���RB�       zYR�bF������RL��Kϐ�e\�"��~�+�uy����s��)PR$�? ���'���1J���g�dŌ+�� Oz�"�'>^��G8�*{�����
��J~�  R����r~��V�[k�I'�$�������{�(�������j׮]�m����?�����J���W�}���%}GCQ�v>x���-5:�p{Z�~�RRR�����UZZZ�m˖-s!�W^y��ƀ?8_^�i_�S��1W�-�y۴���Pv��I�t�g�n���1Uvv��l٢ŋ�n@w����w��B���f�5��׎|D��{]�Ii����w�l�       �Oxe�<�g�����Qc�9�5�Gk�w��Sf��XW�@���y������V�2]�1������L;N1Sg�3nbD��t�{�:q�d#��^����f�o^~ �T "AM�Z���U�K���Z��w��Ѯ��\MMM���Q�6r���;���~Wyyy�m�7�k�.��o����l��X~@��"%�>N�X�}�kp��5U��f���~���ۻ���w����B��|>�r��[~ժU-��|��K5��o)q�d�oU�K�)i��$��͓;���5ea�O�:U��~��wD\\����zKIIIZ�`A��h���ǻ3=��C�L"���yW;���~�_�㫯RCa��W|:g3       �7y���q�a��c���>���䔃A���)K��́�|�'l;�)��wq�kD1�:n��	')���fJ��,����^pc�����߷ǽ0������ ��4���66�,Y�H�kѵ �i��&t���T.��{qq�aۚ*����j�WW�Hx��5�g�W�݂��Y��f�뮇�t��GJNNvg2d��56n�H���***���@�u�]�B�֐$��|9�ko*.u��U����y�K܇%9J9�f�(fM�;�L��;�n��K0�B�����&O����jӦMӭ�ު_��n�Us��Wj��k­��ؿǎe����p4��W\�@�z      �O�����~��ZC{_)�m/O�p7��+����_�@n��hB��/!�5�ǜ�P1s�3�v��_�c���ƹ���kx�����Q`�w t'c�v>t�k��Np!8ky�����{WVV�A��9(ל}��w�;���k~n�6g�v��c��g剉Uw��W��p�C�X�m\m�bS2��痷�r�-nOHHЧ?�i�3F�:������g��,�8}��v�k��n�IUUUڱ�e������5�vϯM��r�;	��M���.D��������v��ѣu�Yg�
w�/����H�v��ܹs9{�ܜ9st�UW��'�l������z�_pO��~���vF�@��ƒ�=�       t%+ʍ9i�bf�(όYR,q��dR��%Rp
�������q������Fd�����*��[�y�i��w��X�\!U�˿a�|kޔl%VS� ���y���Yvۄ	\k���-Z�Z�C�����]�V�s������o�]>���^�a�*6��ܧ��1���-_ۚ�-ps�0�=9������ڼ�(\�c��u��-(|�7hҤIBױ�5�������k������;�����=����^��?���s����|�j(�v��#YCql�@��'	�%��U���a�>\�{�bc�v���Z�}����5���,�D�:�3TRR�W^y�Ŷܧ���qs�>si�|mS�
v��#y��h\m��/       ���+愹���bfϕ���f�X����n���
��F�w�)���4��9��;�bN]*�����!�&�Bs�Ynت+��U�o\�^� �X���JV�>�6[���]Zx����i�2�s�NM�L�bO�2e�n��F=��-���/|O&/Ҡ�˺��j(�sX����F5��)a�(!�T�|[9��\�m�]vY�B�h��{�r֋?~|�?'99مܿ��o�����v;VH��@�~L]"87�A�[�%�ƒ}J>E�U[^��g�v�C�w�y���_e%&&��z�j��fϞ-��,[�Lڰa�a�|^w�����V�C't���V���vkkoMCq�RƤ�x      @d���)3sʙ�]t���*t��8�7[
��koV`�փ����vGd ��^�I���OWL���3u&���|���
�T+��-�W�&�\H :�z�*�>uo�mIII��:5��7Z�b��N���={���g���7�|8p@/�������ٿ��5n&fM<���5w��Xw�}���I3qi�,tᵀ��Ŷ�O>م6ѵrrr\@�g��s�����<ؽ����o�����2y�,%��yL�F�Zk������>���B�4h
����ɵa������w��`g������5}�t�3F���c��o�Y���3^X}��4�ko*&!�ؿ�-�)?�������kr��)       �j�y�bN>C1���!��}���T���ߢ���{��~�e��B���3a�b����%gJ��z���{N?G1�a��R���)PR$ h���|����.q$o�r�-1bD�ϝ:u�k/�aaS���u����܃.��R�����w�=�v_m�v>t��0�1���~��=\�/k&n*�U�0����=��z�Ks[l��|�������YL�Av�c1q�D]��z���[l��W����o�Qlrz����X���]�L��X�O���X�\����r��G��v���w�ys,l�F~~�v�ء��X�	t�-Ұ3^���������V��=�}�.M��c�����J_CM�?�����IO|�,"A�tfu�v&��,6^@�<V9��T   @vrM�6'Pi\��h�|_wFU�2)���s���!���8^q���6ֿ#߫/*@�.zw��־�TŜ{�<c�dp�b/�B�-S`�F�����[R;Cv ���X��8�e˖���o��ǎ��;w*#�F�Ϊ��U]]������g�6n��Fr��{s�{�k���Ѹ��;�@�摼����8*���U�iy��-�i��,���UTT�kLUTT��3�<��Y�h�;���/��b[}�6�}�vM��w�_ou��s�Ӧ�C��oj�(>c�����+���z�mK�.UVV�z�-ȴ�$��m��Ŋ���Y�p��[oՃ>(���9���Ǖ>�le�|m�������-�x��-��$��>/o-٫_f�#䎨b��[J�jpY   }Q�������#����n��y��a[{��3o���N#�'>^���(&8��_��^����
TV�	��v1�&*悏ʳ�47�!��ì9��@q�|/�]��/Ku����_|@�v����{�G���������w-��8k}��$���IJJҧ>�)}�[�R}}�a�
W�Li3����k���v�����w��^D��8�UoSy�V��-y�m�i���B׳�������t��.�L999ڲeK�m%���9�?��8��;��fb�tɎ)��N�mv\9~�xE�Т�7�xCÇ׌3tִi�����׿�ض��;4`��J:�C�i-�Me\X�3��劫�RlR���B�цp;   p8B�6��#\r��P�y�ȓ9T�p�G)��O(���x��������N��m<ӎs��1s���B�!Y���-�������ۋRI� �ڪs��r�m֮y��׷�~,H��E�ĂV�����j��X�����}����<�IFJ<�����v���T�B�qiC��c���_ܨ@���\y啚2e���*++���"�_MM��,Y�e�gA��o�Y���7U^^�b��7Ӧ.Qqm�O���ٻ���{}��93��l$a��}������ui]��.�����ڽ^[�{�����zۿ^���+Tda�({�@Ⱦg��?�(���s&3�<���t�7v2Lf��������#�@޶S�=��7DBv.(�Zj�]�"mi)������}Cv�y��1s�Lcm@��>������ �ۛ��?���G���0G�8_�^�N�6œ#X�A֒���u{�,C��n'""""��!w���.e`Գ·z�砤�������EP�C��C���_��Sŀ;���k�B�~ʨ� HJ��K�:�BW������w�șB�6����F�;����n��座�Ν�����S��}�aÆu�'󔔔]�W�X�e<�ވ=�|	�z��}���U�V��k��;5K��*(������V���&w_��SS�fXoȎr�I��w�q�x�	�]�<$���7_��o-է�ȿW�o��"}!s�'}(w��%R� ]����̌�y2;;�'˚@ִ�:����x�سg����v�A��~���?v��bGo�N��!o��w�d��J��S�c��������r�X�p{lR�N��ˡ�9P��\���2i�>���]F�0��=  �Yp's��PK�u�uP��{�-�c�ig��e�h�w���e�_FgUEğ]{�������I�N��wtt��F�U�2e
(z��s�NTWWwo��6j�=��o�?i!xk���]�����7�'�k�XҰ��.>l|�����@����4����>+,,��Ǎ�K.����j��Z>z�^������I��W���"EE��H2�V�/�W�6.��E���s��v�׭[g��9s�@UYpF=';�ȎO>�$B�P��|��Șy>R'̍������5-3����=` wc$�1�N���v""""��aȝb��G����j�|��hS��qP�z��7"���Cp�ۀIM���p�S��P�K��''e�H�3(�g���/ڰ���Ȏ�DѺc/�uğ͚5��vZ��wڴiX�x�ѩ������8q���w��q뭷�'?�	�*�+�t?ҧ-D��	���5�B�gM1���ܩ������Rp������K��[n�))) kHȴ7;���x��-���?�|���G}����ξ�#��k��ѵ=��l�m�#��j"�����P����g�����B<9ֽ�_��rss1i�$����eG�7�|�˸�`���[����P=���R��Xe����{�]/��Ad5��)�0�NDDDD�;�S�a�=�(#s��z�D�ח�z�U�����B�6i!ga���X����g�ݑ�:�j~BkW ������e��b����
D����v�݈�O����J��H:B�Y����E��.��R���+]�C�6�~�6L�濌�e����ܮYX�,��o�FB&�e�`ߟ�G��.l\�k�m�:��6d'����|�uo?�Xa��?����.?�>}}�EL{lőB��Y&�7�R�D�c�3_2�Ow7~�xL�<�J
6����d�̞=;���dM)�@{���2.�g|�Gy�w��e�)�v�Zz{|�\�N��'q�H@�cȝb��DDDDD}Ð;�
��c�2b\��j�FƐ�G<�H����!����`)���'�S�)S��}�PFskwb�9�A-�gl/��?Akj�Kի��Hn��&#�~*�����S�'�.�dg����ƍ�s��.�-ۖ�v�sH�;���ܖ@s<�C�Ž�5mzu+�7l|����K@֑��{���=*�^	�J1��~������\�C�?�ϗ��iֿ�hob�~V���\�fظ<�8��;)��Cٵ������GB?أ��B�/~�����o�q�������!i�Dt�e�ܭ&�#�R�.�5�Sc��������0�N������jtlw�s���!I���| ����4B۶��7�~�����7A���ۆP8}a�:��sNG��/!�ƫ��ſ��M8���F��駟�3f��{�̙���r$%%�zo��X�j-Z�	��x�aa$	�^�Z���P��x�.����d� ����{��;l\UU�|���xֱ�toommEzz:�g��}~~~�~_AA��-^
����e�]�=���֜<�ӆD��!q�xP�;���/����t����'%�.�ʕ+����u�NF�~/�����k]Ƶ` #6�S������o:��˃� EC��_n'""""2C��_n�.7\΁���4~VG�1����OZ���~�D�I �?��%&�u��p]z5��tr�T�]{\g�����5NLD�4����K�t�����M�U���p��49�����9r$(z$�t�E��W_5������wމA�!ݷ�O֟JZTn���0�C��"�_T����;���9��3d�͛73��KMMM�<M�]w>��c����;��ƍCcc#~��_b�ߏ���7��k��0 ]^�6�Ua�yyy1Z������ŋ1a���$�a�TVV�K�ǿ�ۿa��"p����-*�%�!�R�.�U�S�1�NDDDDd.��)�n���Yp�x��� �,��$��B��|�/@g�N�)2:)u�p�p��Y �a#���w��{���V{D�V����ޏ�3	ZH�p3cٲe��� �����֭[p��w�ѕX��n���9	����@tB��tq8]����O��:�\r	�Zuuu<w��L�2%�W��W^y%>���v�m�%Hؽd��-�W ubiTn��� ��G��
tx�o���[RR����DMMv��ats��D��dgYK���?6���hԨQ��:���i�m�N�$��S�����*��{��_�un'""""�C�-����C���P�@�+		p]r%��g"�ǧZ��N��Sdك����F�ѩ�ǐ2uB/>��;� B!Q|y۰�/G�Yaa!f͚e��@�8��+�Mvv���xƌ����x�	�qW�L?���C�D�(]�=CEEϾ���` l��k�������}�v��{���EE���W\aI��]x�X�����נ��oU]���P=I�(�B��?wF�'O?�t���#k]	�oٲ>����<GP�ѣG�[n���ӻ�^���srP��6*������ w*_Pte}�trgȝ��p;��r'�1�ޏT������/ 	� �+%k�_�&B�Vi�[���)���a�JQ�Zx>\�}H�v�d%)��z��<��=;AD���o?���@ظ�,���Z�~�I��x�b#�C}#������ѝ������S��X%h{�С.?Ow0;Q��Q�=���IQѴ�u4mz+l\�yyy k�ݻ��^�͍�6�rN�s�t$���4v�W�*!��/����}�s���m�/��ef4Ծ�<Z���0aF��IHH0�+V��̙3At��J�CYY�Qq���m8�8�:�/���1��3�N��X���\��b1���v""""��`ȝ��p{�Qr��}�P&L�Y�¹P��@��|��l�K]0�N�P����֯@��V�ʘ��|�I_������&o�nT��dğ]|��HOO���Kw�;v��eI�ZS���5p�@L�2���رc��s\�V�jT�ةE�v���p�-ľ�|#l\���_~9�Z���7���s����N,�$�qRt�qRR�ବ�������cيg�y>\�֮5D����#��3��B�Nx�Ѱq�'�Ν'KMM5��󎱞���9��d ��cE[cƌ����?�4��a����� �!��@����4Eۑ�{%�eȝL�p;Qt1�Nfc�����p]x\W~A��������ۡ�9�g	��>	�8dtm7���fi�"Kɢ�+��*B�~m�Q����7�0RwÇǙg�i���~�!�@2MMM��� YCh?���G�6
4��
�P�\��;�\��o��	���[��_�C��-a�R����VEE����СC�����'��*"A�Ç�܏w��/������k�mӴ-5��N�����.��H���Xу�eee����3ϛ7���I��I�12_��@���]�[�!�Nmæ�d4�vD����p�~3�!w2	��DDDDD��!w2���C=���e$w�%�)�����_"���F�M_��pw��p�q�6&�&ٶ���/|�O��n/BC$�Y��ň?�ꪫ�jV�3g֬YÀOIWԵk�����KB�'O6�h�6�����w��Ԁ��PժD�f��\̀�Ť���+���K�}ѢE k��԰���$$�`����.EQ�"��#GF����7n�Q�v<�C'�Kq��
����Ns<Ì�o2_�����Ӱqy�N�6�)Y_Ȏ�����������O�	&�fw2Onذ!l�_Y�����+�wE�&"��y<�N��$����T1�NDDDDԿr�S�p{?P�λ굷@acB����o�Z�~�shu �b���Ԣyp�z/�f���D� ��R���OHO�D#�����̜9yyyQ����HII�Ɗ�>��؞={0f��9"u��N�Ir�wmjA?�%��˭c����;�H֩~�)�k��?���AE���͛p�%�â��Xd������H��������^��x�y��aXM��@{#�)�	�
U�|��w'��oG���l\.[�#F���)S@�$ρ����IKK3v�����2.ϫiI�xo`
j���Z$d�Qaȝ���v""""����;�����s)(�g���_!��S��W����'JL����:�|�e�,���bD��24��-l\�،���,Y���Q���mǎ��dȐ!�8qb�y'
m�r7bx�������h6�ݍ5
EE|��j҉�;|�Nkk+�ϟo��P�re'���sT���2NI�����d���-5�[�[����6l\Χ\�|6y.������F~~>�
�)�B 	�y���Յ���Y�3&��WV�F4�J�YCaq
��ܩ�n'""""�-�So1�}jq鑆�����%�Ք�xx�%�#�³����8����߂�3D��8!=�(��z�?���D}G���wL�;w��A�?HWC�X(]���233�~�z̞=�7h;vl���B��P��/{�#D�N�[�D��>l��+��|���=
ҧdW�w�.�&L��s�D݉/��|<��s|�7a5�xa����:Ⱥ�zN��v�ލm۶a޼yF0��[VV&O���9Y����z���.�Rl75�����]�����l�'�ܩ�2n'""""�I�SO1�e���o���+d�r���}<��!��@�>r�D�]�]_���
�X�:�(�s�Տ��Q���X��Mo��K�⢋.B���Ν;������������.}�7�5������뻆�sZ12%�mև�D�F��5b�v�Z-��Vgg'�^�����в�w�\�����?Rwb9�OM�CU�^$��k���2��� j�{.l\v���.����1�5k�k���bS�)yH�do��䠺��P��x���8c�yxe��w!s%וr��b����"+�p;Q,bȝ>��Q���=߀:}�b��;����>�P�J�30���bTW���IZ��(֩S����_ �ԏ�Q"��C�I���U����k%�}�����+WK까�#�,���=ztX�]0/e?��-� ]�D2W�ۿ2���.��b��֭[��$v����o�}&���M����u:��2~�E≗����|V��#!k�����?��ؽ��� �wǞg�/6
C����I�v���R�0dȐ�yR��&�F��{�ۆ��jB2��C�t"������4���Dn�.e�����AC@����?^F���nMa�~p�;yR�� �BnN�E�׷�/����Y����h(-l\���{��o��50�~
侓�}�8�ȑ#��5555b�Q��J���VX.�ي�����`3�|�8�Ɠa��Ǐg�0
���qP���g϶��"�M	n��c݉ú�h¡��p�Y�ƪ ��wJ&��Z�P��ٰ��Ç�{�Idm���dݥ43���X&�A)�<�B���\>|8��{G�F,�r.^^�� �q� �(0�N�1�NDDDD_��ܟ����	�G����N	��(nH��K���3�_�Z[B�o8;٘2l$�=e��#���������iV]YH�lB�����X0�|���{HKK������q�9�NL�:&M�dj!@�.�� �Takt�i��z��\�����"vo���KA֓��+�\[[��#����G�G�e^�Q��ҝXB�ǻ����7_A�Yw�j2W2�~�����U�;�
-�J��l���0
A�͛g�c(���&L�j�'��loĴ�f,K���vX-�ϕ	�#�������ۉ����Ⓞ�o����Y��;��Q����N��.Q�RgA����;Ъ�쉟|ٔ:q*\<%�� QPϽ�a#x�G@g��\��è��Oa�ҍ����C��P�������	�	A�ر��Pd�4�˽t�B����.��N���?|�N��O����ۿ
7n�L���t�nmm5=�mg��~�̙�_�̓f�ۏ�.�ҝ�{�\�v��ڡ$���MF���[%}%��Ë6.ǭx�Б"F9�/_n�JGw�R�#��(&��y�=�.:*7a΄yx�|���v�����X��;1�NDDDD�2�~������Q����!��K@��#�������Ul�?��!�d>�w}M>��]�3�������w��:�y$���cРA�%yyyX�x�Ԧޓp�޽{�0�]$����1b�Q�a&	#u�����s��2��B�:T�RA}״�MtTm��ѱy�f��{������k���Z��@
x̔��l�=jjj���u�<<��Ȝs5�$��@[=<���gNQ���F7��f̘�ֱ]��,Yb3�2Կ�0W�v���Yd��������?ڇ%z����j�ŝw�5�;��DDDDD����s1�=Jf6�_��1�Ad�ip=��w?Gh� {a��f\���o�6� �%w,<���߅�w���I���e����XlN�6���7=���	���%%�Ȏ������cǎ5�z�(c��hoo�2>3���=�F��	����~6&��g͚����e������;�޽ےвu�˜����^)�RQ`�k�`+���߄�I����fy��<)��?��X�0��ٳ�(�1�̓��"T]����v�!X-�� ʵ|N&�-�ܝ��v"""""{a��yn�e�h��.��� �����#8|$���/�>p�U���/C=�ٙ�5�o��'�V�Dtj�^���`ظ�$8���vEE�:��������� I᪪�0|�p#�g��#Gb���]Ɣ�LJj�F� X-�ֈ��i��΃�i�[a�-�Q�c���{���EEE�]��J!���]U�+|zz:������Μ��v�F��y�R��-���Oz�e�2t��6>u�T��|�)��$]��l9�y޼y<W���g����k�u�� �+e'��y���(ۡENVҴ��p๙bC���p;�=1���G�:}��Hb>�lLQ��z -�?��@�0ځ��o���@�JJ*<����!B�@D}W����،es��Eyy9�}$��W�Z����:{����ɓM��!C���@��:ljN�>��#�m��.�}r����4W�1)�(--YO:�����ѣG[�;v�څ��(&�H�݇~�eL��K��8�.�����2OF`���z�X�޲eˌ.�3g�E߾}�0t�P$&&�v�R�+]�����Ho߇�!�[���p��Ő��1�NDDDDdo����ѣ�*�����\"gp�{1��T~�$
�������������$$���#��OZ������;ѼuIظ�pg̘�X&mv�<5r:tÆ�;|��JKK3�:�1+�&��y��@Fg�Ş� �&A��{M�9׭�sظt�e���������T__���B�O{{;���M?�dgg�����O�<�etb_[=�)Y�RP�+p�C��-l\v/���Կ����ǒ%K0m�4c��)�����ĉM����EF�';��a���p�7I�P���bC���p;�30�n_�G�R0�{�]>d����g���/���/�㘢�|��IHNFD�$�>��ӿ@��% �ީY�LX7bq�駛މ�
,�n�M��[�C7m�Ā�IH)//���@Y���tۜ�t{0V3��9��i,��ڰ���Yd���KR�-2WJ��k9?I���u�����@���a�`g����0\�վ��q�u���E���9�u�Vc)x��b ٝ¬�8)�������˸��&��!#%	Mm����a�-p� Q�b��~n'""""r�����葀����/\ r"�Ժ��_|��xŀ{�JL2�W+�g���T�;�G )�w�"�	#Ծ�|ظ��%8$H']A[ZZ@}#r�mۆ�S���I䶶6����v�j�.�MMM]�'�vD'��#�m��h޿�	$��ݘ1c���b��������f,X� j�����^H��Lp߻w/����!�K�1���3�;���#��[�B�XBB�1WRl��������r���ĸ$k�\&E�&L0�:e��p��a�ةX�e?�lod��bC���p;�31�n�G�����F���ɔ�B�z�':;@��x���?�e�t�p���;����	"�l-ۖ��x0l|�̙HKKC��4i�y�dee������FwU�/n#ڷo�L�b�uJ�{�=�|�F���v43����Ch�����.�z7n4:S�IG�h��2WJ'a3��{<�K��7{�(���sf�J��\��rt��6>n�8#LM��X'�w�}�(e�}�I���\���R��������.�ޚ�(,��w��R$d��>W�ce���?�ۉ������!���p{���.<n��QQ�P�N��k�!��G�x�O��σ�0�=��Qw��яF��4�������
���n<���ʥ~d�Ǡ��r�%���떻�y�}�Dtr�+�q���NC��={6v��� UIg�U�V�������"I`�,ҁxǎ�]��kQ�5$��8�3u��-�2������"��d�3wPp	9Ο??꿷��uuu��f&)�p/,,��}���{g�����=P���Ǐ�}���C�F���b�F(2���;ִ딿W�����3��
#�Ӱ��V2v�u@MHQ�c�=~1�NDDDDD�!���p{���/�����Ftȇ��'�ŧ�B�~�i�f�������B�c�V��(ҥJr���i�м0Ed�����O>���&������e�l�i$��]?���.�أ�H��'�=>�ooii�i{Slܸq��������c��;���˙���	�T�;�G��Eh�
QdBh(�kظtȝ:u*⍄�6oތ��tP�HgG	��S��hڿ��[�Y���t%>|�p���P��@Ms'���m�ŗ=Q���ac��ERR�Z�ׯg���\.W�|UVV�p���t:�_�}2&ߏ֪Ф� źN�Z(����$�OJ�;ԯ�a�2G�b�x";"�޽�XWK��s֐ݓF�e�Ra�����ڽ�;�?���v41�Nq�!���p;�!���p{��sN��������ZQ�͚�}|,O���n}|oAAA�Y�dŊ�			�����8�G�y"�T���B��o �ԏ�P�j����נ��Y@?��O +���妖��.\hm����|I�ɱ���V�Z5��r��o�E�m�ʣ@�������|�M�@D�6��@k]ظt#V���μy�v�ZS�l;��֬Y�E���I}���F�n�H����`G3&%7����7�$ %�˝j}��x�ك����KJJ@��z�q{N�/������@[[���i�uꯍ��|UUU��¼	���H�͇�d��O�y�����7���8$2RX�z�j$''����x�yd��dmi)��.����]�}u��/9o�W���V2v��xq,��Lv.Zr�i�Q$���ۣG�]��_g����ӏ��Q&���MG�~�;ڀ�����ҥK������/g�k�~�*�2����Z4�@�7�!ۮ�b��@Q��P���>�ˉg�~|�O�k
���Ν[�_�s�0�Y�&G��t��_��_N ���ml+��ɣ�*������eSH�%^I@�]&O�t�߷orrr@]I �СC����Ǥs����WSR[��:�ŀ{�4�}Y ]Ƥ�fڴi k�[��WR��|���B	m�pR�=��������>`u�������a�+�%�N�+55ո\�x1&N��1cƀ�#����\ӊd��p�](\��0zp:vW7�J!o����M�(~H����}x&+�!��p;�C���Q�ς����{woIW��C����}PRR�1�h��uG�ƍS�~�td�/��~H���a��g���"��_�e(�pf���o�z�٠٫o�'�7𯼼�Vĩ�'�?=$�3A�w]��\/�/�ԇ��9��Dx|�Ǿ�@%��	4m|#l\��73��
�z�S�I�Պ�
�O�� �\Ovv�q���5ap�(n��&/���le�={��ᖬ#�m����&؝����������f����Ҍb����O��52T�f-�O��u#	�:�P��pd��������Æ���dee�����Qkv�S�|>c�����zdm�u{#�{x7��,�<�.�WB��tœA/C�1��v"""""�	��c��ѣ����<|o�������
��(..ޅ8���߆#������Ӓ������%[���NJ]x\���ߟ@�����8��s��*�II\�G/J�v[������ů�X�bErbb�T=\���.�/S@����������D�n_�@k�󡨨ȴ�n������{a��[����6mڄ�3g��2;�$p��cBz ��`�P�M?��wB��j}�\6^PP ����둒��mo���!##���/�̽����26s�,>X������5��s���.��~ظ˩��6�o)��m۶���g�q�Lp��A�֕���ݘ���. }�1�x�ܠ ����`g��$�~a�a���X2�����^hpy�nj6l��H���@~��o�؈_Q�N� x�"fd�X�V���32�����u,��	��sZj���g6��v& ���h�GV�k➐��E���| w-�%%�z��v�)��p?� ��QOB��/�4�%�����N;͖]����^=z`͚5y��\�7�ߎE����A��C�_o�b?��a��B��t(�&���'�����ٳW�5�~"���Ҿ��r���}E�/>�����/ ����Ap����v���6�q<??v0a�,^���%O����s2�K��"	�m@_�ݪ�7)�+`���Dr�����{{�A�+��ɓA�jii1�z�32�L�>���/���g��?����{����h\�����+E&�@9�/_n� �'Q�544III�\��Q��e����LÁ�fX)�ϕ�K0�C{��׌��)Uƒ*OR��vg3;hry�,�UƜ���TU�ik ���۟��]�,r�5���rY�A�yr���?3�a��b�>}=qK�>$2����%g�}M��qTL�(1�������r�t�u]L9�IFjЏ	�6�E�����c@� PY�I��������]C�'SRR�U�تi�w���J�ݯ�~ ۍ��;8|�-@��ɥ��̅랇 ��b�>�>�v�_8�݆��'��˱~����`�K��7��P�A7�<����B|#���q�?��$D8f�؅tW�裏�����BK+W��駟��� ��?�������`�	����nmaV��`����6�WjO�:n�g�͛73��Kh:4v��V�x!�&	�z��v|����X�&�mE�P�Zؘ��F��/y>�w�y�8/���wRd��0)ڵ+|G]_m%&o}�]B���G$����\��c��M�������r?		�?�p{L�$�k�Ì�r?1��c[��Bo��O����V�0 ���'r?9��cW�ˍg�G3��$������p{�����s�9��q?&w�=vө*<w��q�.�����<[XX����?�c�ҥ����]��ݮi�"����9�}߷���C�*w�b�1H��|�q %d����P�����[@'4{������[�n}����
�~{P��m�t��b�n���"����CǾ�a�ҽ]�ћWYYYF����������� uU]]mjgZy�v��aL�dl�8�.�)2�x�R�nظt�&k>|��݀zF�4L�4	�FB�f܅̗�����e����	�d��W��Z(���]�j�F\W��ɬB0�mǞ�۶mÜ9sX���֕f��"���dtttt��Ub���Xf�ir>
z��JJQ<`�=�1�~r��>��O��������1�r?9��cC�'�p{���˟�b����R0t��ie��(��rQQ��%|�eee3���~�>���p��p?�(��>����>�0�k�*�އ���ҙ�9����Y�f �X^^������I�4��^��\?��p�w)�}{Z����is����3`7���3�����X�/�8`�ڵ8��A]��Ԙp��a�r���d�R=��An�ŗݵ�Z�`{S�1	��q��%;v�`���dg���"��]�@�(�2�̗����3�z�j��8V�Цt&fh����F1b�9TU5��6m2��5����zE�r��Ԭs�̓����fO�b@R�;��0<Ā;�	���C�1�?r�����{8���C�1�?r���������\�^uх 9�)K��_��+�}&���q�Ƈ}>ߗ����{Go����F��o � (v0�c\7�	e�48\��i?KHH�����6�)�OJ����k׮����c�}+AwǾZu�t�{wA۵DNӲmYؘ�R&O�����t����e_I��]�va�8nmv<	���!%Ŝ��:`� ��w��~|�O~z�ǰ+��dv\�y뒰1	m�;�����ˀ{/��� I(���C�5�:�!�&r����{���e]�]0�����Ç��G:��w�}�fAX/�N>fܫ�����1fH:>����B�m���4���C�]1�r����Đ��n�O�w�p{�aȽ+���C��Q'N�����pr2Y�o�NI~~�a�Ɑ[�>���!!���GJ�0�x���(v0�C��΂��`-��k��Qqqq�T�}*R_)AwEQ���Ġ���}߆���Bk�Ì������1	/'%%��fϞ�%K�0,�GR��s�N�;�ҧ$�dV�]�c�{���Q��CP�`�=Fh��0�[��M�2d��5�s�%����J�J3��Z�L���񆹚`��>�e����w��d�0l�0�s�<.]�e�����CH1����MYo��/k��E����;8���;���n�_��p{�b�����C���;�܏`�=~1�~���!w���އ�s����,�4�EEE� S������[�n�ώ��������]�g���Ν�b�:n"ܷ����'���n�gϞ���Ѡ���֭����?׿�����!�G vw&���솯�2l|�ԩ��I�&�СCFЃz/++�ׯGAA�S555=z�i�'���6-���B�ş{2�N�Y��W���q��XRQQ���^�.ɱL��@ n�l������f`�>g���*RD���_�ްqY7صp�zG�sٕc˖-(--5v��Ȥ ���ٔ"/)JMM5����h8��3N��B�����X�p{�szȝ������;�����;������;�����!w���C�@����w(Y�}㖇B�JJJւ,u4���+V<����-������u��e��섶w��1�RR��t�v���/�-**������U����[�N:��L?�K��u�,����?�7���eۻ��ޑ8''۷ogW�S���jo�0�#:::���f��">>�F�uXg�r=��f���k���9,E2'NYC:}Kgn�9	/.X� �L����z2Ĵ�T!k���nDZ�"X�Hh3 �ŷPD�K#��1D�Hq�������9s����<h��9�v�K�N�ǋԤ�vZ��O������é!w���é!w���ŉ!w���ũ!w���é!w���!��q]�%�S�Áh��͢��?*��������^�xp�����?п�
N�� �����-͠��Og��~�v��0ؼ����6UU�RPP��o�. ^ڸq��~�������p��ˡ~���� ������x<3f쮰�[�nEb�c�7S���`�ʕ1��6	"���r] �����76կ��=FH�*�e��ͮZw��F���ڼy3�$ss<Ee�43�.����:n&�~��2�+��Bvwp%�q*Z?^q|��� �.99ٸ\�lF�e�D]�\9~�xS��D�S�A�������J�\ɀ;�����i!w����i!w����I!w����i!w����i!w���!��Q���uޥp�NEQ~��zZZZ��7�g�ޮ_\�nݺ�4M����c��W����x�q���?L��39	�3� ~�x2##�;'N�bB~~��o}T?!=����ֿ^'��d��nh�� ������F�mk�N�!��ޓ‚�<tDCC�iw���pO� #5�-־n���P\��#�"�ǎ�F[[�'�G��Yc�������F��b�hr=2_655u����Q�����#�v�����fذa :Y�Kg�7�|�(@��S�[�Y��0��T���)�����(V0�n_N	�3�n_�B�r9��!w����	!w���퓐{�~$���+����)!w���!��Q��}�W�0(�r[aa�6P���o-]�4?55�a������#ެP�@]t!B��	�?�O��0ed.\��Y����b�~Bڡiڢ�����˟�C�Op���u����QV\�mI�΃���7NQZZ�w�}���H��oذ�s舖��A�\.S�O����]�-5�9��{��5��c�v�c��:eeeFWn�9�w�@M�I	�K(�,��p��΀�����&!�Ⱥ�"l\:sK�={�#�H�B��;w�Ķm�0w�\$$8�}��$Af�e�.�c]�@K-F�Z�M�s%������!w���O>����N�v�3��r����mrg�����>W�5��p���=��p��1��T�;�R��|%�5�ǣ����R��c����ceee/���G	�}�m��ھ=����ۑ��W�8�<����]�~v��W��ա��y��i������tt_ �Sg�)���쨽r�o�9)��/ ���Nv���L|��ǘ4�1�N��t$�.�r��!R�3����t/�.O�D:��x��}a�cƌ�����V$�r+**B<�0���H�jcǌƇ5��4|
�����{7@��eg Y[ʱq�F��0E&!l9V�Xa��KJ�>�I�sfĈ�\�����ꑓ���.R
YW�/;���~�p�s������d��;���aא;��β�h'w;��nw���nw���nw��O�u��N��X
�n*))��yEEE�_|������CӴ��!�L2�w=��w�������~"�ە�1p�
EQn(,,\�+�	�R?-\�nݽ��?�ͷQ���7A��"�i߳>���yyyX�x�i�d�������Ä	��:D2��$�.�_��]Ƈ��K���7C��j۹&l,))	Æ�O_g]f���~��'ҕX�{�%R��������vk�~ɉ�ݑ_�K�����|��e͚5���"9V�"ktYc�qpA�̕f�⒚����� \^}횚��f�B�R
x�z��\E��p���mrg��y�rg�ݙ�rg�ݙ�rg��y�rg��yr���U_��5M���ݻg���r�������C���׶���/ ���E��@�>��?�S�w�������g١�vsj͚5+TU��Dؔ"W_���Ǌ+����ac&qb�[B��f��8p ֮]�9s��"I�}��ں�K��?K6�BV	���#��m�n�,�0_0D @bb"�g$�>kV�u�b ���>T��tBB|�O?���3�u+�$��hA?�����=�yn�~�騭�ņ�C:y|H [v�n��t9'�:Ќ�"���C2����;��nw.���nw.���nw6;��nw6���nw.���nw.�܏#٥�<l\��6MӮ/..^�[e[�n-���|J�{~6����6�Ch�FPt1�m	�p��o�۩(�]��� �BII���˗&%%I)ҕ�)�UA��j_~Dv�����T�����QQQ���tP�H������8�t���FH׬�		4u�'ڐ����v�B�؄�O�|ð�j[��ȑ#A�+//7%��$2?�c�Sv�hii1��+�����.c�FX]�������6&E@'�+���>�XUUU!##D���(;;۶m3�Ws�΅��-�x���Ќ��f�F�R<�rb�6��)�C��S���n'�!w��I�{ȝ�v���;��Đ��˯�2*6�7������	�����	��u���KӴ����$QU�n��7���=���(���ʐa����\QXX�	d+��vZ�~"�Z?!ݫ�l:�.��������]t�(l�ɁM�>.�J��J�'���ի�p�B8�t$���Ya�H��`{3���4�.$��&�9�QU6&�1d>y�ب�$$>c��+��2_v�g�;Qk��\�T8�~��<�=lxȐ!�D�2e
&M����2��>�at"�C���������|8�̕f��.�9)]�lo��l�{Z �>D���p;�!w���x�3�Nǋǐ;��t�x�3�N�H���A�񥺽G��n�c��ܯ���)^�ܕܱp]t9lLN��*,,���(�m_N�B����f͚�����;6����|����e@5V���u�Ű+�����~�̙�������Sk׮�P�����ٰ���F�_�$�❿����q�vp�y�i� �&��C�0l����z�̀{�����&NO��jX�"9=அX%�6mb���P\\�x�}w�S� hhV:*���NɂU���5V!�sNO��CwII	:::�b99
ُt!���;�cH�����̜+������u`��	��'�jZ���4�>�p;uo!w�۩�x�3�N��Sȝ�v�����[��D<��n��ZT7~�?!w�۩;	����������� �ms��quQQ�R�m���lX�bEqBB�d
υ�ο���A۵��c���m����3���_^�pa d{�����ѿ��~L��+F	�����P�E��;K�e˖1`�GR  U��"%%E���tY���t%vz��[[��7���ǹ�jjj����3�[�t��gf�#u��b��,��nN�y���]W����3�DUU>��Cdf2H@'���eVn߾�X�G*p�)��;T�;��YX����\p�������s%E��t"�rg��N$^B�����Cȝ�v:�JOr\��n����;��t"N��.���	�����]T\\���JKK�_|��ǎ���(w�nT�۾
����'+�d���(q}�(�FÆ�s��=�$��Q���v�X��4!!�U���a3�knB�|5Pcq�\"�uVG�<N�/�1b���6�Mvv6�lق�ӧ��,��2`��Tc	�+��<�i��;v0��K�����F<koo7���I�E
�:�]���3Vт��aP4xE���H�brlݺ�(|IKKQ$��������KKKM	���'emi�s!�<)��i)�hl�U���EǞ��CV��tB�rg��>K���n����;����rg��>K���n��⤐�2x(\W\;�4m����\AAA�1���jY<�SVV&��'��V���;��.G�A�c�=���z�U��EQn(**z�HRu�t��s�����{%�$1	��D���(�u�6&��۹�aOM�<�/f��Sp��aӺL�+3C�r?&&&���6�7=��bu��fOؘr(���T{����K����wr���Ҭ����BBB|�O?�IMM�ڶV�~8Y�	v2d�)]o^^��Y�z�qN�s!Q$�B۲�GL�2vcm�v4!c@��w-��-�PT��DVa��z*VC��SO�jȝ�v�X�3�N��!w�۩�b5��p;��SB�/�md��FQ��ddd�<q�DvZs�������ʪ�/��[=�]�_�Ъ��>��Q��6(kCI��MӴ��h1��.\���/^;nܸ���~	6��.��_���2�+��ac�B����|�ڵn7�D}!�4W�\����é$����a��A��w�g&	��ﲊtvhS�����4d��{{/544���v �M3�$�y|�]��JN�+�5�#�K1Щ��ܼy���҂�k�_'����T攷�~3g���.�Ȭ݁NT(loBfJ&��Z2_2�NV`��z+�B��So�Zȝ�v�X
�3�N}k!w�۩�b-��p;���C�J��3��9��4M{����.EQ�����BQQ�Kk֬9�����o����u_B�? Y�i.���gA�]�i�B���� �l-�/Nn+++k�'��F\�ߊЖ����m)>����:B[���%��$����P�Hf�#���HKNCS['�������p l�wsUTT0��Kf�c�tp7S��2m��'1����� ��%Һ�����:묳��~c���t22G�ݻ�X�K��Y��d�\)E���m�2V3
�<�j�C1��v�X	�3�N}u,��_�k￐;��t*b!��p;��X	�3�N}+!w�۩�lrw���V}D���WQQ�WE�@�+))yw͚5�TU}S�66��B�>ږ� �0�n%��n��4�'����g��star�ڵk�����PF��u�����⑿)|;��*--��իm����_�`ѢEp���OEBB��!oR�<�܃��j+���6�t"Oc1Q�477c���3�J)���
ZpR�x�D����,y-h��5j�qlܸMMM�v�'{����|�n�:�𥸸ؒ�d��5WJ�I��B�v�'Y��$�'�l�ө��;��t��×d���!w����rg�����!w���T�wȝ�v:Uv����0l$l�'����������eee��_����2��v�����~�w�g_e�h�H�~�����At���1��$���;lB��zW,�_�5�(����1�ٕ����A}������J���|>���poG��A$�w%���ac��&s�_�����+	'څ��H�� ��oIA�#�Suذܭ���o�gW�Xa��#�݉ıb�%K�`ܸq���.����Z �v -3
�w�#�0�Nf鯐;��d��
�3�Nfꏐ;��d��
�3�Nf鯐;��d;�ܕ��p]vl��EEE�����G��u�i��6�䮌̅��<�����QRR��z�H�>���p;��~B��ѐ���y>�.���~�x"]�C��/���=\AA�-[��eI ���±w�;�}�HM�F)���7}�ᝉp7G{{;w�襶�6c�;1�HHع��d}�f,i��h��?�Ec��s�g����:�XF�5~�K' �u���k�.��k�����J���ܥ�{֕2�N�`����;��d�h��n'+D3��p;Y!�!w���l��3�Nf�K�]��� [���p;�Daaᦲ���/��[l���&�V�����p���k�T[<E�����Q�'�����gj��E؀��|�5���㡈���N�cǎ5�SL�Mvv66l؀Y�f�i�mJ�;-�� ��	�G!���>�TĀ�9֮]���TP�ɹȌpc,�Fw)T�5��1Vqj���y]����=d�q��gc�Νسg״tB2�J�]
0e�x��/�٬�{w�
�k܎�L�p;Y%Z!w���*�
�3�NV�Fȝ�v�R�B���U�rg����!weT.\g��P�w�������V���}N�����x'��/��?�7�|���<F(��PϾ6��OD��'��@���F{��o?~|��iW ީ.�������ⅿ�&�8C��I�]:=���<��<�{��`��� �/�.��Dq3)Y��Vb�q�6u�8�[oi��i�=N�>M�OR'��8NdY�Ty�]� (R7��b�w�r���%f@b�w0g��{���� �9������R���ׇp8�4L���mz<����z
��tq):ҟt����I�T�5%'�v�� 2�t%���,�)���p��w�Ε�����1O��1�u�ts�t7j��ѣG����m۶A���͝{�,�<iNz��0�+�d����vr��!w���iN��n�Tp2��p;���!w���iN��n'��r���OK>d�o�����d�@4�`��P(�	��SȀ�~�曐'��>���?8ґ����*2į����D����G_|��O,4c'�o��'`\�"����345�guzt[@�.����7���>7� �����?U�N��|H��A��h�{N���󭱱���ɜ��ϙ���:�&{y�"=�~pd�+���ו�U$��ȺM
Bd�!��L����s�8=t�V�^��˗#��U<9�|����xtD"�gFD��p;��S!w��)U�
�3�N��Dȝ�vJ%�B��S�8rg��REŐ��d9�z��S��ZXX�s����@��`0��B��gͻ������'�;��)�W�l���C��02�a�S__��A4�����mE���j�L��y쓈����
�
"�0h8%��ng�΍$\��Ӄ�����ۣѨ-���Ç���{d$y ����fO^2�fe1�1]�H����T���.�3���R�g�Gᨘ;?���i�t�޻w/���q��I����h*������Dss3�n�jg�#9�a�u����8p7���f��vJ5�C��S��rg��惝!w��i>�rg��R��;��j�C�꽁�
�ܽ�&S��7�����j��:'W
�
�֚w��9�D�{��هw���Ih��4����~D60OF]ǎ��y\I�]�ģTRj�V¸z	D�.����5%FS۾};�=:oIU'AV��|��A�I̦��T��Ttpws���Hbw	�q���'Np.����A"S�l������|nn.bag?�vkhs���ҥ���=�Ξ=��7oZE�D�H�9>N�:e�;w�L��V��J}�eF4b���5��c��f��v�/v��n��bWȝ�v�OV�]��X��Y��n��dWȝ�v�/v��n��"!�P 䮯���e+2@�y{����D6����Rcc�r��ǡ2�ޏ�$"�� �0�n#�����:i�/h�f��&����?�x,���Gu�b�����O#�ǿ�tK|�����&m	J�a��y��%�\�na��2U)˓���ޥ_���~vo������G�7nD&���*E(w�e�cLt�Y�+��(������cݺu8v�ulH�w�d�ؕ�+�����r���HN�+oupw�B���+ivn��6א;��4��rg��ҁ{�lB��S:���_�끟ﾊ�Y4�a����\C���|S!���V�HqQ�0~����D6�4-v�ȑ�deeI�D魮�}�oпt��������?.-䠸n����-[��}?N�Ijkk766�����&���U0�p�F�-6>�0����?�7o��Ç��s��7 V�}Ŋ�}7��+�<gƤ��'*N��K܍H8a̗�2ͧӧO3�>C}}}R�Lfw���	s�0�ҹ2:��q�u�V������ܑ��$�})�x����%K�������a�ו�>n�t1ې;��.frg����lB��S:��iȝ�vJ��3�N�"�C���j�5Ad�/���?"��ܹs4
=n��7u�:/��8"��_ {0�f���������-[�\�Cjkk������1��\{}�?�#��X8q�yܧ������SC�{cc#���x�~ON�u�����iӈE��ڟ���6	͐�w2�������8�d�4���H��7�*//�{�����bݔ���h*%%%�y�&.\���۷#����|�=�΀;���)��4��p;�����n�t4��;�픎frg����LC��S�Iא���F��𽺺����!�`�����g����GeO,�����)7��?(m��ߪ�����i�
�~��+�+��ѷ?|�o��.��$�ܧo�ҥ�x�"
A�3<<���Q��� ��ڜ���o�~W����4^P����f��g���uuu�tvϕIÛI
V��ֹ2��[���-�nMMM�����4%y�$k��Ǐ[ޱcǼ�v͕w[�8��.^WҴ1�N�j�!w��)]M7��p;����n�t6ݐ;�픮�rg���U��ܵ�
�[wBqgsrr>#�/9�����P(�5��W�*���@���;���������.]��� J�`0�����I�0��T�
����F������1�g����N����͜tNmhh�޽{��Ѩm��,�t+��p���~'vp�=�}��	��o���p����K��aT��ݪjӦM�D"8v�Չ��;����̗_~UUUX�n]J����ʩ��;�7��)ݽrａ���	_g����퐻�wg��;�����n'�+��p;��wC�=װ ��k&����)䮿�#��������b�ڸq��W�+������Ǐ�6c�� ���30q��P��r��g� _�`������w�
ѿ0OF���j���Ey��(�O}e���|+ E�������,X� ���n�Ɏ9#�t�]����X�2��g��͛(.��ř���uE�v'$�/�-�:7L�Rm��bO��=00�P(dus�4����ts��~��c���)[Ϧ☌9���+���I���C���*n�ŝ!w��I%�B���J�
�3�N����_�k�_�rg��T�!�� <{Bq��u�� JM�b?��x�S2��³�}�����0�>W���Ce�a|����*�R�<�~����ywT���އ}�I����b)	�f��۷��W_���4s>�'N��C=�L�t�=lu�t��n���9OE��Lt��Y�����n�����̽se&�`����q��5\�p��ݕ�ӗ/_�vvڹs�ޝb׺�n��Q��r���n'�L�3�N��rg��Ttg�]V���j&��n'�M
�3�N�����V�]U���\[[�u�ضm�.;v�ߙ��7�(�C��IP4{�ϑ��Z��������� �Rq
�~ּ{
�V\���0�?|�'#JO�v�x<(//���hvJJJp��9�[��ʮЦ����"Qs�o��A$ݗ�0�A3����b��.�{�(��ތ�ݕx�|)v�4E�y��N��t�t�R�v��q!7�AJN��K!�t�R��X��T�Z[:�s%%q���3�N�@�7�����A��z| R�퐻gs�q)K�p��r7�f�G�Q��IA��ҥ����*n'�H�����t��b���H1r�����gzo�:�!w���Ms����%��yP__��P(�A���PQ�"�5u��u4{�ϑ��(�����{ͣ`0x�رc��\�O(H+-�~-b'B J7z�nR�H<;7nġC�P\��gC�?7n���5kRؙNwڌ��[�$���Iݟxqwbb43'O���"��I`�E�=����:���g%�X�)�@V�y��7ߴ�̲Q2n��`��娮���{�5WN��O֭Q��S4vp�$��.d���%�b��IYr�o�-B��"U5��Q�Ț��/�\��vRր�>�[�1�"E���x�0�wms(Qw_MӾ�}�� �_�ּ�7oeP�������sa����BU���jjj:@4ς���766��yw��}�wJK�?/a��ٓ����׭��4sR �1�M02�]A��vY��lw:D����$�����>####VX��oxx;w���x�F^����9\zR�'�l�IseVVv�څ��.�8q��֭i�=7���E���Vн����BX����֕��g~m��k���������\γ��P��i/������Y0�jll��a߀��-�ЊKa�v�f��9��{���.���	��A�d;�cǎ��������nOF��<9�	c����Y�p!Ξ=���B��HN�����4���ScZ
��l	�ʍE-�
�2��$	0�5w���o�����'i.�<��yg`1PYY8���f\�z�k?����l����-I��\�5W�-��:��Rc�n""""""""r1�in��P�g5M��9�����&
}Ҽ{��=�w@���͎����Iס�Q�5�/F�^�gA�F���ϛ'�?4�~���у�}��A�N<ى���1��I���Ǐ�K�,444`����4v���ea�p>d��8���Iǥ ��� twV�Xw��3Rp&������x��LY�$[��Jsk��w	�f�U�VaŊ8v���uQ2~�ߺ9r���s���+�ZWj^���������������<{R�i��kuuugA�^$�zڼ��}�C�>��ҕ4s�ϒv�h��P�nٲ�
�������fee�+��R(F��~�d�l� �t�'��.���� ��H���p��H��7o���
�B^Ovu��D"I�G�)	�x^�*ˀ��H���?3#w7�e�>�N�N<88=����;��itt�L��۶m���R�'�[��AS�p�8|�0֬Y�%K���q�*��j]	O�&��C��M""""""""r)i���!(�y�c��`0�
��ļ�e(F[P	m��0�N�f��Y��{�j��| �4�s������_7��9���C��� J���P������؁rֶn݊_|���������ӧ3*�ng`s� �X��e������7?y vddtw�V:�K�Z�y�����
m
	�O�8��]�s��s��H!�H�޽{��Յ'N���DS)**B[[Ν;gH̴Xή�������	���:W零@+[ E��`0�������~';;[�.�b<{F��Y�Ն��	@߼*�4�K555�MJ��������c�����c��Ҋ7�4�6p�=�\�ŋ[]bivJJJp��)�w�}�v�e����Z�����H��-��������ܜ	z��偦O�n-��3��,�944���.-�$�0^�s7)++Áp�����s���t��5oSS�&߱cǴ��;p�t�D��H���3����^(�����'@��v��5��������wX�c��~d�x�a����SAӴcQ3�S�<}�<�b����7���(dUɋJڶǍ���[���5k��СC��9�U��v�/YY��ϓ������p��;m�s����ޛq�2_���sT�-�MB�7n�I�)�K��R�<˜�u��U&wk!І�~�z;v�
ggg�(��;�����(//�V��]��$�˺r`��u%<.^W�ki>��mP��iگIfDi�����666��ywT"sÖ��y	43��0���P�Wy""��ս
��5�~*�̓����F��緺G�z��ش��͛��ܜ�� O�x�������%lz�r�xJ�t����Iw������Ԥ+-��3��ׇ��z����d�͑�(�l�wp�n��h�,����:��I
6�n�jV444X�t�&JF�Y���V�Dee�9��*�Lp����	��ݼ3��V�P�a��;Q��4-������1��o��Y`"k���<�6C5��H]]ݏ@��_7o��7��{a��҈�haB�}`` 4w�_����ّ`X&t�3�9>>�0�g9D��e�
�O����Z{{;���@ӷz�j��]�oK��};jLE�]:_��l_a&���s���<p� ZZZp��Y��Cw%�ޫW�Z�#v�܉@ �u��J�1$y� ��Rpw�\IDDDDDDDD�&V�<�o�HuuuφB�7̻ۡ���[0#��y�x�a����泦��f�o�H!�`�ԱcǞ�4�'�=���VI.$�_QFo��cw�H(E����W��$n��V(LeNwp�N��#�p�VA�dnN������Pww�|�����{������s�f�� �WXɀ�],Z�ȺIp����E�4%�J
!�?�ǃm۶���߮�2�)<�\�9���'��������ȅ|>蛕���;���'A���2oJ5{�d��ێث�A�ǫ3�o��_�z�d��yӠ�� ��jao Q:�*�J���#++���9�.�׮]�ҥK�*;C�ccc	caݏ�1g��e�/X�0���J����]�ghɒ%p3������X6��.����/ɺR�aX��eӦM�D"V��}R M�DNN��ߗ^z�*�X�v�mse�9R�Y9�홀Ӹ�$""""""""��7o�2C���7vo'����B��̻J�y�m2�>C��0Zn�5P�a "���7�'��̻�B<[@�wJY��Ƥ�$�G��>|���gI�U�?^ـ��n���J�H�X,a�/셁��{��v��2_JH���ۦ;���qΛ!	��{��� lrxSB�#Z�р���2{����p8���a����#�]�v����ڭF
�X@S��ϡ�!<����ԧ>e�cN��]��8ܽ,� """"""""wѷ���@� M���0���m�s��Q��0�1ڦ̀z[�6�'��HQ����Rw��Z9�����]�&a���d��+WZ��\�����8q�7o�j$�.!};L�i�?*�a8Ic��$�M)8��{ee%�=MMM��>C���p39?�v-�<gJ��W'�wϕ���I�e�d�=9):x� ._��K�.�8��J��R4��ڊ���9�1�ZWz��v�����Iw���C۴��L�U[[�lcc�����녾i3b����Q.�=��� T�i���S�������B���C�UC[�ƕfͷ셉���+��d�SwY�bCKs$N%������Ύģ�ɫt�!��逻n����hoog��===���M��w���7�5�]�@B��OLLčutt�����$���2��:�̓˗/MM֊r;y�5'�]�A�C
�d=,�+�	��|v�;###I���n�I���J""""""""r}�h�P��iǂ��� R�db��0���B��:�g����4hҕY-m� "ř'�?5OJ߆B�� ���M:.]ܗ,Y�O]]Ν;�\@;]H`��ѣؽ{7Tbg�}x81Įg�7��� :;��WXOv>�c�q�mmm����"�L�=h��w��ιRHpӘ�[��A��Nr�nS�e����g444XkF��NR���uk��}l���X�ݙ�%��^?�&<	��4�+���������e���"�|+??���w@��M���Ӥ/]�X�m�5M�?���� R���������݅P�G�����7	k�
+�IP�w{I�v	,1�4{��Iw蒒�"//϶�Jp�
�ї����4vڴHQ���Pܘ̗t���rrr@�'������vvΕ"Yp��g���_�.��"�t	t_6bᱸq).�� �>���.�8q��� ���~���}������.�	��ߙ�(č�+u�DDDDDDDDD.�o��b$@���o߾�P(������0n\��Ӥ��A1��o@�̓Q����[�1�E(B�^���C �o��$���$�(]�������*f�M�n�ܽ�%��lI���<,��e5	�k����P(d{'n7`�l���,��5������Ěe5F���nmm�\YY8�����ƍV�$��ؓ�������g��+**������&��.���(����;�H~���i�[WWQ0��c�K�]���"ʀ��0�>M�z[<�A�!"����x<_�*'#]�~���xD�-����^�c���.,,D4͎t1mnnƪU���� �^{���e3�q3��bd���4v�|WΒ�Ƥ3��� �o7��0�b��Gm�z[R�MB�v�dA}ȇ��e:w�@�-	���6k�`1��]����V��o�S�{-Xp�To���5'����;M%/��䖠�*w"""""""""��~_��RH��e����K�P�E��~(�j��ܓ�{c�}4�H�j-T"�) � ۶m{�������Eh��p�4X���t�$gl޼����4s��|�2V�\y�Δ�@��2U�=�m������{� h�X,f͙rL��/�{,M����=�]Mt�?؝p@8o!�d�t�)��#˷ �}3nL�I)�\�|9hv�5�u�V��vCC�UDǢ"w�c���dZ�_)&�������5S�+}�����tO����bI D�0���4M����f �#��1�>+�o�����Q��
B�d�N�}�z���$���~k�{	D��֭[���V�}n!��5�X#���X�L���4�{8p�
�n	,��*y7~��5W�%D�.�3�D��'�w��)\��t��U�,�'y��+E`ٖ��ׯ_g��ҽ}�޽�y�&Μ9ÂI�n�3-j������I��ۻ(Lp���00�'i/4/�DDDDDDDD��e���e����'�����.T��}�j�.���Ӡ�� �<�q��	e�h4����4��C�%ˁ@.02���]��?���cQ�doٲd�ŋ�wޱ�÷�HS�I�+]���Mp���} �i>%N�)�	!�t)&��ƍ777[�C�z뭷�.�4}�����ě��.���v��-��޼
NҲ��|�JV�$�@p'�TUUY���&tuu!??��***f��d�#	�www��8��2��5'�+�ޕ�����g��Vť�me&�G���K�ɽ��{����\kV/Bv�R�fd�W�w�2ג��(.����a�}����JP�0s?#���g��@$e�@��W9�s�|�~���̳̅��m�b(d$<�S]]=
��o��WP�&]�p�'ܧ��@!�B��@���o�>`��~d��T���W�C��F�'M� ��C�č3��,�>~��)+pB3���������o�m��ʇ��Éy��p����tv%���z;z&�/^�7�ΰ,ؙ�X,��z�����c'Y��eX3���o�>�6��d�Vb��9n��%�f�M�6Ys���w��\�-����zó��L4�xaݛ_�˝�;�ۉs%�{/,��MUXX���/`hh��������˱xqth�4m�h���g��X��>_���#�}���w��*�XZ��ܙ����H$��ϴ3���֬�Ć�(+ɼb#��s�|7n�t������4?*+�͹��|���Ѯ\��x��9��jU?�q�FN\�����w4MS(�xt�ߋt&[�
�z	D�K
8���_NF�S�]L�3��,vڜ���l���Ϻ������,aM	�M6�-D��a���{Y�q��5���č���������p�ӧO3�>Cr�H��x��lǋ�N�1����B��������Y�n����ر�Z/H�]�d]��V�.$�eee�<��D�%�~�J
�+����ڎ��K�����z?I.6�7�q!w	�_�z��K��Nע��ڇ��Er�p�����}A��`���ל�J���9�o	��<݊H��rn02ԇ.eT�]���uch���b�!�hEƅ�%���v�:���X� ��i.e2M����t)��aô��7��UVA+P'�a�P�ܷo_Djll����Q�WMy2�t���A�����Ʈ^��H$�n�?�߶m���+�X?�9�χ�'O⡇B��3��ߟ�[ص1�~vN�$��PB��5���Kw7��[[[]쟋��j�-v	�x4��{[[��+�$�ȗY����ue��7&�Z�;���j}��)�<p��ULp��Y��d���DGFF���
*q�����%ʴ���p;�H���o��a�@�!�Q!���0Ν��X4l�)3�-t/1�����͌���p{x|��kS�`dTȝ�vwʴ���p;�CW+4�i�@����`8
=e��(@+,�VQ��s���]�=h�j]�5�π(��ڵk�<�h�}
�W���Q�����_��V��x�
[��I�A<�H�Z�>>::
����R+ĕN�9�����Z�=O�ge�eBB��uCH��,���DG�D�?�u�+W�0@9C���t��Ǐ�ۣ�hܘ�6s�|N�$��b�wY��$�h=�[�h�ukjjBww7��޿��VUUe�c%�Kh�k��p'J.SB���X���nw�L	�K�����!�Mf������dFȝ�vw˔�;��6�=�V����4�p]]��2�dg�c]����] p�;��A[�

�}�^Q��!	�ßm�aܼ���-(G΢���7~��9��a�:t�!�9��k׮���Ǉ����˦t��܍X���p�eN��j�M� �z���Qܸ	�Fª��ff��Š[��u�S�/�vû~!��gq��S�µ�V ��7~��P�lڴ	�pG�AVV�u#���֮s�����C�d��J\�v�����BK��:Q:R=��p;�r���W�Cv�N���n'�C�n��v�S;��p;	�C���O�Zd���X,��2\VV֡p8<n�U�ũ/[�ث�ASc�����nun���� +�(�y<�N�ܘδ%�p��P�a_B�]:c�C9KH׮]�:�����;v�@:(++�����dќRt�;����sA����J�K����vkW7��;w*p���>vo�Cyy��)��d�Z���z��!;��!o��}����f+`��+�aF��|سg�U���S��  ��IDAT�h��4�6����J�^3ɺ�_�B\���@�s%ѽ�ro�܏��6�rg��nS5��p;�G͐��p���hȝ�v���!w+��΢e�IH%��Q�����B��w�C��#��{�/�*4M㉈\a˖-̓�E��j(�Z�6�����~/��?�Ʈ\����1dg�uqU5\�b	��Ha���0rs�7�-E
vv��.H$�8��X�ـ����J<���F�_M?s�k�ұ���g����;���IQН:::0^�����f���{��9Zv~ظq#(�� i����t钵�g��:�/_n�cMp��p�J��Q-�.��N���N���n��T�3�N��
����nj1��}t�Z!w+�~�C�= �M�����v�kb�iK�C!gjkk���$Ck�Õ�kj5ߞ�߅V\
�D3_�?�{��F��'#J���@�=0b�� �a	^oٲ��۷����,&����������6uݾ��?WF�C1g?�׳s�.��(wE|�?u���ۇL'�����A�744�ݻw�n�b�@���帜���ɓ'X�+p���B���=Y���O:.�@�ϟ�+WZ7ymHW��.���5��ŋm{�dw��Ck8��1�Q?�DӥJȝ�v��"!w��i*���n���r�n��p;%�F���p� ��H��;���R���9�1SHn"[�����@/(9��F�J��-[���K����4Ms6�b�wJ޼R�U����W���~�m�S@�>_�~P����<���`ѢE��3�����Xґ~tt4a�_����i!݅��྇������;w�
���M7�d�}f�����t˂l�dA{���8[���3 ���b5���X���q	�������vi��@)��z��_:�5��?�0>>n�0YV�"��>�I1��󃈦/�C���=�yȝ�v��t�3�N���!w�����;��p;MG���/_@{{��җ��B^�K���6566�Z,+@r��S�O�W��B�P���>�iW%�>��do�R� �|S3�qh��~8!�.AF�jgWjJ.⥗^Baa!h�<������Ċ��m{�daM�ibpdNӳp��G����ӧQ__�L%~�413�m۶t��Sp����-��gTΕS+���M
�߼y�432��ٳ]]]8qℭk�����mJ';�$�U����4N�N���n�iKӐ;��4]�rg���/=C�����gȝ�v��t�3��<-7�<�B���K��{�����<�?X�A�:J����-�*x""�ټysK(�f�M���A7���s �o�������7&]����Q]]r�,^����w��T%%%8u��ﾔ���J[Og�i��E�8I�:��U�}���X4n�����耻�f?�;��M.x�Ձ7�����|�ysbb"n��ٳȮ��1�9��-@���0.œ����28p /^ĵk�Xh�&�\[UUe��%�k��/Dk�8��@D��n!�����p;�D���n��J����P��v���
�O��8�t��v���
�3�N��n!w��SD2����{9���Eb��뚦)p_��w�-�7��0n%Bn�:T��Op�4�X�����y6n\�:2��k֬��C��Es����N���=U$^QQa�㍍�%"���p�cNӲr��6M͛_���	�^455YA�L4KGl��13r,��Ձ�cw1�HV�t���u?NF�t����(����>O�ё��в�d�=�H��U�V�رc�|��:��>4�.�ɺxt4q��+��َ0b1�/fzp'��t	�3�N��&!w��i��%�.��s�1�N��!w��i��#�n���uah��v��t	�3ܞ:Z�B�B�4f
ɍ^�"�(��w��+s����) �1�d3b���r�B�DsUT�ᄀ{(��>�1SD�Ν;��N~~>�=�]�v��{JA��������G�+��=�yr
@�V��	���q�;q&vq���<Ό���r7����q��kr�].6]�.�ӗ
<9���(9��C�}�����eg����\�n$P�u�Vk'YK��(��t�����.R4i$�h�U�MWz�4����@D6��;��4g�ro��U��i�;�~;��2�N�5�!w��i��?��t��Cο���5�!�+�nO!�lTaFD.B�����M�}���S�OM�2�U/�A�[$��x<o�b1(A��-e���O���ߏ����ŋ����<	�ej�T�0V?
S��/^l��uvv&�:Ύ�0��4oNj�7Օl������ƍ���p�`���}���V�H555��TUU�����B�;�9sڲmp��b�{*��S	w�O�?��{��ғ�8p ---8�|��St˲e�l-�L:-X�����4N�GBG�sij?�����nќ�Fq��#�!s��tv���v�+	�߸�CK}hgG';��b���EW�?�sq_� ��d�[!�+ù�Q������d	�_�3g���Ñ�y��u���B��X,vD.�q�ơP(tټk_��hť��D#�D�OA+��BF�xD�̱�/�Dj߆M-w�Vd/\����q��d�=uv��iu�d��ّ�cǎY�,���������##��g�,Ź�q8M�=�9M��J�}�g_�ojjʸ��F�c��O�%%%�[����]В���A��O�i,����G�	":�7.�J��ߢE����ӧ�ך�C�[�n�m�%E����̛_����)h
��\Id+)�F����N1��8�}��	LL"���!��Lz�<��v���. �#}汜ګ�1^%��1<d΋�)����Dv��@$��5����k��
���"w�\a��%���������0�>��-�����v�B!i/��+�r��r�ҝ�B�w+n���?�S?��˃T�.�&5�aìI��ʕ+X�|�������mm�ߘ�T���� ��eSK�V˪*��xB�]�d2g�۷�"�;"d96l� z���������7&��}1�4g�u�����E��⺏����7��܌��,X��A*ظq���jhh�^w~?�}�TTT���̶Ǔb�d;�eWV����t�cw""""""""r��׷m�����D�I2��AڂJܧ���ʜ���fRmuiN+]pkW�Xj�&�J�Ϡ���W�-�O�8�`0J���Z:t��Š���y��ŋ�ܳ��m!I I�i�g��`�Ncif��~׾�9��{��2&�~����g�������[d>�.�v������D�ةS��[����H<}%;>�p�P�>�(H�:ޱc��C�����Ά�X�~���'����H�2\��y���<�x���������\D�XݖU�i���k�qJS��_FM�W ��)t��b� r/9��>��ZQ	��.��r�U���;�Ǎ�����ؚ5k���� �,Iq���ǭb'H�v;��H'�H$�0�e�&���fzO��͙�,@aͣ�;�t���7p��e�X��kmmEQQh�V�^z�t$��ʲ�q��x�x����Y4}�oA9"�EZG��#�<���(��� ����q�.]���F�\�Y�F1<<�0�U��o�!s~�(ΕDDDDDDDD�6Zq�rW�a�ȥt]�0�����Sb�}
F�:���D.�i�UNF�/ p�4R����ϟ��K/X��S�,]�.\`xh�����v�+�{{ee���)�ɴ`�F�4����f�|�/&��+���|��ʕ+�fH����Ձn��%K�������V��;�%�N�)5M�''4=ҽ�쁟A��7.kJY[�[��9����ɓ���Gnn.hn6o�lk���^�}�]Q��S��'���������m�Bu��I�
D.5::zY2*���Lf*�OA�W�bvGMM�0�\*�]V�#�����K��������w���믿��{�:���8}��#�o�@W�%vϞ=�>��y�A___¸t�|�_Bc�p�7�4s�5� �x&z[��C�>�O @U/^�vB�髪��G
��~��+A�����~�~N����w�2���5�~�'����݁pW[MM�UH��o���p�:K����vop�L�f��(C�@3������,| """"""""��S'�*�*�Ԯ]�C�P�y��.��d��4u����t]��Tw�4"��J�it��q�p��?��]�S��� �h4{�����Cv��ɱ}'�����_(]��'��
� �̳au'�������ōK�O�̃BEmmm(,T�}OZ�0!���ǩ����s�ӽ^d���b���^����`��Kq�o������\�6	��ڵ�Zk��Tv�P��<]�ݽ}ttccc	��Z|�j?R�ù����������H����"w�lm���iƝr�OE���*�\,�\�.r*��x2��S����hhh�B,�:;w��+����|��!���x衇ly��˗�B2�W���H����i��^8��υ泿˲[����|�w#7~��a�߿��G�$;GHH����W<�F�D7���N����jq��yDV�ӽ�5�c�A3']�'ܥ��ȑ#x�G@�B�X�\�v���$;],\����L�+�������kH�+��A��1WHn'���^�����Tp��BM�\l۶mݡPh¼�������?�������A�5n��?�1x�vfL!�[VV���+))�W�W����HXK~vjmm�-����+���1��l΍��
��'7���kWlݺ*�`\^�:��) ۽{7�	�;ѽ]ܼy3a�ȩ����&;�@�A3WR�1\/X��@|A�K/�d�t���#�L!k��+WZ��GFF@����`0h�cJ����@�xV�b���D����t�z�DDDDDDDD�>
e
Ƕlْ�mĉҔa�J��4wJ��8�\e�nQ�y�D��Ɉ�Ԃ��6!����nu�ݴi(u��>t���D�ycr��U+p%�%�NlO����E*����U>�����x����K(��@��҂���ܒiV�X������V1������R��XM{s���t�y�P�������ōKAM(����A�C�ú�:����7�@NN������}�yM%+��^���]�#8W�k��ܒ�B"�*�g�ܩ��SZv��̨��h�ƓѭEY��s�%��Sq�O�W\�po| W�����������Hh�$@t��1��cV�������mmm���H�U�X�߼�|�~Ov�<��)�t �e�1r�D���k�p��Y���鶛������Q��$��yl9Nv蕣���8M�=���c.*������?E,�;��$�f��e9��ݻ���8y�$5� ;]�������aX��L��k����N�Ǆ�����������JSg�df
��T��j>��&�ώ�F�w�e)�Q�ʄ�A�ɨK.�;MNDDiH��P�������B���s�p��E�^��:�-��{�;=����%�f��������m�Y���,�)����j� R�]6�#������&�?��3�ܥ�rnn.h��ѨT�[�e8�6����I��1�� E:�N`ω��%;?����7.�BYߨ2O�̕�����V���q�X�v���NCCC��	�%����N����c݈��������\ɧ��"�0R�!QzS"�n��;�	pO��*b�X�\�\���:�rʥ����g����#2_7��s��s��(�v�؁�Ǐ#'���ِ`{CC���7���r�J�=������v���%�{Ex�� z�4M���c��.�;>����	�^477[��u��!�E"vP�!)�����RUU���|G[vC�셗^A��_#�堹[��/�땿5ߨ���U*�ٓ߱�eG	b�uǐ��2�Y������J�s���qӳ-=��
�|ΕDDDDDDDD�b5�?��9!�(�Iw��
i�k��1㦚Z!���/�\J_�?�*Z��[q�O�f�y m���=y�{hee����1����֟A�(]�~=��F�V���}HOn14�Ǔ]4o�9_~7��儯=���ip���3����x�:�M:J��˖-s�e���M)�x{���28M��g�a��kQ��Q���lܸ���;��~)�H!�֭[188h�eu��V�u�`��2�ޞ�p2g��x�Bj��Y8IDDDDDDDDn���i��F���A����pg�09>+�(t��/�	���T�D�)�M�ׂ�~m��1��q���>?�mۆ�_~����S�NM+�.!���j����֤!$)(9�S�h,5w;ۮ���|၎�q	o�9s6l@:��b�1�S烷y'�͛7�nY�j�c!իW�&���������/����T~��	w������<�d�����������D

�`ӦM(,,��q��wR�»����ڌT`�$����"�J�q�\,S�u`x��,���d��>�^/��z���q2�rʥ���-Ƃ�E�3�7.]�%���]�3���-Zdu���)))ASS�2��+VX]���F���>RT����Hݗm��^֮�|>i��~��X�~=ұ��ĉVؐ�o``��K�.N=ҕxr��p8����n\ ��#����>��M0�t(n����p�#�e��dM+���~����+Fqq16n�h��[;]L��x�9ӅT��������������M��l�K�N�\!s�"��S�i�d���N�5^^vK��W��D����X|��{�����/C��_�X�f:dehv:::���R0��<�UUU�_�T:1�xz�d��H_iʺ�{ٽ�1Suq�q��}�v����>G:�f*�;�U �R$�۝r��儱�/����C*�#�3��̤��x�'��t������7ް�f~��Dv�x����Bִ�i:���R�U��U8����	DDDDDDDDDӢH�P�u5�TD�x<�r�W	^u2˩�g%����A�r�a�+���� a��~-O�f���+W
�P__J�͛7���Yvm͜�y%D�s�΄��|>�]����)]�%��PQ5N7��{�t$��#�S��{������B�מz�)���Y�X�8{�,��3$]�y޳vK�vqq"�)�y��;I�Pco y�wo�H��U�PT�!�&n\֕o��jkkA�#k�]�vY;d�������)v�(**��q���166�0XV���������s%�J�f
���j�ƹI)3㦒f���?�� r9]׽�
�[U*���*�O�|�/1�Е.�[�la�:������Ԅ��|���9bpp0�9��N��q4M�
�zO�y:HQ���h�^���௠�?F��-n\����#�<�t!�
p7��q�c�J�-[��9(Y���_|��_@*�� ;;h�'������y2�/$�@555�NP��`����q��5\�p��`x*-^���ն?��c��������-Õ�+H��w"""""""""(��1�����b1�2MvbQP"&^�0"�0y<���ϙh̓Q�'��:s���%�>���7��ݍÇ�������q��1��egg��7������w�$�TRbw�!���'�ZW�j�=��p��V���g���W������s�a�֭(--�|� 1��3���cu�w;	��|���VǍ�<zrt!r�ˑ
��J�sr�܇��GO�?ō˹��W_�޽{A�t�R����h����P���;v�p䱥hNv��,���t��"�v	����@��������7iv��s�?ij1���B!TM�x2"�3_Jza�Ie{�?�3������g�"��&Ж͞t	�~�:�,Yb6�/_����x�b�q	P�Ж��1�T����x̤B���G�����Ƹq	�=����_�%�79.�(��d.���ygݺup��4���ի	�O��v|��{�������'}ǟF,<7���O[�ʼ<v�'XEErD�1ʉ]v� ��޽~��K�<��ٙ�=�h+GK�5���|@DDDDDDDDDBU#��L!ѭׁ*w��r���D�i�ϓѭ��
'#-�*�;ߢǿ���Xܸ�N�x�	��/�2(�$���/Z�l�9]�q��9�^�ڱ�f[[�`~���J��NM�]�ؽ=u4K>�G8��}	_
�Bعs'6n܈�"�%獙��������f2g�_��р��,�T *�HW
�"ߗ�T�v��鳢0����x��h}�w�ƥ[�SO=�O�� YYYصk���p��	������;V�+;Ēlw���/kC�xr��y��#�P���aJ4%rR4�k�\d�ܤpO&<UȋD.�ŲT8�"�H%�uE��G�⹸��Ǐ���	�6m���W�X���h�x�Q^^n��lJHS�x�W��K�+���s�g�n*�ߋ�������	_��w���~���։�����ϐ
�J�I1��]������ɞz���oH)��嗁R���_A׫�p�͸��^{<����!�����v �v�
��֬Yc͗N������q_Q^����h?R���DDDDDDDDDwP��23��z�����]m�'�Vw�U����A1T�P��m�~���������%��v��yl��ʕ+q��%�1�	�n߾���R�n{xUX�$�L���͑EI���!^���ŒO�!�O��|�����>�,{�1��t"w2���d�ݻw�͖,Y��
����/\��0jl��ڏ!��HoA����^-���å��Lܸ�����/}�KV1ѝ$<�j�*���V1aNNjvw��'e�%'H��dE@��Z��j;Rœ�=+ """""""""��4�L��!D)�ŊUil��s�Q��b�=	C��a��L�5^vp'��+V��C_��'�k�xGG�������8(�jkkq��ydee��o����v���qee�m�-]�����~m��o�F��lx��ٕ�X��/���~;�k?����e�R�3���[((( M�̭n�J���˗;�=�_�nup����]A`-RA�t�
�R��O�����Ѕ�q�W�\��Çq��AM&<o۶���hhh@ ���ןIv�سg�c?Ggg�5/NXr?�8?�p4�T�ڷf&""""""""��d��-����%�tpWfnI)ܓ��\EC��4�'#"Ue��8٩�C_A���X����C�Y�a�H�SRRb^p�>���q��w�,A)��C��.�ۓ���?�(�D4u�h�k�LU��_Go�?c��ٸq����o}_��WRʓ ��ϝgB���[�­�Bvgq�<�p���g~��m��T��Y�p��3�O�~�/p�A��m�p����������{�
O�81o;�ϱo�>���###V��d��y,Ņ���������Q&��F�P"g�C�06
JĀ{2�(�d���!ݱ�;�E���� �T���X��?�;��pܸT9~���W��U�|��Ҏ;p��Q���Ze�-^�۷o����t�\�hќ_�����_�t�1V�jW
��g���W�?2_.�������U0{	�>����G>�������
���E�Q�IGd)r�{�;�c|��ҥK�X����	�Z��ّx��ޏ��"n~�kq��p�*���?��Zt��āp��kW�����}o9G�߿����<�̏���I��/�ǏBH%_q���������h��A(B�,������
�Sܧ24 �*�Ɉ\��_�6����e���Y�%(��!�>���~��������������h{�a;q��h�$Mo�.ZZ(��A��2�-�e��=.�{)pi��(���h��.2mgڎ�xｇ�q���b[�t���s8��X�t��G���ZZD��[n�,x(\CaY�R
���L�ܹ�gP����^ѱx�(TEAy_�������#�����[�i��A�돎���+V�\�e˖�>��<>L��y�fD"*�X�v-,��~<@E4�^��
��R�]�e�5!��?
	�����G��p��Q?��7�xCt�fl2�V�+D�'���j	��tl�s<�����X��Ex�ކ����S�v�#x��1�c�1�c��B��$�

����.0�$	�s���Vן>�ɀ�L��`,�EGGgC���I.�C?A��71�Q7��{������E8�ϦM���k�!11l<��I!$��������L�Ե�����e��D�ܙ�!g�ބ��Ѱ��1�܂��G_���y��)t��_�_��E��@������hhh("WŠ@(��ݹ��ۚ��q?��W��� X��	��9�ՁE�J�v�60��F���Oc�ҥs��
��ĥ�^*Ƙ#G���@�DA�I�W���#P� ���{������'�L6���X�8G�p��&��^?���GŰ3��0Ϊ�E�Bo6{��cX���Վa�l��1<4����q�����EΜ�m\��3�sb6gF���}��3<�<�E{��@�W���%E�P�L�_p��&���悱f6�s!�~>1����{�/p�{��	���)���O���l�a��.����	��,%%W\qŤ݈)����.���A���ӧE��q喥8]�
[["����������tuu��'���w����z�"�M�1wq�z-�_���B�nt�c
�����;kkkq¼qI�2���&���b�lG��E�?�s�˅G}=��V+�

��ܯ�����s�e��ٻv�+
umojj�y�e�v����<�[��}&��1vz�T���F(��f!.��?��q�,8Q\"�[|\2R�m�|0��׌S��mG9b����Kҳ��p���V�u�!��f+�e��j�9�����!T�T�v�)Rf�<D��f��7����^o�'�))H��!����l�X��,�-�8�����'����SO�o��V�i�����"z�)��b� a��H��>����Q?����?�8>�O ��ɴ�4��梤��t.Dyy9�ΡΚ�as�݈)HG_�����Kuu����p��Z���#
P�����_>�ֽ����СC�C�Ν;��v�?.�I�h{��Q��ՁM�^�TI֬Y�������ٳgE���h���������l�%>pݗ��-|�w�[��G���/��o��Sq�ʕ+���)
.����?m�N��kL��B�T,�{�ndee!P�0���^��rd.ßk���fV���XHP��d����	��;�
��M����uj��!w6sn?^R�p;�GK8��fL�۫�Bn'��ͭrg��p;��ͭ�rg�B���%�	������9�2e�^o.�P���l�H��ǙB8��<�V���\�打+,")��Y����p����#5���yqq1^}�U\u�Us~��������֭�
�G���|�X��222�gϞI;�_��ö��N9�Dݷ)��9.i�İ+�_�ْ�xO�~��;�&��O�����ggg#''gNo�^T�AE�]v��ߏ��0�苋+V �P�=��	�2Bc�XO=�,;?-V�Z邻�u�λ��(��%Pݣ�Х9����E!F Pq ��i@ݿi̬��&6ႎ*�9p��x��Z�x1�{��
l��I��9����8cY��:ߝ����-���
u�]�!w6SN�9��v���L�:ܮ�;�����V�����)hjw�,ܮ�;��P��ury��R�B��Ռ@bb���#G>z��O��������,�Y����{�T�
c~Q�b�}O���wC��F]��ϊ��U����(�B����?� 3��(��v����W��HC�uÞN'v����a��x"t�ӧ}��G�KQ��/�,��09b���du`�=�3��v����_�җf�aVܖɄ��X1^���;��`�Q�

E
:���I��@��V|w��@u�;��5x]�M�(X�R��':w������G���P|�����:����C�E���y��<V��v��%�+�9�T?;� 
�zu��������D�����kap�)�b�-y>c�e�p��C�l�΅�KCn�qȝM�� �v����)���8�Φ�\������pȝ̈́Q��:����	�p��E,�׻��,�Tp�Cmk�,�f3�4{�E EQ�BjO7�c�"v�%Xp۷P��ύ�9�}�Q<��CsF����Xܤ�^YY����v�؁7�|St �D˖-Ö-[0ӂ'
��1���}Q[RR"BɾtĮ���.�!%q��(�9�=_E�S����m��կp�����p��#7������.�������u�(��F��D���DQ�6�B�颱��̱Xt��Tڏ�+w!�l)��-�MO�u���+�=�ꨟS��?�)���/�IQ�М�_hy޼y�vΜ9�Ńa���V�����b,�ͧ����WS��.�#{=�_�î�~�nMʂb|c�z��n�qȝM����:���:n�2L�]�!w6u
ʪ�n�qȝM����:���0Z�]�!� ���@�M��L*c���Rd
�����w?�v�y^��͡��r{OO�2ȀOD,e^� ���FW�s�~Na����gx��gF���Ē%K&-S �B�������A���!--Mt�$tlP�úu�f���S'uФ�
_�s�8�}��/����x�&kb��ό/��/b���
�w�ɓ'��7�|�~wrr2�/_.^�t�B��6��ޡC�8�y^gg'6oތH�����K�"+�@�����Iz���!�ʯ �,щ0;"� L�I�vq��p���������p�w��&���Ŝ������R\\�+��k,�-Z$:�ahh��@��_~����̖��DCC��˨xq_w&:�L&���t0ƂG��K�n�qȝMƨ�v���d�p��� ��C�lr���8��&���}��0"����2f�]�!��R[��,Z	�,..��^�z�Ei2�*�
�※t"����}��1	uww�RE�q�OD,,)
��+���p���PWW��������β£��Tegg�0}EE���)ioJ�w�^$%%!�qr饗��~.�q���/�|�=f�����w������g0��v��kB�$h���/1Xwb�xI^y����c�Ν�����-\�P�7h������#V|�ϱ���	�K�~�uH�����Ͽ�������s�^'��`�gM���O�	��yT��`�[o�����cϞ=3��4�R��TW/�b���׋�;�Y������|q��/z����9�VE
�*���W�4٢P�G�7�N�X��|5���=ܮ�;����v�ܙ?F��8���3v�]�!w�߹p{�A��!��,D�xf��p{�q��:�5Ε$�nZ��O���#M��ƞۇ��А��D胍���(k�ɵI��E혗����,\����SB�W��;2: TPP 7�pÔ�T�k�B��ӧOGl�M
�S`&���P����ݻE��D�`
�SNG��ou �t���Tw7�N�B��?��K��r���O>���(�9
�Q�v����6�Ժ���W_}��S(>RQ ��+�@8�s')))A�M�H���8��DE�ՈI��`�$d@	b���N��˰�}�F�o?;�zJtצ�[��
/^�y��ќ�V�(++�=��B�L**koo����E�v�Gz�ZA���>߫h�ݗ��Ot �_�����<�1���urgc�n׉�����$+�ܙ K�]�!w6�
�����8��Ɠ#ܮ!��&��Qd	��8�25�=���;�(��-,,\	��bc�q�}޶�rC�ǎ����`,�h����tj�;g���s�OP��w����_a��۷O�{(�GA�ل��q�Fr���E��plii)�222D ��p��S��:kZ,�=s��+*&TE�Ƒ���P�� KLdt�74^������.���G��?��	;���ƊB��_]]]S�#���Z8p�oG��� �A�P�p�U�fT06StVUU��9���6�!~��taK��.��$��0PY����s:??��x���X�1��JZ�e�h.@����z��6�}Q���\����K���>/7/؈g�x1���b����Y�16��~Hn�qȝ�d��z{;���;�/ܮ�;�����V��s�;�'���:����n�q�= $궬�c��o�X),,\���ٚp�pBp����������;�(�$,�)��h�DXxK�u�O�����9}����Ft�^�l�ϿK����\,X�`N�u�^�n***��ԄHC�EEE"�N�8������J�0[kk�(�())�:_���o5�����!$ɥ\�TF������u?��E�S��~1
�Q���_����颿s�e��"$3d)�}}}صk�UZZ�.]��<�1����Q?~�����͖��+]Hjѽ�a����E�~N�����'b��(�N,n���2�Qi�*��b$�`�
�����+���o&�Չ��H�[�y�[�<ې���௬bM��50�����΅�K!+��s���҅�urg���urg���urgno�F�d�v���5ܮ��ܒ���<�*��e
eiv���3���'�6��!�K��	0!���O�͍���P��݂۾��3�*|n��)Da�x 999�.��ъ+D�x.�D�B��{���#*�D�z�}2�S��;�Աu.��s��)���H�<ߔ�a���BH�eꝺ�1e��C8�k�]���˨��?,:��ݷM&���D�}�������X�hzz:�~�mR��ٙ�pC��E�m�����x\Ѕ��ǞyQW�lA�OָT�q`r2٢��SO��+���](Lcޏ~�#|�s��B��B��@EG�6mBYY�X��m���b���8�?����2*v���\G���~W��&fa_�"�m�D��k���X��n�q�=r�3�.��kr�\���ur�\n���6ܮ�{$;n��3ܮ�{d�p��%������ Yh���}��9���3�"�e�e��_p��ZW�\
�"��jݦ��H�@�lcaO1a��~��_ߍ��#�.���ؤ0RVV���خ��@����3g��ݍH�u�V����v7��EW�@'�@f]]�N��+Ħ��lt��<���X���6^��x��=�8<�b����#�����xS�Ʋ�(�7A픔\��8v��P��m�6�:�R�X�W�
�h%��ї=���Op_�YX���O��k�|0���a��_�敗��Bihh�O�S|򓟼P�C+����A����U�h������3.*p�U�|����c�ޯ����?�ߙ�����C��i
��n'�Ԝ� 1��%ܮ�{�p�ѓe҇�u��Yd�p���;�z���%<�:^r��_�	�Sx��ur�L�n�q�}n��C�@T4$`������ cBQi��^�2�A��	��U������'�ر#4ߊ1|�h,Q�KD��O�	%_�WW�����E��/|�X�v-/^�`,	Da$����z���DD�W��K���(��y�fх5X(,\[[�7�n�I��K���p;=�6!��-K?�/G:��]N�O���+��׿�7\���&:���=����{�C��yH���+	�T����`/�G�v
�S�Xz�%t��0q�6[J��3��,�G�'���?�	�@/>��c��G>"
<��WG�@�9Q7w
A39P��+�zޤ�6ZY�V��ɹ��흝�?��yj�7aoIhV�&d�d�c,�z�,ܮ�C�,���v�ۅp����v��;��.-�p�N�'����7�an�QȽ���22��};N�v��!w��M8~��F��c,3��ކZ����$(c�w


R��RHB����[�	�����$�������Y0E��Pk��X$�%/��_7���.�Pkk+,X� �&u)��hOOh�$��|�r�ݻw��FEa�-[�-�F&��c�o0�	�Z2E	/��,,��q�?w�3�{��4>RG�n�A(W�^=�S���9
Jgdd�ѡ8�����pA]��cuLL��n?q��p������k��ύ,щ���w�c�%n���1j�ظˎ=���~>����L��7m�$�TD��n�EŮlONN��ߧ�tbb�xC���T477�p�/�Ɍδ|��Ԡv��[D��[�<0������4W
��M���_��y}~�Gtv�0<����
����Xܧ�b�z�w��k����=J������,���5 :�
���&�M_�-]q�hs��<�[چ�����fC4Ε'�G۾�" e
UU��s��rAml �O��v�x��T%{d��0��Y8~�x��咦�;WZ�H�`�}�%��֕���"N]���>4�PuUw8��_QQX�n��TTT�����Y�~=*++���):(,F���I���BLLV���XKh�k&{�B����^���|�ZxG����;��ƍ�����(--ŪU�F�e���(x饗�@ us���E8�06�ReG�999�?~Ћ��D��#G
�߻����~Q�v[j6X�I��~�tԢ��߹�3z�t�Mعs'Ξ=+
���z�ۣ�"�q�>�x͌%33S�+�J���k*���ο�Ґ��Mtqkn�<(&dn�ӥ�x�?���mO���1X��bcLVn���erkh�E���Z��}&�[wπ��������-�25�T�򂂂���|^�����Z94�^�r��B�[[�$w͵T}��EdXX�R;���Y���ۆ�<���]�5+�ᮻ�Б������y�CHԍ����� \������Xt�52
�Q0��l6[Po�:�R�U�v�bC���CR�i��`�+n�.m�|C�(����HMMuygg'N�:%B�ң�f���>�(�w�u׉ۦ�=ݦ��oذ��q}ѢE�!&
�;~k�D��w (����`�i��߂g��{A||<��^,[�L\F�c��;�J��P����F��B��
���������������������4�jQC�������34��T4ir�_��c�1�c�1�X��WC"UUwk����0F����« 	�N�� ZPPP�Z۟caLQ�k U�Z_�"U��=ȹ��V��B�]�t:q��I�Y�F���*���
us��cm߾G���u����D
6
�����j�|Ҵo�Ϯ��lP7b� ��_t�&,��+HL��ц�t4�1��LcX0P�x
�S7��G���(�'
���@V�y>///$c�N?o�_����/�F#aۻ
��t����uK��������%Q�q1
�S���vJ��¨[8�/'�<��sssE1k ��Ĉ���C4�9�΍��O���OV8�?�"�#քL0�c�1�c�1�fOtp���$iT�(
u��;kG�Yo2��Ajg
'��I�g� ���w��WZI����X�
?,2�7�mU�Z�e�x��?�}�m�u�k��c�D`3T]�)4�~�z������{2���( �M)4����ۧn�n��|S���}��(U���K���\6E����Z�����
<S�[��a���F�9
S��`�~Ac�Ν;���*��z�dP�p�ʕ�=���٢�~(Q!XP�}���r<S� ��!�Ȗ<,���;��/����?���� 99���4>��n�z�
��*���o����+eF�X���=�B�Y*d�������z����	�F(�U�Rs��1�c�1�c�167ԁ~��Ȕ�;
i�V�͔�l�N�fmj�i��q�}j���o� ��t���.S[EɁ$�e�`,yG�l���}�;a��kQ~ʂ���I|���8
"Q`��HIII�I[{{�$�S�=??���C}W�}X�v�l���*sn�_�e��x��o����,6�R�9ݱR�1��Z	��]�[S���郸m�6]����DȘV?�N��F]q���j455�%�^kt���b�	u��V	UPWG���i����O;��C:������T/�m�pt�p�����������;����N���ի�t��SV�X!�;T@I�K6��9�b����{(P��
&
���V��Dt�����+k���1�c�1�c��3OY	��ܗ>|x�֭[���0���{!	�傷����Hm�����*(��BڋtKAAA^~~~C�����gJ�X�q��a��c�"�׼ն(�����SR7풒,[�L��C�BRԍ�:1N��Mnn.���B*�����`;qiojkk�)ވ���ǽK�z�j�z���f�"�E��/�P�X�V��3c;��<�[�Z�4����$����
(���DCC�(R2rН�)˂��1=���z^O�>-�c�*.�s�6ą(�Nl�a�o�6w���sE����c�	(��̗��h\'����8qB��m6B��h*��3�?:$(
��l���G1X�P�T�*����SU��]��V��&�1�c�1�c�16���R`�; ��t���;K�Z��6@�g)�61N�Lu`6Kp?�����UU���!���B�5�k���܉]v�~��'q��oޣ���( �0"�)����!�H��������B�ŝ�G�V��g(��BH.�Յ���v�,�?Z��U֤�09b���	#]�^�5i=��-Ż�w�aФ� :��5����P��4�i�����R1^i�7��y�f]LL�x��+�c���������Rc�݊P���%>�Eq,�<�ݢs������d��[���������O}J��t4��U&(�N��P����!Z!������>G�Ĩ`A/
e�~B�Xqq�ߢIҗ�OUơ��u�����`�1�c�1�c��=	3A����%EQ��ecs�l6K�4�[&��p�q2��&H�Rpga���`�6�ʁ,z���4��H��G0�Z�sp���.݁z�?�q�s��:kR臺�/_�<��k)dH�i��;7),)k �B�TD�N��999X�b���n�����Q���g%4����D'��(�9�V�`�����O֝�{�Z3�K5�)�L�P�~A�R�h���{uu�X1!Ԩ�ƨ�C]��͛�⣉�qU^^.�|9x���� a���s�My��iҎAQ�=�{)*H���Z�������}�c��$������b>rq��P����ҥK��:MMMb�( �Ή���v�����̙3��h��+a5�����3t�B�d�#=O�z�c�1�c�1��{jc=����C��=J��
�X�	]g�P�i�p�}
��Ӑ̦���U�6m�W+����p����8۪|w��#f�V��$��!��C�Ctt������Eȝ:]��vkh��&��h�<�o$�����{JJ
�,Y"B[��OGWW�x��v��Ec��R��m��du������a8[*�~:z������������13ie#��@��m�DAMMMΞ=+�����Ӄ={��hǅUB�y�m�@�ߪ%���G�[�~7B���M��ż�34ŕs�1/�Ggl*~�����܃�k�^��V�())�w��m4O�����<���YQi�P�����tl�^!���������ɂƸ5x�ʆa��dO[�j��R�1�c�1�c��%U���i�6n�,�^���;3����TU]Yhc�zV�LrHp�}
ԮхY�Ȃ,<Ͻ��3`,L�7�rܹҊE WO3F:f�w�K��x��o�#�]?��f?�����P i��b�  7i3B�⩠��;'�/&&Ftk�P�Q���($F�MGG���x��swj���
l�3�Ğ�w'F�k�crfE�I��LO�w#;-��u���Eȝ���͡?�(����'6
�WUU��{___����t�%�x�j �}�H��/�w���M��?�싨�~7bs6 �8���#��
����h�|��`rD���>���p�%�\������bnI��C�B����h�מ>��Xi$���cA�%N鹢b	Z	�
���%N[W�
���(�[�6�N c�1�c�1�c,�Բb@����}��}qϞ=���Ř����aHDmn��3�U�#ܧH=uT����(�NF��'#Fޫm�L��/cኺk��W�=�3��c�K���o�g��^�/�����S�D��:o���}���"�����v�n�			"�3Sj����|Q �(ҋѿ���~�.���4<ב����vn'��\����U�Hg=\����U#���+������Dޤβ4fe�BcΆ�Fcdmm���߽k�.���)���ڍ8V�D��������A��"*iB�����ۦ��u��`��񝰧��O~^�57�pè�[[[�8I+EEE�hh�F]�i���hu�[�}gb�1��J3�P�5=n�{�#�]�q�^E���[�qҚ(�g��1�c�1�c���{�(��I���}���=�������g
���S�9V ӿ\����&m�$RUZ��jC-G��fk%�.��>�-q����{�qm�n_�LA偁,_�\tP7
-R0�6�J!���.��B��	k�L���;���<���@VV�]QX��(|DaM��
:�s�|Kz�B_�`K�s�T5\l
T�K����&�-1xͻ�%{�gU���P����z5�k��mܸQtoll[KKˬ
oƢsE(:���ŉ��:�JF�'Ϝ9�#1���?���/��C(Yb�8��T/��p�w`.De�G��˿����}�ݣ�T�v��1,[�L�EF�p8.�D�Sz��ܒ6* ��8I�%���ԩ},:G�y�V��+&/�/AI[���Eޖf��`�c�1�c�1�ZS	��J�q?sKQ�{�w&���oQUuj���/ ��OU�	�.����NF���,��z��B"�c��X8r�wb���:��-6���%���Sh|�y����](�SXX(�F$
5�F]�)�D!N}����� �`J}�(F�٩���Q'bP �:��+*P��)��Z}Fܡ!Y�RaM�/��~�V���\SMV�H���ᝫ�a�����
�Q��5d����b�
n�n�����Ŵ�t5�w�*��k4~�X��;h�J�~���eee�(�g�⩣�y�C�?6�� �=F�t��9W����kM^�E�ʞ�"�������aj��JJJD!��c�p5�q��r�h|��OZ9H�[�{Itt���8I{#�2�'�����4�����sg�z��w6���%PL���c�1�c�1�X�RUxO������G�Y�e˖20&9UU?���@-=	65r$�@�ZVe�H�NF[��'m�Լ^�g@�v%��DX��ޔ�t����ЛI�z+N�.G�O��o~���L�$B�p
U��*
&Q�w
']��gvv��dff���}�⽢H5�p,z����7�X�*B_d`���-%,����1�Qؕ��gC��]��+�IqQ>�F�Aԭ�V^0z��l6_pz�(�I�
b�{��L��S��6����r
h���\�(�.�yh,*����������7�ߵ��oC���v�3�hǽ|�5��3�g{5TO`�?�x�|�a4��0���o�#��+�$/���$�*��״h~�R��N�N�(���$����B�P�1��X)K����7��=�~��h���/M�6@�]#yP,s{�c�1�c�1�c�MN=Q�pW4���c+**��z�;!o�	rgS#�7L!&�r��l�)m�0&��Ǐ��\�; �ޒ`,\���?Q��1��������]����(�HA%
d˄�Iqqqb������Gmԑ���tm��S�O
�{��!B���m���"E�R�Q������a{^��AC_ C��`�E���'��,L�^8۪��
�M��/�zҰ�����)�W]]-��2��4V��{�i\�׼��EB�懶~Fc�t�H㤾Q8~�x9ׁ�P�1�B��
�\��^F������F�n82��=��&�t5��Ld^� �s7���p�\u�U��B��cǎ!''G�	��4V�F��訐e켒�ȋ甴�N1����R��1��R�xnC�[UU�(�����#�E�_���N�W��ܞ�X�/�c�1�c�1�X�'�^�h�!�;<���۷��1Iy<�����7͝��x��`��=�̭����_�$�v�?������N��@���p{��k�c�K�冯���W̯��ݻ�]��:'O�ȩ���!m=(46�~1
!Q�r���)�Cv}���vʤ����hmm]6�2��l��_Z��7� Q�V82�@1�}̲��X�	~�\�-	/{v���kxǪ�c!�TB�w3i���'/^c,
pRHU#i���S����I�����	T�@�M����f���b(;>�#�&���A�{�6u�׃��*�{�z��+wÞ�/=� ���p�=��.�:=���ގe˖��LVz'���-�I�m���s�>F��qŊ�n����d���Q)x�7增�����0G'�1�c�1�c�1�@?ԳeP���DV��ߴ������=���xn�d�p��O��P��	JF$B�1uq�,�����c\.׿A2ޣ��X8p�4���8�Ύs�bC����p��O���QQQ�F�<�林�����3
�̩�'���.���u'���t����_�Y��uvxU���Mf82�B���x3�<�ݢs;7CE5�P�q-Zʊp�~$����J��+++��>))	��W�y`��J�uvv���B�����a�kK@���@�P��--&��ܠ gk�.gHnߚ��>�8^�����ᮻ�+F]����=���l��P$��^ :� �
�=ńL&4[��Lt��w"��LX���c�1�c�1�-o�!��
��wk��߿��;v�~/�f���|��զ��`S'�l�Co���[!��<�]^R��fdd�c��ȕV��c�S�#p���.�~�إ��o�
�詇q��U�[�XԱ������"��7���[T8�w�7:
!Q�v�9�K2�֝��~/�Bt#�\
�-
,L�^�P!������M�Cov�Ś��W����"����������pH��O@��A�M3����w/�C����m)��KL�aD2*�U�]G�eY����\�G~�M��-����Gu&�W;��͒%K���]��Y[[�(���rB�8�AAM(��[�|0�c�1�c�1�B�s�-�o����D��v�}��G`L"���v�B2�o�Mܧ�{Pʀ{��b���;�Hqqq��АtǬz�jG��(�;�t��MsL���2~[�4V��3n��Z�]y���E�M�Iw������� ��+���-�������1�cP����-�q+�n�\"�#�h����a#����Fyy!�1�Ѿ*�S1��SSS���,}�b#�ȉ����׋m�⥒�R�P҇�]�a6N��=%�X�j\��쩹���{����R8���x�8��o��;�ļy�F]gpp'N��#ݍ<Gb�G�?Z�b��I�kK�_�rU4Ih���,c�1�c�1�c� �Z�V����8��BUՇ�~���.��>0&	��������%e���p�}�ԚJ�uP�K�%�������������>���!��X1٢��Zf��;U:�oy/��.���3ܲk��E����Z455!;;YYY�7��\����|�(�D����ă�T�֗��nZy�8!$zL��avā��l�0V%�N�emB>o�������|^��Kzm���"33S�� +꾛���H���.��O4^�e��T�_���`$��������Ĺ0h�0D������� �����?�.��t���w���N:;;QTT�����˙\\.jjj�J&��Te����,�oN1T�$�D'��c�1�c�1Ƙ�x�	�dwM���_��I���h����0$�6�Cm���π���0������l6Q��\AA�����zd?'"�N݉�ˍr�X���z����c/a���q�;���:��,X�3#�sss����`'B�֮�.�l6��А�RՉ(�X��᭖��@�p�-5����%B�b����F�I��[j6�K�\7�>�G����j���"##�P��T�}�d4~�sH�J9z�^��ƥ-���b��ٖ�kB&X;_𥶜�g��`��\��k���©o~Sts�U�.�v�E�Hcc�(��qR��I��j�����N<�S�aNǫ��h�y����x�:��1�c�1�c���Л0�~����}����?ݾ}{/38���EQ������:��q�}h� 	��콇zx۶mg������%A2jY1Ԯ0nL��3��l>U5H����o����G|׬M�ڵk}^���%%%�������T0�(�����%�SD
�R⾾I�o�	��,�힇�>���p;u�e�O����8rw��0��9u~�ٍM-E�ω�ہ��ѴbBRR�+�f3d�t:#vl���l�陸#vww7��{:���K�h������E ����X"�'=��0KB&�?�c��~?��q�ƕ������XS^^~�x��Jflԥ]��J��X����,L������2p��Ij�p/�E%���0��U;�l�F�ن3���?ԃR{,jlҭ�Θ�A;���G�����|�06j��K�P��|b�nl�B�Ձ�W9d�1k���cuюvxϞ�i�JH&�l6?������p���wAB�T�M7j}�X.@����L&����;��A=zt����$$�9�WfGܹ�{K�qB�Kl
p��Ru!��%�t�v���)�YZZ*��RН;��GaV��`���l��1q��('���0�$��i�`��/\"�b�Ñ��x!w�Ӗ��+Pr�(�HiCv��1����"���(��P�L�V��4Ա���V�'B]������!����n�/l�2KbXюC{�m^y�0!w�bb�p�/P����{��.��珻�SN�:���x1�䠻�й�������pr2�K�P�d��I1�E,щܹ�I/�9�;:����rȝI�������v�єt��`L&W��bW�t���8\�!w&��C����	�6W7i��C��+��<�0��E����ų�PyN�$�q���p;����qm>�T8���A���w7`�38�G�������:t��m۶U�1��z�����}0��TBm��>c'����0��F{��XXXx��͛����v�@;Nm��Ȉ6I}��3�10k�[�B��a$Q��џ�?;�<V���k����{NK�$��N��y��!333��n�IOOGcc㸮��B$zN(PK��'e����T�����F Q��H��D��#B�Y�Ewb�k�P]���n�s^�*���yn�8|�֩s�t��frr�!��ԑ���H@�eGG��D<�B�'O���(��B�A�#[�X2�"�b2Ñ���J���5g�[42�����o_�.�|�M����GV��"*0ᠻ�PQ�l�J�v�G����{�n�·ƛWZȞ���v��pȝ���p;I����3�P�}w���g)T���8�!w&
��������;{�ŞC�Ln��|���v�=�ܙ,(�����v�32�;���ܙ,�p���>���`z��P�ҽotX,��i�[��\���<��63�K(H���0���2��(�_�����|3�����z�7BB�CoA0N�A��d�9ߝ���`����߃�+����ǥ�Tlݲ�ox���WTT��������_N����\�}~)�D�Y�B<��R,6�y��fw��c�FD�=Z�V=`���Wro)��9� SMV��݂��~�u����fX���)�N�j
�S��:���vE$��4F�����#��9��)���3�]q3�-�Q�Ss`�K�`��==h��{�FB�s��_T���06/���7ވ����w=��œ�C�dSS�'�:�R��v_&N%�k�\�`�O�-E�$��ܙ,Ɔ�urg2�8ܮ�C�Oh�p�ܙ����=pȝ�bl�]G!w:���;3���v�ܙ,Bn����r�.�FU՛�9r��-[^cRPP@�� 2r����>����LI|2��:(���/z�����===�Iy��J+9L�(D��M��A�`�N��>����^|��ڰ~�:�קLMM��K�)螘h�N���������9�R�a*,��{���L&�yppp1������N���h��1�l9?V��g(��M�������Z�1�X���������.m���b����+�
��$Wԥ�����S/��������N����q�F�c�F���0��(up���hb�"f�QQ�w|�������馛�88�^<IsJ�Or�d�����9+�t��
�Ɂ#=�8�^�a�q畄��,�qȝ��p��C�L���:
��C���|��urg2�n�m9�ɝC�̨���urgF�p�y��_�I�L!}�����śW�^=�e2��j�rH�{�m�����g�#��H�

���ϯ c����%m�R��=]�"�b���N�\���Ȓ�	l���U�Ͽ��֤cI^���Sx��1�QΌ�����Sq0Q�f
��ER�8L����S���n���#�Q�g��k
&�Mt{��.PLphǅ�����+>E���J�[��1'a��������8))	��FAi%̾��1��Ա}`` SA�a�=R������c0�YK��� �.fKY(����f�v�Ư�q�/C�����׿�˶m�u�]�3�>22"�'i� *��;ͫ��zN�*@mmm� �
���e���''�9t�����v[�|X·��1�!wfT���urgF6Q�]�!wfd��urgF6Y�]�!wfT���urgF�p;����%c$�fhh�Am��`� �=����|����o`3��YP�>ѧU�PU�_E1zf���#G���vBR�}/S[S0i���ep�V�3l�jC[Z.\iǟ�ˑ��k�tqV�����:pVWW�->>iiib��.�V���q���]j���S��,h7%�P��Z ��j�G���_h3_D�7h��{�/�Cm0~1��b���FK5�Ώ�p��!��i�1��Kڂ1V��n1.�z;;;E���ݩv!��r�*b6 f�Ge�/�������7[�|1鬇)VRw����Pp��8��`��سg�ςHz-_<FҊ�\<9�cI�$�Ni��F`Aag,N"Cn��`d�V�ȅ%6�E�3��j�]�!wfDS	��8�Όh*�v�ܙM5ܮ�;3����urgFc�p������|ۇ �/=�iӦ0B��*ڱ���G);�-MP˸i�lp�}6�?�),,�Wm��Dd�ND?��6�������X�R̖s!w	���̥ж����o�bK��7��4����+++E�b
T����f�sؚ�bO]��V������D7����i�k�18��Eu�^cg�.0GŋnĊ���R��rE1�HG��'f^�"(?��R�X��$� ��i��!��A�%m�+i̡򲢀>�5;::�F!��jhh��3���^��� F�/�huQd	�s'�kBLV�mUP�S]���ԝw�܎CG_�߿�ClY��k��F�{����O��Ɗ9V�O��)�B۩xr:�Vt�ⴺ��<�ơ�Vb�G�$rgF1�p��B�wwԊ�{���rc�5�p��C��H�n�qȝ�t��:�3��n�]�!wf�	���y��o��vǤ|�h�z����z��(�^��������c�JH����r��Y�r5����=��~)��Ç�}�֭�Oڰ�TXX�ym���zjO7�hzp�j�HW#�Κ4��᭡��+�׍��L¤0�v���]�������(�JJ~�H����t�탃�b�V@�[,�{�8�Z��a�ª��4ؒ�� cSa�O�#m�ژb�ς�IKpKP�ԆU���t �1��Z�6
%��#������
q1k��H64VR�v����3�N�S�%8P�D���a[�N8 sT�Xŀ��T����ZgK��酚��bC�� qӍ(9�y�qlX��+��Btk��B۴Q�$�'SRR�F]�#uf�񑺴�x9�P;iuZq�/U��W��齔=c�(�`,qȝ��L���ȅN�rg�2�p��C��fn��!w�F��;����urg�6�p��C�,Ԍnz��=��KvAR�?�����@QQQ����d52�ͽ`�ß��[=o���k!�$���ۧ�zjϭ��*IO+.


6i���y��,c�X��X�7�Q	�{/
=.<��=��di:��������;�8�iKHH!�pA�E�[��n!#
�Sp���.�k��UA/�p�'�J.��囂ؒ�.��M�%&	&��-P=3}װ#EHñ�!,�;��=X��2��K�m�B 
p��o3	�S�s�S�f:OPX���T4]4�8Z���d�,���ɐ��%6��.b�f�E�1o��{f4����%�ښc��g��,w=.�q	6o��w��"h��;��T<���$��sQ$�WҊ��X9��I�(�Pqڛ�&5�|F�p��{���,�Q���]��M���������3�����/R��k6��^fn�qȝ��l��:�=��s��;��Y��6ܮ�;�ن�urg�b�p�y����9�N�y�q�10D���
��� Iy�xjo���7's��ҳ0_~5�9��v.^���h�����c\.�o�?ʔ�E=ujuc�$cp�BI֥�Q�ݨ�Eb�A�O¦5+a6O��,�-��$m��L����f�l��7�F)lD{��l��(�u�Q�]�g4�5Ք+�N�#{j��.��L��1���í�:!�%
�I�P��9��+�5ؐa��6����Ի�wt��❊g(�%����:�wP�c����4N����=Vghו��FAubV!jٽ�Ac���;3X�(>���x!:��U�=�D�l�|ms�w��#�s����c���"�>}U���z1���]��\r��R���^�C���ti׵zq�7��<�2����+16�g?��YPQ��z,�w.�^�G9�΂h.��:��P��p��C�,�*ܮ�;��
��8�΂���v�V��Zz�ʵ�����߿?ǎC`,H
���.���^x_yl�����h��=v�M� ���ݴiS���Cm����90��Ӄ���J�w�Ú��m��qᭂBd�+�:̈́�KO��&�;;;Ŧ��l"�#�����;u��;��ui���sA���0l�g
*�i�w���?&{4i��X�`l��������;!���8��(�Bf_)��ڰjA�(�
��FAG�
���H{}��S���B{ǎ����f���	G�6�ܕ��kE��(�G��ӵ�#�͚b�����&��m���`��R��\~J��p�� u��ׯƖ-[�|p"T4�ww'T4B�B�џg�
F0���Hڨ ���Lhs�S
*�l��ӡ�C �a1��۶�lq�0�F�;����R9�΂h.��:��`��p��C�,��:ܮ�;����8�΂���v��?�"o����Z����cAPXX�]U�/CbޢCP��f��s�NF��m^��邂�|M; �8�]�����5�(c�7
n:��c����VH�l�y�v4`;�]�x��,��c��(�f/�ѯ�P���;��&�5) ��� 'm�=��ڹ�B� � �������0)4i�m���r�4hFijL9�q�^�n��=5[��3�L[�=V/�	n^�c�BC�&m�ިm�g%�$:��7��%�K��&}����>V�Ax}���2�/}h�;f������|�Z[[q���ddl�m�������+��
y��&f��	gk�<�m��Y�/6���[����{�M]�߼�6m��dh��W֡b񫵱��ċ�'���0���k)̮�� W�Ӎ�vg�,���k�{>F+^�3�`��c~qȝZ���:��`D�]�!w���8�΂!P�v��Y�*ܮ�;4Y�턚���PdCV��|����͛7�������UU� w����3`sC��H�ӧ��-��d9$����~��SO]s뭷��xڄg�v"�$'ND��*E�-e!�Qqp�UC��yjQ�`�NTi�t�z����X=������lP(��JSE�Q�Q
?�U�h�<���^T�$����n���(��~��l�a�Oc�BǗ�#V���ar0xc�PK��gkC2ʑc��X����q}��l̤b z���������h̤N��;�*��p�e5�$�m�u��ٝMB���������@0;�5�U�F$Z&~�Ubsk�o�~���+��4c�\lܸ���S�}4�09mc�\�
~h�z��E/���n}\ԋ��1S/�ԋ&i\���A��6��hs,��_����Eq�2�&����� n�_�9�p��C�,�n�qȝR ��:��@
t�]�!w(���8��E�p���_����|�' 3UU;r�H�-[N�� Ў1Saa!��Abj���`s��M�Cx�|�!�L(�\�x�W�?J��3�'N$���<��Q�OCՎ6x���ٻ�6�����I��#��@H$qPa�jh���
���UJi��2��{C����XvHHdǉ���t���g+$��8�%ߝ����~�$ْ-���d=��u�����>#дq������{���7��,Z�����X�ay��]�����%CD�
�
E��"�aQ%����z�˽�ܭ��;��&��(�d�D�W�6��������r�Z6��ey�K�a����L����tu���2�����X�x%�7$`��?����:,;�1E��_
?,�蓫$�P������d5�H�]N-ZY���~���e*�)G���Çw��<W��s�ܢ�9���뱢)kј�H�g��r%F'�r?�!w�F�
�G0�N��p{C���G0�N��p{C���bn�`ȝ�����/>�z�)P�;^�āREy5N(,,�Q7+..�Al����o��>�w#3�5�K�
����J�`���Ɍ3����������)"����BV�L�;B���OPh����s���"d6�Fo�C�}2�TC��d*6�(m`=rQ��M[|����� !w�Ln�(VdP8��P����,�+�z������}P)������#�n)z��S-����0�B����˱�lʚ�٨K��C��5x�\�%!w�7�~�ru����RѼi,����Dߟ2x�ݤ��J,Y�=�^)Aj�r�OW0|�0��HKK�WTTV���e�l�rP��;��*<��&���!w�.��G0�N�)����ܩ;�2���;u�X��#r���p{C��]�n���0ߚ�?��v�,�юW���g�(6�˙�Ú3�}p�Nr	�W���R�?�/..>dܸq߂�:�Nq�s$\�ڸ��>u��"�3 ZR�7��e��)2�W0
U��i�*��T�L�y�$�蓟�� gذ��6�M>�[��rQ�f#ln��&x+��3z����+`��5VZ/T�&����Hk(EFxr�:$��'���dgp.+ů]�e�j����L��J+<|��7�#,v%�>-���z������{"$�+�����9H�����������~Dj�:d��2�0`� 4p29�g�r��n��f�8�LE��B��t/��[��&9��sL"�<�ܩ�z*���;u���GDB�Of�Ǌg�W'��p{C��z*���;uUO��#r��ru�����Ў�����)�rLII�mb�uq<���$ZN�]�|�Y;CL݇�nf�̂��'(�v��%Y����@�;v�JuA0�LO��$Vo'��a��R����2#)���e��Vm@Zxҍ����fd����	�/6�ga�DE]3*�-T�	�E2j�4T+���2`�s�-���Y���D$#�����@�^�j���P�05�U�יk�ظN����"u������G��\$$$��g�!�M�6acy%��,T�>�	��D�ȃ/o�>雿>⋪?	���c���)�	��A��d�d�Ї���K�F�n��M�mQ]��	�ϖ#��{d���lBf"������| %%6��UYY��*P��~�k'��L�{/��2�_�W�4I��r����p{C��=n��!�3*r����p{C��=n�`ȝ:����2�Y�!w�^���kQ�%�ξngY���`pEaa�� �Y�f6M����%P��a����Q`Wq��u��с�?o޼�G���"EMqq�1���&x����W����N�|H�����U����8�����c}�U�uH�"�lD��#ٯ"�gB5u|*���i*dP(�OL�M!@Ua*~�-�@ShOoHMDȗ&Z*B	h�Z>N�߾����ѶKQ��J��-O�(d���^�b�p���9�Ԥt�D�$�7ms�����J�e� �jB�j I��賠�!�F׀f���>1)1��-S<�!&6M(�46�ai�76�Y|W�@�� ��d4kIhR��e��/7������������k��B�$��\h�ϐ}����9:������ d䙴��ME�	?V�!�n�%墟,������
!9 �)-��A�^B}ed�PRR�8�����Eӡ����K��t�&�)A�����RР�BK_F�=vm){_r��r'Mu?��iW9%���;u����Sg8!���;u�S���ӮrJ�=bC<noe~���)@A_x��`�����u�8~��o�扠���3��ǀ{��a�� ��#�#B�Л�C9RH �⸙dY�K�H1KC.#bz�" QO��Y5;�i%�j�=2B���:�.koNk{	̞�,�1d.A���U%�PS[V��X�p�F�;5%�h���E3���HBB�@�	�/�@&�ĉ��~r�e��8X~f����P�mI��5���o�`l�!M�:�f_�BN�d����Q�0�N�p{C�+�n�`ȝv���������f1�N;�p{��{Fo������#r���Z��f��_��.���s���G�7�킹s����eY�����a.��~�G���S�_us��U.u�h�/^����Ç;�̗K���'!9�*	`�X
s֗ ��h~$�_C5B�0���MQ5���_�\AQ�j���l4˾2��hS��Y_F/2�x�-��Ҁ\�B��	�;!^�r�u�/%��j����C�3N�G0�N��p{C��N�Gȳ�c[+�3�N���p{C�3N�G0�N;��p{+���`�z
����ɖe�3{��C'L�P��9sf�,��(�Dx�,&��S���.Q"+��0��߁���kjjf��� ځ������]��
�Пy؞IIDѣ%g )i$BUk�W����E�Ok�܁��
"������p�F�+��2��E�&�5֔�ۉ�F���	��/`�Wr� Q�1�N���p{C�#N�G0�N;��p{C�#N�G0�N���p{C�=^��L�3�w���tUU�[TTt�����h���߲���L�G�I+�Ⅰ�`�=���:v_ б%��Nt.Ǌͳ���Ɛ;m�8a%���Įg�䖓U�烈b@V(��kW@m*��\������ ����T(N�D�\V(�Qw��Y}��y��	��k��l�J�6�x����f����zC�-���#r���!���;�����ܩ=n	�G0�N�rK�="r2�?B�!���sau�~��LEQޟ={��	&, Q;d�]l���1��P3�� E�Qdm� �נ2<d�h)3g�<qҤIM �Bqq�8˲>��IÄ��d"�-5���>{@�وP�X���R4����O˳��D^��H�5��Bq�*�aw�Ú�I��O�53
���<CN���_j�]��pI���KNƕǔ����1�Nn�G0�N[rS�=�!wڒ����Ӗ�n�`ȝ"�n��!�3r'�O�=�x�(��A�{�`/UU�(**:r���A��ŋ'TWW� vO��o�T��}��0�eƛ3�8JN<�贴��,Xp�ȑ#���b�����-�zG�z�,��6��_z��l���A��U7Mu��Ĺ?��r'�
������*Ŗ�Ŗh���1��ş "�RIH�;���*V�5�hW�	�H}���
"r��ɭ����Irc�=�!w��n�`ȝ$���#r'���#r�x�Kֆu0?|گ��C�E���ٳ��0a�� �Ν�R]]���=^RQ���@�ŤO���a�x��.������^0<����׊����,�U���\Z��0�~DԳd�@V_���n�u��H;'Ú2�.�lDqAN�H˅���IA�a2�)�X-�SsT�vH�I}F@�݄P�ZN
��R4��+���,9����r5�a�=�=���{|ss�=B��O��ǳ�c�����7n�G0���n�`�=~�=���{���p{��Ƌ�~9Hτ�d���aII��cǎ���͛��e�܉���G�l0E�1`~5��G@1
s�h_��h1 �ť`0x�eY�����ܣ��XՏ�)_ 	y���,@X��+A�--1��>b��x�yRPz~K_YWq��-��D{<��\�%9)(=���k6 \���?Ħ�'W �g���T�CU"Wΐ{��J�=�!���p{D�8�>�bC�q������W�������#r�?�n�56@�1/�M5MS�=����)P\***
���{�c������P�y.��Hb0����������H1 };{��c'L�P��e)�D��{<��.�����G����'�����1�kl'ښ]m6w |2�^������l�_j6�vhٟ�2�C��eUw�~A��C���k����㋗����/��#r�/^�G0�?�n�`�=~�}�����0�;�	�hO����ƍ�HQKq���h����%v{�kB!��gg�)�p��ue0^����A���Ҵ���7@����_'���<.���Er�������M��޻�l�C�j-��P��RZ��I� ���@�=)�n�ÛF}+��!՟�lOɶ+W���IA9���I�f=�������*(2�.'��}"r/�ܽϫ���������/��#r�^�G0��}^�G0��}�o�x�A�{�'Ӊ���`�̙3ϙ4iR�󊊊�(�����B��ga�_��c�x����2h(<(E��Āt˲e��1u�To�$̞=���i�Z�5e�x
(�/��ci�8I��� u����Ă�0C�W�gx3N�@����%g��v�^�"o��>v_�*��AMH��Jۉ:FV�d�����u��� ���M��Kσ/-��v"a�ݻ�n�`��ۼn�`��ۼn�`��ۼn�`�ݻ�n�`�ݻno�ڸ���@�v�HQ�iiii#g͚5e�}�]�3fh��J���=�q�+��|�MP�0�K����=�_;]��=�����&:������S'N�X�`08Il^�,+e-�	�����d�����$}��7�;v��A03z1��Q�|�9�����ѮS|��*�?�M�M�_r��W��N�h�ٕ����O�E�f#��0��[Z&��/%����<�!wp{C�����ܽ)������Mg3���n�`��{�%�����0ܾ}ƇoA�� (�G���h�VWXX�_��̚5+G�}���ë�����]�Ū�b����-����P�:^�(ʑ�@����䤱c�A�'gX2�b�xt��d����SH�fJ�f�����z�&�5Hr9YM՗�k�~�K�-�k) ��@V�WV \+����{)�
_j6'u'��ה<1���Xr7N"�/�{G���#r��x
�G0��-�n��gǵVrg����-��rW�FFrw�x�G0����iB�^��}��l�3G�����U�ƍ�YQ�<@�=�������k�Ply�7t2c�SPF�e�`x��4�)**�a����O�:5��%z��ٳ�k���eY�㌗����D�2��(��"�ʛzC5�=쪚iyv`��Qt�PtZ���P�=)H�-��Orf��刾2���(
Zr�ݬp3�r�\�U:\CN�}�_���Q|a����5����7�c�=�!wo��p{C����������!w���p{C���p{�X�V�x�h'�	�D������o�������o5ȕ,�R������-��aVY)�W��?��v��{oi�q��kۧ(�5�>|֬Y����A�RTT4E�R6<Κ?�^]���IKJ��?�d����9�GD=G$#�;~��{��/�a�~��GQ5�R��	jB
�(v��I �/���sJ�_q�s:ENLHʰ�J�^ ��5���+�����[<��#rw�x�G0��n�n�`�ݽ�=����{1ܾk�w_���X�#���M��|���������())yZ�z�`.Z���@�ǀ{��:d%wm�9�:EQ~�iZqQQ�E�Ǐ�xbʵ,�񷛆xP[���rj���d��@v?;�d�7�2�d�W�RqSZr�]�]��>"�Yr�Id��{m9t�WrbP��AM51�%�Ε-�z�+`Ȫ�z}�}nɉA=O���W��cQC���p��rw'��Ɛ�;1��3��݉���1��>�o�!w�a��L���#p���H��e��\0<"
]<q��
��Y������!��E�DП{V)�:��{����PF���O!�@��(O��������"�#���ߊ�}�8�?r�*�#���cKUw���X�R}��J����O��R��%g�Ո��y��9����T�R�]����P�h��v_)Új9������m73��v�-�Ġ�Ye?��f��DD�Ð�{0�޾H��������c��-��݅���rw���ǐ�{0��>��݃��.�(�����]t%��i�@�Ȣ����x�s��ϐ�����a��� ̏���{�ȍG�z�}@Z:�eYi�6'^U[[{��I�t�#̙3g�����#G�OރY�-�(��V��2t��0Dk�a���ٕړ�j'r)51�r��}��+u���^v����ډ\J$!�@f��������KVv�~���sJ�ډhWɐ����x�!w�b�}�d����Ux$�?C��p��ɐ���~�!wGc�}�rw��w�!w�c�}�ZB�x2{ C��p{יE_���#h�M�8_�m-�z~aaa)����oY�����/q1~���T�x�;�K=��&�F�M�5nN��E�=--����Ǐ���̝;7%_aƥb ��AH�ˇ��>
"�E����c7y�j��dཾ���NR�	�Ӡ&�×�aO( �ğΉ�'�Lq���i���(�o�� J���G��-�8ȵ|~(� �Hax/��d�։A��+�,��Z{� {"%�!���dI��ʾR��3_oD��1��X�wL��̐��1ܾs��;��;'���^'�#T�$e������a�ݹn�A�F������c>��a{@��q�עR\\|�eY�6�z��;)��E�xb��w��*P�b���9E0^ڔSgF��￢#�Xl�2v��@1#E<�'���[�Ł�3V}�;o B|SHD۱e()��p7k[�IMu�X�vH3!ZR�����GN���
����!z������\'�N�k��%����Wf���_ʠ� �yN�--�^%�l�+�W6����W�$C�+ ��R�c�!T"�F2����՘/���c�c���z�ε��K�EJ6�9���P���;"r�(5���$��qH}9�]wJF)S��F�,V�r���H�L��ɐ�*��R��Q��|��;D��O��%���c�x��'-w�����#p�@r
�H�eY��s����,,,|FQ���М9s��q��;�q�x�iX��z�a��"�!�A3�Ft���6����a��QJkAQ%��#JJJ���w�I�	��`��FD����Kϳ/�U8e I�9�U8M=�x�h~h��-�4�6�"�_����09HN
���8q�}eBrK_� �ʄ�4��\�!���2�RN���\E(+�ۓ��+Ŗ+ZQ�稲�U��	��@�V2�~L�z���R�Dn6���nDn58�`7"�ZW��;��˕���R_EQ�*..>����������������0�l���;f�o�rܝ�5p�\�^}��e] ���I�̈́	�_�n�����eX��rQWD�p"��C0C��5�N3���Ū�}UK�f;|��b�6���G���,@6�����OF�K���M�
r��9R�^N��d_��,�hGu��76�l�'�9��>S���>'��[���RN&'�m�,���j��e1mi?EQ>*..�Z�_5nܸOA�*��e��_(�񻴋�P���b3�pw����7���@ n1 �+��D����4��o��V�:Ͳ,������\\��`�d~��� "�n�j�&[r���,��"��Ko�C�r��0����`�>v�]�Z�G2|ED����:�)E���ɰ��'M�O��ҡaN����vp]�}f$��O�G"�.�+�����!�e��W6ړ+7�����'��[�-[�I��������������c����:d�Qc�,˚(6�}"�7�?�#P�����\$��s���1����� ��'�c�.���]���x�Z�*�e>��/bPzIt��O�0�;P�-X� ���xJqq���^ X��`���bQ,�ʔZb�ݶeW|�8e@���p��*��n
��0&T�����}�hW};�Ɋ�Ds�9[YF����Lڪ�G���~�#��+[�IU�3V&�}��I�ې�*�Hںܢ���IC��H�gʉ=r����G�L 
p�$Qw0M����_�x�(�d����Larr�#G��:���h�x/�S�s��e�x�Xe� g���@�7��(���i �Eg:M61(}*:�G233_>|x3�]%%%M�<����lq��Em�[��WJ "r�H�w�~�RK8�hٷZ���k$�d��&�E�V��T�u_k	`�aMDDnc�e�߄����
ƛ�J���Gn�Wʾ��}����W�+�!s{՝��8��-e�h�KZ[�����}>�:���U)������JN�!"""""""""�-;�t|��JJ*�Ey����Ƣ��G��ㅅ�L(o��ŋ���~#�'Y��`�fƌ�`��
�<�;���P�s��+�f�������*1(��4���c��aƌ����'��4������a��_oWp'"r;T�,b����}v�22�DD�.9�GN��J""""""""""7�֬�q�����o(~��ު��(׈�U��Ų���b�����0�`p�9����,�<偶b~�_o�r&�`L�A�����Jfk��\�� ��}>�scƌY�8"~oU���oE;Y�|P[����`-�DDDDDDDDDDDDDDDDDDne.�<4��/�j�[S-�:Tle�,..~Gl_�}oa�`08@ld�\�+��.s^1���9�Nf���	�kn��w �]{�X�a\#:��b��4�?~�|x���Š{��=���qgU턽��W3ADDDDDDDDDDDDDDDDD�v�7��ѻ�)��ڕeY���V��`�UEQ�jnn�|�ĉ�� �;�%~�_��z�؎�U�����4@�ŀ��Y�u�o��%䞝ڡ	�s� �[D��J�/:�D�9f̘*�Tqq��.v%��'�:���}.!BDDDDDDDDDDDDDDDDD�b����|�ڡ|�γ,�@ �X\\����.��oaa�p�y��e���I2�..)Z?EQ .�v�|·^46���w�6m�~�?����P�3@�_t���\�0�`0�����i�_���bpZ
�9sfbjj�8UU'�����h���	�ןA�~y�eA�n����{ �C�Z�ɪ���kѾ4M������I�&5��������Qf
�We�P(���W@���
��*�A�ǀ�KXe�ZB�����T�.QE%�Q�s���BN�b3_��E�����-�{�׈���4&dOOO,����^�1G��l�D�q&Uט�o�?0]� """""""""""""""""�ӄ~߭�P�L �<ю�MUU�����`p�����(sMӜ/�_\SS�<�w˲��s���;T��h��%��-]Vh�.��C�� ��@�����X+�������o 1	�%����M���݊���� �R\�B����^엋}9eG�*��)t]���C�5)�Z�/K�g�]Y}=G�O���/���v�����s��~�b��,vy��C��F�.��Q���D�iG�fY�T�����4YPw���\\^!چH�P��*�U��V�;0M������>!M��|��z�[��b�ۚ)�'��P�kl@���Z�������G�o��+�]Y"���b7ٶ���^EuM��\��m����G��x!���+����o��˯�:b(*dA��b;q�`d{�A�1���^��먛�B�v-�e�A��Y�~�~��]�O  �����45������������������(n���O���]e�� "د������q>�}pw)s^1���i/-��d�39 �o���DDDDDDDDDDDDDDDDD����J�/�
ʨ}@Ϭ�Fӯ��`.ȝpw1���ŀ����@j���]�]7�K�ŭ�&����e� �GV}�[����G�{1��r��_w9|W� %3D�������:�������������������#|׍�9�	��(��T���*�+��܍w��J���
������x`~5��w�DDDDDDDDDDDDDDDDDD�Jס�s|���/Q\(߄ЍW��@�ǀ�GXk����.���! �2�÷`<�`� """""""""""""""""�m�&�q=�)���ˬ�+��rP���{�U�	��.��¿C�{�<G�t=� ̏��e�x�yX����g@cd��ǚ��w�4ԃ�����45"|۵��'����WX��6��"Qǘ3?��i#|�;��"�0?��c���ܽ�4�?~�5���z6�� r39�P��ZX+��������������������v��}	�����^����ZW'����w3>xVu|��$�ȍ�%?A��;�NDDDDDDDDDDDDDDDDDD�c�Z�п.��⫠"7��a<|'�Y_���w�3���K�I��Dnb~�)���B!QU�øN��C���X�ʠ�y�=Y����8`�Y�����ǋ���"���aO= s� """""""""""""""""��c��֢�;�  �әsf�x�vX�u �c�=^46@��Fh��m�逪�ȑ*ʡ��oXK������������������������W���@��"G�,�
c�S�5A��x"_�o�b/͠��(� rkn1���ր��������������������Z���C��eP�"'���`<8�bP|a�=��a]�gh�\u�x�8��ͫ��x�5ΰ""""""""""""""""""�!����WC;�X�'�	��QO��ρ���*�A��8%g��_mґ�~H QO�V�¸�V�+��������������������z�e���M��ρ�ˡ�������>}�O���W���(f��7��<��ADDDDDDDDDDDDDDDDDD=�*+E�ꋡ�r�ÏD�"�?�>�%�	-���K�z:�#�TD�d�o���=0��������������������DV�~�!X���Å@v���4`�������?"ܩE(��G�|�	|����a �v����=45����������������������.��e�B;�hG���s)*�������E �`���b�\��՗���hS�~?�����LB��Z�=���������������������`����o�;�B(���[ȕޚa7�:��Ā;�%�zx���o��I�c�:����A������������������ȵ�����B�ǝ��>�O������sׯQ{���vYkˠ��
��ӡd�hW�%��?���DDDDDDDDDDDDDDDDDD�^�ة�ʳ0���i�B�{�vIE9�����′@�=�ӎ����������)-3�툜a<�0�� """"""""""""""""""�֬F�������ߟ��@�P(�÷`��"����a��:&���a|�!|'�u�I���hKV}̷_����������������'���H��?6fYh\��}��M����Q{cȵ�n�v���p2,=��H�c$
N=��,T}1�_~6���|���ǿ mL!��:lx�E����}��l���EH9ZRrT���^yU�����1��������+n�5Eߢ+��T�9�<�칗��+{���������<&'���=�M�K��/g�ڲ��?^(�����.�B�a�;�cӻ�w�>��r/���������}]��}���sҼv�<z��v~%dN�_p)��kB������&4�Z������O?��ꊊ�C����y�$���ڹ^]���?��',���}���2dO:|������]�(�����<h2��:�{�q�/����SU�:�4dN<P�i�n��#�q�8���/��8�[<�'������͋�C�5���s�y��N���9���=����^���Xu�-��_�ه���g<�ڒ�]�O--�λi{��V�����hZ��y�/�IC�����״j����+:#i�p����n65�?�$�M�
�8�O;��|T�ֿ�d�ǎa7ݍ��{�;��Umڀƥ�Q��Gh��P|���������C�z �C�m�sf�xJ�#�s3��b��v�\�ۡ~���N��۞ ���̏߅.gW�ׁ����������'eL�%RF���c��;|����ծ��Obޑ�#~ݥ�f�>����P�-H�I�V�xbe�{�@����/gx~ll���551	{��.�����/簣��o���o�ҩ�H�}O��{{�?�ߥ���z�-�q�,Ѳ=
�lO��U��a��/ٯ��PAm��w�'^F��cc�x�Κt8����;u2@���X���pWU��������W�u�;�scGr
F���G�Rf��	�;���w�Egwz2�����;ᤘ=^�ă��%W\ة�O��o��p�8V�>����AW^�޿�yRO�1S0�q��[ҩ�z�m�9T��O9���BS�rēAW\kacE�q�{��O�ѩ�����c�]���v���\t���͗s�q����pg�s�O�jO��틬����D�v�s2���~.c��o�aމG��l�.������uyǞhO��,9iyԋ��-�ٓ���[��K:uI����g��K~B��Q)'ɑ���O߇Q���O�6�(���0�}���x�IX��hW1�N�b.��ڿ�,1"��;�f@��0����_�U?��""""""""""�V ����Xq�?�r���oW��οds�}�}N����rD��ln��u���#��cbn�LQ���+:pߙ�_NF⠡hZ��Sߟ��6��#d�W�Oe��]%�Ǯ��i�2�;0f��-���˱��G���E{d�+}�~���!Cz[��%�RC���F��v���~"���-��}�'_��S��QW��vbn��;~*����;�W�\I%�7��|�N}�\1@�;lI�[�;����i�|	���$�����z�M|��_ui�7��(���łܦ���ys����$@Y����;��rrP�s.��:9)����v)�.�s"����+�2�K�a��$���W^�h(8����N������7��#d_���;:ʏ��a�c����W(Y��?C��Ł��<��W���Dh���A�8e-�	ƛ/�,���b����^bD4;�~�P�C����`���N.�DDDDDDDDDD�5��E�eHHVѭ-�ݩ�Oj�����Dq},�ه���2�)�JfS#�g��>=�y������w.�WV�]~��;��I���{}��᝺?n>(z�
�d�˗��p�ƨ�����t�}{�pRg��\�Z��=����c��GO�c��{G%�.�~x�Ou��O<Ğ���!����X'��!�ފ���.Xߓ��q�������Tp�X����̔8`�mTJ���	�~�}��C@���u2��9� T}�Y�����vZ�="����;X��SѼ�'*�a<��w_�z�I�>\�I���U+`����_uz2Q��-��UA?ڱSt�(+���0ޚ�`;�6j�\�JVq�l�}{�&Y�2����a���@���~���Q;�(:��V�SNƪ{n�^U��߼��^'���v0N�`4�͟�r,�8X)W�V�]�U�e8��tŮ�v=�����8�&Y%����a�B��eK�J�ZjZL�h�G���Q�����4ݩ�S�w�:;i�U=���*㱔��C�UR�J���d�T���+Rǒ�꾏޹���U,6��ڮ��Ή}]�O)�vƻ�v��M����s;p���u�%'�x��?�(Vr�3�877�����B�xp�������`��2��7�S�a�������ٔ�GB;�X;��S3��5����q��*��M """""""""��U|�>�<�`T#��_!�� �U��a��U�dЌ��U�9ֿ�4z�tZ�3�a�_׹��%���p�G�COkZ�R��WbЕ��-�{5,Z�U�OG��/�Y [������>����Գ��?W���~D�]7���]�n5�hђS�4lw���=�L��]s9��x'Ԅ��<�/��
��UQ}9a�S�nf��`�U�b�w@MJ��c��3..�r"ג\��n fϱe�Xy���[���s�:pw���F c��`�������>�b��˙X��Q}��&ف�ƥ�O�{�����s~��k�֯���0_z���\!b<���@���sa|��(O��Ā;E����)��@=�h����l\�7a��hn�����V4.]Խw���R�usKm�*_��gb����M�&���>+n�'hk2X���:jh�;�
�ء�mɪ�k���մ��_}�j��6�>����i�g<���B��#��w�9V���0��u��{oC�G�!m�x��v^�U����/m�������>V󺵨��Q��!'i���������q'��3�0��t7�m��ed"lz�u��-FƄ����������=�g[rR�^��+�U����K{�M�e��@��1�?.@O+�M��N��=y���:�d���}�Y���~�9G ��������9��v_�k�yᝬ�WW�z���jі2r4��N���F�w�T�a���K}�t�r6�Z�=|��׽w*�ׅ֮�'�E=|�(�}�9���S����]���K�@z�~�;��������>�(q��.(>Y�U0^{ƻ�A�ԣN�һ/�]��4k�v�v�eE�]p���g_=��7^�:��DC^/���&��������o��)���X��M��gQ4�m���4EE��PS�-ܬ�o�a�}�a���-�:t��'��āCдrhkr�DG&O��ڻ��{M��N��هe��@��;�/��]���v��n7இwk)�ȟr
�>�� \Q.�7Q�o�i;�bT��	�):�������{�)ǭ�R������	�1\����y�!@;�x[�^�v7�1�C_+W�i/��Q�p>�D�Fീ�\1b�U7n�2�<W���Xv�e��%�P���p��㦢��@�����0ߞ<�����?hO�jπ������c�x�����a|�!�q��z�PG���1�m��`~�_�>�'+E�5U0�|	��_���hhN�:� Vuw���3a|�]��(V�赛@DDDDDDD�f����ņ�r,�:�{�1���ƚV��N�.뗇`�3�ǋ>g�瘀;Qgȕ�=�(,� ��3�V�"4�Y�����߱X� V��'Rm+u�������5��({�nx�������a��_F������C��Ѩ�?D��Y��ݔ�\��u�QPX@�9t�.�k~�)��X,�b�w�-Y|�w�ES�{���t�~@�g/��l3?���s """"""""""r�>g��_x����'A�@��L;��((>�����ڹ� r�����uȑ���]���{�|V�{��J�4��L���_�
e;��jB"�{
���5O<`gw�F�NK�v�y�+{e�me|�ԆU�	�ۯ�x�5����z�P��q�	��0d��/?jk@���c�T�x�5�)}@�� ��8J�~�(����s֗0���(���[�)?�'�M��2u\B��<�PT~�!�.���:�u�������z�~.j/�#�ܪ���0�N�Vp��X���0C!�U���ê{o�Q_"�	� �c����E�kV�����{��mnK�}Om���>��nJJ*�����
�˰{�m\�d�/>��|	�z_��VY)�מ�[$���xW������|��
�
����%��I>��hQ[K~�?+���6��*����]��C_������G�g��������E�볏8	���ym��l{�pz�~H=u���ɶw�󋜣O���_��m�8��ґ����9ZӪ�P|>��w[}���g�R휢v���|u�U_�O���Va��c� ��kw�6m�Y���+�~Z "'᫜g��{~�Qc��4���������Ü3V�,{�'""""""""""��B!��i�;��6��O����P�p>�*u�}���xp!����{��'B��}�	[R4
N=+o�DN��'E6jbb��
��K.� DNV����������������U��fO�cd���0��a�ȑ�^z/���M)#G#M�+�ς���^���Ѯ�*잘e��Pƌ��� ;�A�k�O0e�����Z����X���Y����}@490AL�>�P�k��i�s��a�-�U�����ɰN��/�+�oK�y�\q!�*�Cw��'c9�ΞӸb)�����<��m�S�a���a4ԃȩ��
��j���ks[�Qǡt��["�2M�|b�׶�)y�Ș0ճ��ӭ{�Q��6�'�����'s9ՆϢߟ/�����ާ��ـ�����6�_�v���h|�h��@8�ޅPF��:l��X얬�ka}_bg
�s��&�_��r`���^�zR��u�nPv���{���W���XK��i�E?�������������;��P����;~j��r�>��߀���p"4jO�EH�[��e8)i�04.[�O?�n�ݗ����b�sO����>�0�(�V�+>?
N9�w�DN�������K�
���}�p'W����pɕ��䵹M�����5�����(��mn˞�+$���U+AD�`YvrCV"�%@�A0��#[r�{��9�,ӄ�f5�E`-Zk���6m �1�N�U]i/�a�Ē�����bTJA{�r;{����V��r)�%?�*[�
�DDDDDDDDDDq@����ˢ/�N>��N�/@ʈQ�޶��0䚛�kgY��_Nf�݃�����E��ۈ6��>��{�)�Cx"�jX�#����8��m�N>��fc��ʨ�Æ�_���m�	iI���q�R9�
a��O������-}�/�:jo�͟"���
���m��+���ߝ�7�^�K�l�z��DQc谖/�!>xӞ����e���La�A-�T���]ז�d
K��Z�̥�X��<���_��1�Kh,����'�-�lr���e7�w��ظ�������c���M """""""""��T����)����ks[�S�@�#��lrև�v��m*KV8���}j�s������C��ɇ@�#�����6�'"��Q��G r29٨���/#y�L��π���1\p�Yv�r+b�.��,��J9ݺ�@��/�����6y/��B9U��e��b&������Ӱ���0jk�%)��h�z��BF%+��.�ۖ��������(^�-���l8���hg
-��Y��%�.s�e�w�uy��m���	�l�R�3��������r��4�i�־].O��Ե�A.�!O@�jE��%��USK���g]� �����������h[2��^�ݟ�c�7��<�$��C۽�z�WvYro/��V�h�)0�A޲��p��ۭ����sp'ǓǨ�p-+]o�����������hͫK��8{�mn˟r
V�}��*���Z��M(��vW7�=���~���h������ZJ*�O8�~���w�>�vok�&hL���vÜ��o������
���B��j������}�+�fE�]&��v������-[T��d	e�\������b���=0�f-[���ƶ_(��'$�JL���{�^E��}���CB
%����ņbw-��(H�(6,��]]�kD)V\]l((�E�I�齿���y�$9ɜ���ry9�sf'��3��{>2�/���]��0�KM�/��_X�����1�R&`_R,        #o�'*O߬�N�m5�~w�k�������s�c-o��sޢ�����u���{�)��}&��ʀ�p�a�����٣�JV��Z�sl�Wuн��L�=�~�����`�S�=0�����W��?	Ih總�d�L �)���+��&k n��͗*]�J���R����5�}�?�|��քl'y_}!����T�-]�����,�QV�Pa�6�F���9̊v����VV쪕�z�)j=��jx������p�cB���RI���O       ��ƄLء�]�j�zX�o�L��taw��pW��:/W�+~Q����߷?w?��ƫj?���j)�Fk������L���g��C��W�����B��a��`�	�U�Ǫ�I)��u�c�2+C�]%���p����%_q��M~ƚX����;��'l��:�)��������e�yh���J<̱n&|�H�?hh�[2���!�        ��ߞ�N7�W�Y{/��Ƹ&��@���V�|˦��������Β�K�?�ٙ����J<�[-�K���jg� ��-+U�{��~��Zܩg(���T��7nfB�]�d������U��ȗ��a"?R?𸂢�m���*����2�Ov��nщ�������;J7Q��mm5�:��A��
�����[�fD��ԫG��!�����<o�� �w        �*t{�E�VT��jkT�j�6?��*�o��Ԕ+{ΛV�սş>�
�mX����L��y�����_}nuB�[hj{��z��֯�O���J�b����	n���+�y�t'�[��#������L�3u�j��l�u���p����D�]9s���{��d��`�+�J�j��Uhr�=50,����zޗ�Y�U��r��Ě8���V3�8���R�q��!?����?~P]�J׬���=�+��M�
YoNW�����>IQG��忨%u�U����.2��   �w        �*�&�����;���z���Y˧���j_�;�� �(��`�v>����
W:��rπ{��e�ܑ��vɶ�Ɵ6����*^�~^��c{�j)W��)��?hAf�S��(��l�v�L[�~D�y���z���/Lw����*sYP���RY�����l53���>Nſ.UKJ2\���&�o]M������<�̙S��l����{R_|��������x\x�A�>����tU�씛dΜ���nR@��Ob����5V��L.Z7��{ ��A�        `/�[h|�������&[�XA�αՒ.��g����<���3:n7���ן��XW����T�K�׷�����o��N���D%�w�v�yS���1�p7�ӓ/�m/Mj��a&d��<C�1�j.�ݬ~xG�ij?��N���h���Ւ���~7����3�C��3���
����Lw�0�*'	�\��S�&�ٙ���%^8�VK��k�\eV��E]u���zm�w� ��         ��2n�9}�c�=0���/�Jۦ�[-%��3��P~]M�}��/�1��((2J5%ł���l�5Y#�c���~��&���	p����x�ϊ:�X[-����󪫪����r��n�-/���|��d�������	�\�-OtPE�6�sM�������9o*u�h[-�o�9���6��|ߕb�����!J�b��'�S����D�[6 �A�        `/&�]����y]%��P�aG�j)W����/Y�[pl���9ޱf�N���z�&ı���Şt�r?�X�?��9�5u�p��ѭ�bO<���Y����c�	E�I)J<�"�����t���;@��IMW��+��}�jw��/݀=�+y�my�a���E�r��&��!ښ�Ғ�}4-���+AA{<�:�s]�񁻄Vά��B�Q��e*Z����;�VK��kE3���{ŞS���!�2c�  ��        vc��nz�~���Mne�<]�d��������ι�7�k��;�
�����u�����ӻ����p�c�o���7�EA��Z�5c�&�w�j{����J��ߝ��U�����(�/�(4%�VK~���m�v��m�y�ֹx��RŶt����%�)愓m���C�텧USZ����XaȄs/��!(*Zo�]&�&��"��H鴺�Y�`ˤ�:?O-%��>:�շ���f�:	MN�A�?���SU�~���j����GT��R�U�k����m����oϐ�Mm���>�U�  ���;        hҟ}\e���cj�JU�r��vf��r��Q���($1�VKqC�����鸽���T]X����/��1����]]e���c�Ď��Vʐ�Z|��jspW�m\/_�|�p��G���/�U�{>�
��L��zs�:�z��y����u�
\���+i:���~h�������h&X�p��U��/S��ij	֊nԆ{�Y�"���Hk�Nc�p�D���A���TS\$�3����m<߽Wk��g�RB{r�F�ǌes͔t�Z9�b/�E������Z���1�������L���Df&j�uL��̤��wf�����\��䀞c�Mbz�Q�9�|��cVjJ8�"�|� P�        �U(��.�^����RY�����l��#�V���8����j�)�k���������LW䈮�U�n���Lp&�a�.�J�j�~h�|��ϐ6��=7��X�V\y��2g������2�4o�� &��G�����.�L�[6)<���f�p��ZC��j)�*O�|��+]�Je���)3wM�ۍ9��9�Ub���8V��
Ev���r�(m�EkR�?0�7�n�C���֬h�b�=���u55�d��w�o��{���OW�7_6��*^�T9�|x��3��-�աOOV�1��6n�r>���� �zp        �A������[f��PZsܣ�;A�q���'&�V��Ma�l���p�c�7*o��{~�{Kt�ҟyL���E��IV併9�P�T��j��*鲫l����X�a\��V�o��.���;����}6D����"���l5�N��mӧ��#�l��
 	g_��s��_�$%�%�����q��������7Fe�v��g�|�}Ey��ީ�5)���D  �w         T��S9��v����<�
o���C|����M���-�����E�|�P�~������W��)����6J��m�y���@��f������.ў�uʐ���_�Y������c��#_�l��;ܝ& ���̝����QHb���~�~p7��_j����?o[+�-�3��n*۰N����\��ߠc>Z���[���p ԋ�;        ���>�E����}+�k�c6��s(U��������:n�>����Є>��LGJ��?���Z����xm�ꪫ�U��5*�n�bO�k������=���BnUSRl��S�_g��q٣�JV��O��Z���Je͞��7O��"{��c{7��F�R��{�?���2����+�{n���$��Kz�6��N�3�9w��J8�[���] @}�        ��ҵ��p�w�9�d[�˷>�����S|D��^}���2��bO��ys��9�U����)�j;�\�|�� 7˘>�1���K����n����Jz��*f��{�	p��Y��~�-
���o�̈́����ֱ�:�k�^�����Q��L��S�7*o��+c�	�[�������k�~\�pIJ  �!�        ��2�Oq����&���+^=�S�I�߷?w?������ֻ��h��^3��;\/�/T�q�c7��a��~�b[�����ϳ�/�-O�C��U��T�G��%�m��g�kM�����i����u�ה�Z[���}�ӽU`xk�����טϥ���x P�         >�,�^�e��Ӻ�j�îU�̩^=~|�3���8��� �U����Je���:\��}L/E}� W�2g����{�V
��I����vf%��{`h���f�����/Z<�k�ݘ�	R����'��
�]���+٣���r�H��~A����ֹ��g  '�        |Ym����ćl�𴃼�a=�M�bz�,o
m���Ck���p�̙��~�M
	��R��VŶ-�,����4�N���j���(���Y��U��Ey���2d����,��L���U쉧�jɗ]�������;��l�C�R�p�� �5!�        ��ߝ�N�ܮ��[-��1^;nܩ�&o�?} w?W����O>P⅃l��s.P�G��f��e�~g�ڏ��V���G���]�W���gl�C�x�E|A��)����h%]2X���������s�mg��q�|M��s礦�X  ԇ�;        ���))V�{���&�S[Y����฽��*\���/�{OE}�m{�i�m�˘>�1���t��0]WS�������%����}u�p�B�l���/�r|��-����Vc���}[�[o���l�ȞGy��[�t�rG�  �w         ?`��)W�R@P����P\��ίe��z���eL����9�����RpL���U��-����>�V���XE�6���X	��'d0��Lp2s�k֪0{c�g��Z��L|�Vb����~�M��՗ưY�+��k� @}�        ���m�ʛ���<�Y���(�&��uu�[�y��i����y
���c��{�i�����35�0c�)����Y��a�X+����wgY5��c��������?jw�e�eo��|�葿h�  �w         ?a���p��7�q{��e���h�>�jj��͗J<�[-�� �@T�u��:�	�Ef�N�Ku�q|QUn�v��=%�R���))�B�ï��2^�����#oT��7;�j�
U��� �>�        �D��T��WEq�׏���{ނ��߼�������_f�C��i�|���wP��X��/���Ϸȱ������)+U]U��:dL{II�^����(s.Nz������U�U������G�"�m���?Q���(���_��)�VmE�  �w        �*t{�Ŧ����j��[��/�K%+��2�xE]}ƫ�ILRTϣky�?mԾ�~�:����?c�cFv��hBSR�v�]�<�h�������:n��I��[\�*��k��oY?n���u�y��""�z��α���n�>�t=T'������i읊>��������
���?c�2+C���U�����Z���O>T�	�Y���}�	��Ú&�o]u�
�[���o�*�Ɯ[;\w��N=C�m�}|Pt�����������||󥶾�j����J׭V��o��T�Ǽǝ<�u��]����j.�e�j-�C�~ԍ��w�u-U�}�z��j�*��VW��_k�O���D-�\ߘ���Z��琇�RMYY���s�Q�q��M~VE��(7�xmJ��ͽ��ij۬U�  ��       @������w9Dq��������+��vΝ����(�]�׎߷�cW�ʌ�~�T��GǮq}����	I9��F�cM�-�S�zgcB���q�xm�Z�;漩��Fz��ס��X��^@H�zNO�����6���Tm~�A�4Ϝ5Mi�0�������s�i���ά���>��ξ���	K�P��<cج������jW�*a��pO��~��V�̈́X[��xLI��l�~���$��#u�Zu� W�'2�O&���do\����W]슐{��OT��y���|����v�(��xr �op        h$Ӂ4e�hm�x[K��UU)k�tu��v�#�����.��IByy_~�p��u����%�������ڛ\p72����+�{>\�^�|���۽(��no�T�y8}ң���TK˚��:^��DȟD�<Jm���M�%�M��wl�p���?}�"��P�����򾜧��7x~߇x� J��
5��\��P�ApLl���f�Q�1�T�S�+px[��U��Ey���aV�Jq��nm��7{3�D2gNU�;�&_g�Q��~��y `p        h!q�z^U~��������0f����&��$�ܛ��O����Kag�	�k�2Ǎ��(��=��V�;��`��Q�y��~aѽ���\-�jG�Z��æs|PT�js��Y]�|.n�6�����ˇ��ԩ廋{[p|ˌa#������j�6�2g�������! 0�E&m~�!Ֆ��5���+�4����|�퍸.6����T��:�2;Sh>�M}_����#����t�EF�WU{��kƎR��
 �A�        �	�-ZР�mX��-�+<�=��������*g�v��=%�Rސ��J��=���B�⯛d�e׫p�w��}��s>��֠p�7�:�7s(��E
�y�?����tn��mx -c���s?���[�l���;�;G�A���N�&pޜJV-o�3c8�~{l3ݫK�5�Sy����|��-0�����T�y_�]ن��ڙ��Ĥf=��.-�����`���~��VST����@;ޛm�+��c���j�=��pV3u��|��?���ߝ�֢|�fUlݢ��i�zܚ�b��c��kV�x�_���j�˕���lc��9�<��f�<7De�v����w;�Kh>���7�y�ҭ8�^�&w�G~-�<��9�m����t��1�M�?��4  B�        �1L��Y�)���{zu���2J]���ÏTmE���z��F�,�o�s��ն�&���7[����Z�ͪ��l�c��p��=��bN<E�eeV�ͬ��PkP��O���CJww�����������o}�i+8��?[����w�Ҩ�dB�N!��P�}�~s��L|����A:o0]�M�r닓��o٤�O�A��CA��rL3Yh�75��Y��[!Д!#��/�W��w��B�U�~������E5�%�gr���X�5g���ߠ�O<��v��r̪�Zw�ͪ).j��Mg���[�n�[�1�V�rý���e~�Y��P�7�~�۝V'��3�su��2�U���S�QᏋժ��Z���/)�}�f9����a�m�xn3�ƌ�.w��ZI�2+C=��\k6��p�9s�:�m�uNsZ{�u��Ş�W5E�x�+$�f๯3�	2����篽m����E}�uod�3�Mn����ԫF�Zi���
�kW[�Ur>���, @Cp        ~e���h�%��*�Pec�T�kVi٥m����}�K�V�!*wd5x�[�~D�^~Naɩ*۴�
�7%hZ5r�x���mpgq_����@D��
l�ƫǪؚnuym�{l ����C���V(�����A
�|.����APÄ�]r��&���ɇ����:�y��
j��7&xm����h��>s5�[�[7�:���^�9�7�YIc�	��\jJJ��ɗ,�FK�����&h�M�s{��5��(fB�f�]pt���䵥OzLY���K]u�ǅ�~Zs�k2W��VԨ.*ܵ*J+e&��|�IjspW�$���j<c�L�1��a�?̏9w��|S���s�����׹�:�LJ1 mz�~��6˱�D��TC'g����Ϸ�G����G2�}Y�u����U�h�d�5cGY��e>Cf���]�  ���;        �+ſ.��j�@��0�[����P�&8�E�-P�;����D�Ąxj�p���|n~��L��e?˗�sNS��Mȸ��ƻ3�5o�{2�ǒ�Vȧ��5��0a��t���}��b<{�9_�Qd~|HS��4��8F�3�������&�_E�6y��T �[p                �w                �+p                �w                �+p                �w                �+p                �w                �+p                �w                �+p                �w                �+p                �w                �+p                �w                �+p                �w                �+p                �w                �+p                �w                �+p                �w                �+p ����u��(      _YY$        �x� -��毭               �                 W �                p�                 W �                p�                 W �                p�                 W �                p�                 W �                p�                 W �                p��H?#��K�8    IEND�B`�PK
     �k�[�+�sz;  z;  /   images/8883793e-4c9f-4ae6-b420-3a6e91b2597d.png�PNG

   IHDR   d   d   p�T   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  ;IDATx��}�dU����z�B��=��ff��a� E��~���bXu]W�[]W�.:,b �H�!ϐ����=�=�su����ι�UuU�V�ou�Ztͭ���{���p�S^i���6���-��d~���q����n�%�c)E�Q��m2i�΅��Xi2S,��'m��.�FQ���-���Tm�����b0s�;B�~����e�>'Ax���;hW��������߾Om�P�-����sC�z�C�"�"�ZȐ4]PR
��m����5�������(|��D�>u�
e�ڶi2O]�m��$��0���9@m�������+��XҰд�OP�1,�|��� ��r�:�P�����:駙9E�)�3��5Pn�H��~{����mַ_��|���O[�)�٩����~qme����
`q���eIm�ō��!-o��/@Zє��7�dڶ}�|���m�
��-��!��he��x��u��6�o��~������_�$�.Z|��/LW����yf�!������o���h}/�|s�o5$��`qQ�)^�Z�,�̲��n�V4��8Ǧ=�`���e��J4#f4���`ZNѵ�iM4�h�Ry@��Y��3XL��Ч-F�����k6���,��LW���a:U��!�����
�<�.�0�x��N詔<�Q.�f�dw@���H�t5�C?z�v�f�ॕ�g(x����sYRa��]�^��Π�)�Ѡ�fF�Y�o0��C0��+p!�h�Iv;�H�8]���՗
 ڟ��h�4#��H���A<v����A2ɫe�{��caV(�(�Qiy����X����3�W3��@X��?�EI4c��j!]�"�� ,d}�D׮[涯�xSԥ
�3�2�b.CZrbe,�2i#;}Ƞ6�d5k��x�X�F�`��h�o\i:㼹�o�K/<��4�Mc6�*�Y1�g�b�)�L��E��>y�يܺ�652�=/�P�mWHa���H� M��Z
3�3B�����h'K*Mk1\��cC(?z of���.j�X�d�X/�Y�Ҽ���n��iE���1kD�͊��u'�_Q���n8��c�n0e��ym�à]2��ߊ�T�u��=��,�~O;�;=�K�n�"V�G�VB�zR��GV��D�q�[�Y��[.-n���Y� M���1�%B��Y�R3���������Ĳ&X)��X�X)\N���8��������{~���*��X��4#��j藃B�dY֓�P�6�t�H�����f�̥��>�Į�M<�U?!���|�}˜϶ؙ��<�����6��p҂���nz(CT��>���]���߲����[�D�چD".�a�.�߇v3"�8!iU��[ݼ��4j�9����#�x귏����c�觕o,}~�1��WRʂ܈�4�m���$/Ȑ1�6�������ӏ?��J1ޱ��,�u"1":���L��qO�Ik�Ѯ�!:�PuY1��+#1T66b� �x��)�E�z��P���ebJ�p!�BMQY5�=�@_��y����s1��҃ŭ��՚-�]��}��`�Lc�4�E1�8�hV҇6{F�+aAMezN��J�Lo�$�]]���u%P3,�)�c�D&����&�������D��ٝV�J���54���[`�B��2f�V;m-k5�uz0�?.�d��8M3ᯮ��ӅvR��OΨ�l^����C�3���'�(�Hf��,�o�&�^�n�^y�;_�n5m��F<���*�d�[�8��z`��J�`_��D��;��!��VRן,s���@g��p8PQQ!��O��eg�����)Y(��;��o�.X����ΚfX��0x	����k]#�k!;w#�3�:넥PK�C�`���:�E���=S\\�?���H*�Z���Ls�K&��H�h%h]ؾ�!<���(00�L*-�|1q50	}�82� ���X�N����o~�
�;C��W��";f�A�Ě�O���P�a�>2u�R*QP�c+t{0��|r(�F����f�ʈ�g6�^3܇�ۿV[�\d)n���e������Շ�o�C~4�r��U$���i�%I�T���좉�!��:aŮ#�#��Q�%e�����E���}Q�����<�h����4GؿEE"qv�ˎ3��B �%s�%�/- �3s��lᕖ`+�f=+��i�\f����P�I�ξ6}��-v~:����-�CH�&�|���{&Q�b%�z{�EgY�:����:������m�ɫ:��x�x�w�'���]�ǡ�*�t|�܍k�����F�UR`��K<��[0����o��zW�>QgGR�����'ahC�=�ъZ����Qd"���z��ƞy	�?7	�Q2��C&6������ߠ��sz�p����.���HX�2q~>����Iv�2ы�Ƣ/�'��g��iH�;}U�V�
��t�H��)�����0r3C�0������$��̶<p)�m�o�9hi�HN0>{Y�����E��CB�i|��jH6R}'�����4A�kj�*L���V^)�(��a���O��@�k٢�$��5@'"9������D°R{=Grt �8�d��Zh�{��TYEmbЏ����*�4�3�K�ӥzV�Ok_h�� �B�A�C�n��g�gƆ�coB��Y�����j�7�L�����	�W�L�c�]O���m�.[����u��P򳏣���a)��؝�G���!����|U�y��ct��H�1$b���gP���g2��?���J�$������-����v���'�p=���^��@/��%p�{���;܏�+އT�a��䋯��Ӆ���,�u�QMe]���G����:
^�!=Ǡ���#���,�C�����X�H�UP�e�p����lM`5w�.\.�f
7N:;(�*e�I��I#�JqzR�}�t��S��B�ij�V�DM�O�����]�@�O�~S�Q�-�
_K�*�O��Y/�Eu�?�pԏ�6�c1�%��t�sa<�l)�bvH�woC�?��.+��4�.�i�ҎE�J�5��@Z���"�=��Ϡ�̷kl4�IHU.���v��t�LP^�R� �i�T����5H�hB�:!���	!XH�����-��ό�BO&��0��#6��C���T����a�R����Ӣ��	Ȓ�>Mb��!{�P��nc�)�,>3$2��i�fxኘ�0(Ғ:Ns;q��C!��yU���S�c�7����k"@3 ��4�ii3S�y�Nz�J�X��e	v�"`�;���:�B��
A0-A��;��7"��FJ��H�B%]1y�� ��Ĩ(\OO�c�G���DL��J�[�x&�M0I�F�X�'��oC���n�`�D��L���H��hZ��	�}$@D�т�1��y����|4J$#~��I%��f�"ZS��� >�>��UM����f����v�_Nm��5<��`�D�'�UX���H��~*�#�l��*����C�o<uJ!fRC��0�K�����Y���ob�F����cV��?�=�x��&��e�~��%=
3#��U^�:���ue�8�)"��9�"��b\�~9��������i����7�?D�_nw��M�L/��M��s���s��9;d�P�=�O8V-2Z�du/FN ��_/�ȱ!�0՞v��}���%Bm��ϬϨ�0�zF�N��GF7��r�i[8](�X��uE�������$�����O~�n9c7]������Ӷ#��au�浈%�L�o�Z�E�$&�7�N�Y][��HN[��� 95�W_��	��c,>�N��w�����n�yYhln�燈����k���Mm��a�/&�Y�q=�B�lFt��z�G���0�g��9�^���f��� �iaC����!۬8���9h��=p8��$@�
��h��K������o����VU��uo�R��[i)DШ��d"���
�k4{�f����@����Ց4	�z��ڲ�O�'�E@����MŨM�\�v���k�ꢬ��xt0���T�(!�p�ظ}��CH�;�g�����,����K���Yh���!�ӱ��t� �L"M%�CX�*o>�?��C�y�dt6�����ק����g����eE�>-���/������x�p$f�8����ԑ� ���Ț�!�+��	��ʜv�=Dv����N�|�KA���7�B�1)�ljNQ}�=��;d�!�H���3��=���@s$�K�feD�f�C$FL/ll��;����V�<��7#�XN2�˕v2jB�˝�@�����D��k:��߷dt=Nl�p��\�5&�tQ%{|S��3C�sP� Ms�Éd<1�������d,mY��7�wS�_�wi�w�4��~�~0������Oi�Y4L���%�00HD�&R�F;�s�"����*��;�}���e����v���'F����f�&�_}��}�:�Ēp��������n�IcwN���:�r2����l=��X�픭��２�����׊>؅�������쇢1d����1r�LzA#���(�"�P�u�[�!,���сa������rܰe�	?��r�B;�Ey��a9�t�cU�;ػހ�؎��!A#�$��meY��s�5@����2$�	bH�]2�t�1c����\=�	v�����;��=32$�}n��a��ײ��}q�"��8��
�{��@������1V��@�4'8Dk���o���",;��-ȹz�����:�A~��ާ龳�!|����v�a�/ːI٭�myF�$��bV����b��w����A1CF3Sǿ����
s�'��?%|O�Oe*?v��fq��e3����-4���F{���>���^�f�_�������2�nN&S��=��b�,1�E�����F�B��b��n�Ӥ/��a���r�v�z&^Vp2\�2�'Ơ%�0Ek���ԊL$�����Y��U�����@g�^���#�u��{��뀕���2�#ƭ,J�}Ub�����R�B�׳�a��HRȯ��"���J���$�����
C_�sti��2-9$�)��UX��k��D��vH�D�}��C�"r
e�\���F�H�����.F���_q5��
��m@��qq��K�@���&�x2g��E��h�_��I�\04W)�Vݢ��(�{(�� �~qY��y�~�5(�{ 0=��`��P���pd4��ë��ِrb�x�LJ��W�vHn��gZ���Đ�e5,En��ȁ��\�$¿���h�I�7�#nm?�e�����]t����!�~z?�'3��hVL��(+�'�'�![&�Q�����PgL�f��~��AKP�@.f�Ёي6[��\�~Y��� ��K��ٞ"�'q�z����Bv:Qt�F���?���W��l%2�\3�r*��������)l�횋��&
�b�|6��٢������I�e2��8�W�2)5�XA.dk�������0���,>�\�[�b�W�@:�l�Ӫ�8�!C�.��]P|%P#!�D0�³(�~�����
{0�QKƌQҴI_�@xYhN4�0��� �(%�BɆ�z��"Y��j\ͫ���#��+p4��:�t��u#?���V��?�A��v��(m���b���#(��5��p��'VW��?$¶��8����Dp��g!�櫰U׊	ȓ�VY%Dw��A�ܙ0� ����m�VQE�"7��ar��L�@WS�@FB�Zb$$Y�s��1A�Ǎ�l�8w޿�E37N�1	 �z�D���C��XfxXYXD�XQ��fأ��Ӌ������G&M���`	b�ٽ��	�[��i'��:Խ�dB�GM��ޤ6g	z�{�i��썶��iO�<t@(��Ѐ�<�N#������V�
���;���$���[X:�z�ɈP��(�w͜La1�Ngo#�#@���pVz�a�Y��ٵ���2�cN�هk7��F��wb����U����H��B+�1�� �1%�oG���D�o�V��.�/��s�a�0_�
�e���3�Z����d��ayE3"yi�y�V��AݎǬn4�^��[����E�"�cq?~/��2:;;c�_V���w�Ia��~<m��Q|݇�#�X>�vZ��|�k_�/cC��=�1�G�B7�T,��A��r(ⓗ�gl�ǯ�n�:&,Di#��L�W�G�n���?�{�)���"Z �a�i��amA����Ah4I���'�4��p䅃�R�(�P,L�J�*�|�g�A<V�̄��-�i),�憢-`e��f������^�+.�^"\6��g������><�������L�1�q��V=����i��W�{��N�����&Y]L���$2v��D�B����C��'�Z�] ��
;Rezv�W��-H?|nR��6!nu�%{�T8��=�뗠{Z!�H@=F��ƿ��+�<�V5��	�3*I�S<�[u��ۧ݊+;����DҒ�2�� �ǘ�@~G1�~��P�?���9Kt8S1�w���x�[��~��⋌|�drF[�ۍ�r����b�)fw	�X�f�Kb,��C���aܶE��c/l�r��c>�b����!��C�¦�{�|��HZ�yb��V��p�57N#}L+��9,��}R'��>$��ܷ�����k�M������ʍh��M��'0�ė���-���3O}�8�u�pa8�"1�����%m�`.�p=3���'oڄ"~�9h�h�ӆ�n���>M�L�q�	����$��_R!]��5lw([�>4��<#'�K���6v�JvY�hʆ��
��꩘^6��>J����U��'�)�$%Oޓ"�y�Wx`�bC�V��eZ9�2��-�W^u��\�(Y@��сM��b�E��х�9�f��!M�C����ڇ����a�V�qZ���c�A8�[HIy��@�	B�_�S^J�,C3K�Y�E+��bS eǓm/f�*$�����6��d;_l�r] y!��?!�0����g�M��9�4pk;w ��DG�+~���tE#}�o��+j��	�� �(p�%^C�=.�Sߘ<�@�Y7Ŕߡh�W�ؐ���%
B_��͹�"[�Ղ��}E4�{C|���p�Q�dВ1X\ޜ��=�(j�:�&�XYY)`��~���	/��"�2CfIr���`E� ���F��w���;9����p(�7P7N��,%���ɺ��pVT�}�K-�U�\�>��Ŝ���0;6	�{��%dx}��_b�m/�ɑc�����,8�>I�e���R#1����*w�\(++CMu�	j��̙���ƻW�p�d�$�h�����'�R(�x�ڍ� a�A�rF����ņ���`�ß�{��<�JL�~�= _x"0�
N"�ԣ�#_DQ8���/��D�\9�+#!�]�E�2��.��d���
��p8��H���c�/ Or�I[,EQ���x�C�#�#�%��=�Xk��bt�0c������5t�n�v䈱`��K0U��g&̸'��tc�3��D��|����(��:Ay$�e��хzlJ+�EO���a�H�����pCQ,S[60�i@D�0Y�G��!f��8󯺺5U����#����h����Ç�q��֬�v1��*2��xb���21&���o3�~�, ���֞��}�8�2+�زb/J<L�4<<Hv��N��*n�?X��"�,p��!UUU���LQ$=I�B]�BkɴL�k�	��-R'(��D"�λ�����+�PRչ���l�%.�,���B3���hoG�"C�|[+�o-��V�sX���&e0���{:�%��԰̜?3z�V�ɑQ\�e+"�Q2��ˮ�h_m�ˠ0[U#G��{��̲"]ŵ��7^Ƿ�������[��pS�EL���FaUk�1����ۈ��|I@� [�Ծ��ń�M���[n)@YYg�0������,1��Ċ�8ғC`��۲
�S����E:�B�Dn'��GM3�FY4.�ˍ�d���Uը��Ĭ8���	�&�U���f��b�J7?���d�󷏡`7\֮]+c�I����}xf�s(&��,�l��l�㍞�4�5��e���@g�S"��}Y�#X��0���(��*����`���;	�T��d.I��4��@� ��P��]������8����F�57>�������>E�8�����Lx���!�Z�
M�a=�H�����µRc�#u�PS4�Uh�i-z������/��T���F��~�`��b�ϋ4d`` c��|�=Z׬1|\s0�Y�q�Dx�wX-� A���7�N�I���	T�!�h&O�m��+�*��[s)uj;��Иe�p�Y%%�������8�����~�H@�0S��q>��=�^{F��`k��\B bU�z�n����@U]����
l�Q�����"�W*.���D�*u����&h��D�z���3W��4F:�	x�⢘|ԟe�n����*�X%iى�{�xz8G�*HӺ��j�n���2�/L�"�Yb���8�&�M/̈��^�S�I[�I���ҁ�"SXI��e�S3F:�}�#���	|M9M�O{��]��4S�؞K�еե��|~���9��4�	�zpa�	����:��'�Q�NzM���l������.f�[IR�$�.�����!�zc^��Z�
Ȭ��ŃH��%f�[Ҁ6��Z"^��Ļ�}�S�np�EƲL7��PL6�H&�Ԝn�̭��s��%9����"�W"�����>�n�B�m�&l�&��<Y%�c��/��ƅ$}�<76���ǡ�3��7�� �Ua�I�����~�N6��[�R��a�<�^	��):�O��}8j+B�KAM���(F�:�*m9^�n'n�����p�ھ����Ӄ&E���2�W#zp�'���ߋ��h��ۍ`�	|��# ?��ag�x��Fr'!\'G�n>�p�x��L�-
��FFFP�~-���j�oWz!�IhW0~��aTUV���6��MU��?���M�Aó����7X�В��t�3���>�I��`�-��a��j���c�h.;����a�:Y��e�Wxx?�������=d�0�a8���|�)A�އ{t'A͙��YtG��Q�i"
;;N��|@A�P&��:E�IG�<St�2��|4>��b:A�k@(�0��DC��**��r/!}�z��ć�,Q����O�O���&K}�=��1?�)��p�s������y�#�8A+㹗;e�w;Ĕ���G04�4 Y͹]�*xq��Z��>.ғ\�Z=|P�K�rx9��l�_ºj%��<���ݹ�!|E�D���"��Jp�����&{g��{��9��� w[{��}��dk:�O�'��
�A���A�P19�uB��đ+pP��JJJP[[+���ȉ�jG�E6�<��|���R���&�1*�d����OJ�.H�z�
]$�͟��̨&��!�:Ja8hL~�����;}�L~?�L��3�!��8qa�'w�Y6��#�����_Ax�F��4�������L4�e�턪&V��k��N����Alڸ�_v�ܱ�>�(���66`���@��.�9b�X}%�^?��W�QRQm�(
�$<�.!㩟�ub�h*���j�e���+���#�����\e�����E"�|�>LsJ�M�c/��.,��`I���C�xP�_�au"�X<dHB3�Kl#�"�;���՝��34�Pz9M�Ёɭ�D��Kn�-[�o����.l�$�b����[�ك�^Z���G��P�����=�z��`��M��T�JZ����N$o5:6�[O���}b_���+Ѵ��h�x�U�2����=e;��,�d�`Ög���[C��~�$I݆h �FZ�	}3y�\YfH�~��L��$N�<�#�w=�����Σ����w�p�͂<�椩�oooǦ�N��%�}��b�5]�ޯ�iSv�p=�ů�g�^{�G��}�qU�r,�4�e�d6C��T��6�uB������'D���&�E6���14�M�P�#�1��*���g����fiqĐ�-�səL�����	#���iF�S6�['tF2�p9{���c�Qݼr�V���C���x&����g�_��ݮ���\�"T3��=b�o�8˫q4���چP,�DA�a�l4�W+	\alR��#d9��������:>t@���"�Y٧zc7���jY���Qw�����8����w
Ĕ�;Q���Rz�%����V��N�(Ny��{�J�uv��!v�gl�"�w2��+?���"�/kF�nZF��>�Bg��\�ؽ�m'��ϻ�x�`�F����� j�����
�9=ة{jjs��J7-�GFe@1^8A-i�1x_��&�1-��3�5�l=KlSQL>�4<��F�����M$F,(jY�T_����G2)n�8�H��@O���#�ۀ�@|g���+ϋ�
����!nK�Y&E޸|�����>�gt����Ҟ�獻�%��J��)���g���:Z��Hϓ�i#��X��o�.i�Wu<��,������蓄�톯_2��L���[$sv�M:jz*0�\�;׵""�<>��\,E�[o�,� C=��C����aD��`�!��@"��BǏ�H�y"P7���u?�G��pM ��S�˼�e���Fq�v.Ab�cɮ.���n#��!+���6\�!�^���$&�T1ƤQ�;t�C��=C4=��+���QxRQaq�R�s���=�:'iZ���[�l�d섽�A������u(�����dMK��J2�q�1b^�9����Ȟ�#�W����Қ�:q�
�q��%��O$MM�ά��i���x� ���	z�]n��WP�U���v$����b��P �w���%w<�˗§�IZ(�+T.ݶ��v}��O��b��^MR"J�]�+क�	؊��4{ݰON�E2:v�؎�&��(�B�f�N�׹�T�[OB���H���-kB�d��\�lTo1ĥ��2MԨ��1�Mے͓���0c�o~9p� .��,�P�n$��;O822��=>�.���J�:W�3!r`/�$�#���ZS�T$*�a:[�����!��4�Oı1��/�U�\���~��.x��Ι����v�vثV������?*�Qݼ =|5�����q�kP^���ŞF5F�՗s�#���{ϫ�QG��b�J�J��-^�3���J������*D{���E��R\����)	fV<����N������b�����"$߽[����w�}~�[σ�3���?������>�?R҄�n����)���	f����[�
S,���'1�%��r��r��mr�K<��r�6�S�y���c� 4;$�8X�<��� 0&i���?Ɨ��c��|���ouu��F�ܫp��X�Q���h"�,��+���z߻Cl�)�~´J�6��!!N����9
�(Ь����8c����/�燂�V��Õ��V�E�
����bqó�\A\�j���&�����w�,2��kk���l����ϣ%�%`�d��0�����!>�����y��D'�����w���s��>���p:��M����[��Zojj��3�YGɱ�����[k)�+�ov����Q>6������4����غ��<��X���-JHS'�H����Ŝ5<uޡ.�ϲ`�D;���`ǵ�@��Ni������POn�c~"C�H�ߣ-�{xX�>��?���ċ�}%#����
��8V�g�Y��8�ÿƱ�n|���ओNY�<Ax�d0�ǟ~/��Cv�W�ܣ͒�Ęs��/}5�ӳ;�����5��[��}��nNv��F'o��ྀ̽s�y���H�Q�;=����[}����H)(���o5�!��J��H�1�ɨ�Bh���0"�Bm_%��co�����W�2
�3�g����뱬��'wubt2A"vj�q���"S�"�p������GCC�4�]�������H�h�T%��&5Ǵ�[�DL�N�\V��V��kO�ˌC�/��T��N�J.��.��|1���nCI篰�p�8�)CW���KkE�n!���`�-��Ѩ084�~���wC�"]B�L���g�j��z�2�#�ܗ)ű�w@"�u*�0���7� ����2�f��ĔS��X�j� ��{L��s-湓�D4��]9�jxz�{F0H�т$=��컛&�
p{��Đ�׈�-�rbf�<x�o�ג�'S�֪
�%xxx�ؕ~୅�>H@`�.>���"�S���Hv���a��˅b�/3؉u��u�p�}⁹�����ԥ��V��Hb�}�rk������$#AB���1O5�����n!)Kbq��xN^�Yc0_�����Z*�X���l�t��!��.���^ ����rb�˛��ݐV4s���,^���&^��o=.H�{HR�y�Z��� ���9�u�J7�у��Z�hʐ��م�"ZeV���4�d`n�Ԍ5��3b�F��S��S�� ��E*?G���P������˦��=4�Q�ԧ�:D�w������01/.[�=0:�	������II�e����i!>�ה���5��$�1E3�2��դ�V\',vf}=��+�C]���!5��!J��o����^%^��o�.|}7�)%�'�@�h:�}�=��P�~9;��_A��ԋ[x�X"�X�J�����I!9����O[����@H��,����Ѹ�L$11a����,����pd҄G��IBN���"@F*G�,�XWg�{(,��܌6�y�t���Z-	�$�+��_�u]����Q��J�af�n�b�rb����Kj���̯�f��9V�"� ����@?�À֚��Nf$�)��03Z�u���{8���&ie�=D��_��H�S��Ey�6fF���A��/6�#qw�/g������z���p�l�ĺ�:���rPkYC�@asÝ�Ƥd�hξ`�7CK���O����<j�A2��Vd72�x�&o���k˪�%h�U�S���4.�[`#��&�z��T���*¦�H�z��[@c�j<.�pXr�}�b,	��������mB)zV��.�D��{Ǆ(.�C%=8��Wn9y-�����`Z�����eZ���gosh��R�MZ��!ۀ7�Z��;�$⪞J䗳kO�f����]QPJ��C𰴴T���WI��'�$���Cq+�	11øp�>��9�<���J�-ƓP]�VA�ׂ��W�U�}N�Q'�l�h�NXeS.��"��yC�@Y�?ہq\��f?�z������ET1�.o;k1Ђ�>CY5Ը�W�;V�-�O�<F�W�31�ҿh�2����}�����w��V��Ob��^�$��I7�����Dk��ܲn��د�DVn��n���K8W�&���w�Wހ�<⽯55�Ѽn\�R�߭��O+���B(k��k���r�D�-����)B5Y���G�[i���z�O߄3�p1ڡ����E�YMm%�VTQ8b����X�B*�� ;����I����,�Be^�'z�i����l����al�#��<�.흃�b����q����
�r(�t2t�3���Ca%[G�ض}ݍ��
.!yG�u=#�]����~X)��l��.o�U׊�B�3��S�.e�H�Npr��A��$�O�/Oo�K���P���	G���=�����xd2��[��U)A����C�2��e\���À3������$z��X�:q��d�P^b��t� ��G�f���V"�d��#�ә�+ԔP�)o����K���7�k�"�A��~�zACS���$ho�3�q���.~��KjX~/M��km�E�pޣwuؤ��c�W�V\0u��� ��IؿV>��V��SCp�+��2ـ�᰺G���BmGt�V���ŧ�,��&nk/rQۍh?8�J��S8�����ʋ�9m�� ���D�~"�l��E�E,�~R�c�e�H�ץ�Շ,�ʺ<4B�.#��M��&ɻI�3����Z���v�b�b�c$	4e�eR���5��}�m���~6Ĕ���^�i_���O��Ж��fb�&7y����c�g��$z�Ľ�ޏz��`����#�ȐcCLl�5N���ࣻ����bbV1��Lz��ڲ@R��3�1s[��m9�C�k+e?Sǜۈp�OL"�A"vS��2u�ܘ�D:� ���|.$��䤱?�&�B�L��mMNX/6��2F��ߊ����@5ι/���Ǡ�qz�S`9S�C D;FS���z��&fӜi?��|�-��?�
��m.BUg�h��AB�˃=�q�]x�tG��T�����q�\�I���e��c�i�xz�lgP��|���ݫ������� ��D��s�F��>z�7��Czl����`�&N8�','g�6�"�2��wb��;�hX.z��2V�|H��������>�H�A�h��]$����cF!CL�0��G��,Ѝ��^`�Wel�w?�'N�	[f�s�0C�$�rK�� D@�|Z�i7�9��8�ϫH)�%��a����A"f���B�4r��"��Ldm�=��OT�zf�qĬ,c���}�"�ħ��~3�x�
A�,����Z�U9���.��b?��SH�E<�h���"\��8�%���.�i$#p�*�"��
�E�!�sz�ԣ��	�=���d1QO�W��#�uςl�S�=��Y<�.D2���ȰnO{a�t͖���o�-\b�    IEND�B`�PK
     �k�[t���?  �?  /   images/e2e2c934-b375-45fc-834c-534243cbf361.png�PNG

   IHDR  L  	   A_*   	pHYs  \F  \F�CA  ?5IDATx���y������ϯ�i��qa�x�DI<��D��x<j�5�`��db&;;�&3�f�8��a�hČ��Q'8:*���!�A����~[U��B74PU���������#������6    �ݼ�曓�,�'���<�4dȐ�`+&    ��K�v��`+	&     @�      y�	     �<�     H�`     $O0     �'�      �L     ��	&     @�      y�	     �<�     H�`     $O0     �'�      �L     ��	&     @�      y�	     �<�     H�`     $O0     �'�      �L     ��	&     @�      y�	     �<�     H�`     $O0     �'�      �L     ��	&     @�      y�	     �<�     H�`     $O0     �'�      �L     ��	&     @�      y�	     �<�     H�`     $O0     �'�      �L     ��	&     @�      y�	     �<�     H�`     $O0     �'�      �L     ��	&     @�      y�	     �<�     H�`     $O0     �'�      �L     ��	&     @�      y�	     �<�     H�`     $O0     �'�      �L     ��	&     @�      y�	     �<�     H�`     $O0     �'�      �L     ��	&     @�      y�	     �<�     H�`     $O0     �'�      �L     ��	&     @�      y�	     �<�     H�`     $O0     �'�      �L     ��	&     @�      y�	     �<�     H�`     $O0     �'�      �L     ��	&     @�      y�	     �<�     H�`     $O0     �'�      �L     ��	&     @�      y�	     �<�     H�`     $O0     �'�      �L     ��	&     @�      y�	     �<�     H�`     $O0     �'�      �L     ��	&     @�      y�	     �<�     H�`     $O0     �'�      �L     ��	&     @�      y�	     �<�     H�`     $O0     �'�      �L     ��	&     @�      y�	     �<�     H�`�Y?��^Ql<��vd��Y{F����w��/ʳ��E�|V,>��&��;k     �����wD��w�b��E���?���������ҏK?�
_˛{-�5������u�o     PӒ&s&~wX1o�~���J��l��~����;�<�k�;,����s:     �II���=���E�,��J>��l��/ߛ3O�y�ߜ������      jNr�d���}��?d��k�,bT4fOϙ���{��?f     PS�
&3���y^���KpuN�o1�ƿ��1��_�     �f$Lf��7�<�5��K��H��>1�8�x{�     @�H"�L�xeS䅻��������s��g^Zz{C @ɧ�AQ��������TvX,   �:�D0�=��E��>/��;o������\ T����-��'Q��~�X�O���1=    �P���w\٫�;�C���б�һ� ؉�i1 ��c��!�4P��~��t|1`��ߐhl<6  ���5�[��+�������r������l�KK���IGs�3
���������>��_^ ��/���Ē6��MS��g?	 �:�o�u�std�����ڏ�~�lwuL���U������� ;X�|�b<Q��G�g�X\:�g    ԩ�&�ĉ��v���Ǉ`��?�F^�%{m�����.�^��p��   ��������}
�跳>?˳� �@�����X2d�'E[��}"V    P����رo^^�k'ɣ��A�Nȧ�AQ�� �c����gg�cm    ���&y�V�y�$�,�i�[ HK�||,��e ��&.�$V��ã=    ؤ�&Y�3ߩ� � �����1���KG�M\�->_β(    ���IG�Ya'.� �[�B��<*�m���[���U�   `��:� @=�_��#��Jo7�ј��e��7   �NL ���Gk�qo�m�M\�~vx|+    �4� jL�B�y���������a��    �K �!��qA��O�����?Y\�?    �L0��?_�<�!�(|�B%�\�7    [E0���tv�"e�e����K��D��7[z��7�E1�d���  �v$� P����Ȳ�"e}�߱��l�s�=`��#�ֵu됍��Q(   v$� ���^�߾�F��9x��ح_�   �I0ل�=���!�G�]v�b{[�-����+�     P��i���>=z��������b�+���3�     P_�we��G�<'z�6h������"/vĲ7^     �~&��u��>4��_��~*V����X�"     �� ���e�!��/k��=0��x.     �� ���*�wVS�-�D     j�`R���٥�M]�     �n�	     �<�     H�`     $O0     �'�      �L6����-��|SSS���/     ��#�lB9�l�X,     P�      y�	     �<�     H�`     $O0�@�P��}�n�|�x�g�755= �X��]    ��&Ȳ,�������c��ˈ HDG�ϯ    �#�     H�`     $O0     �'�      �L��b��/v�~     ��	&%kWE^숬�Щ��W/     �~&ey�ߞ�{�۩�Wϛ     @�L޵�7�̓��Ȳ��׶x^��73     ��!��k��?�;/?�9�C��X�"�?�@eF
     P?��Y:cj�[�8��Sѣe��!�c�~�^z�M     ��"�l`�[��M}Dc�~�w����ߎb��.��Q�[[['v�w�����.     �{�e09��S�,���7u��g��V�ѶtA��F�,�Ύn���     @���`r��g7�^���Y�}=��J���Q     �-��`���z��5k��eٞ     �E5LZ[[��^�Ȳ�      �J5LZ[[�eY�O���     `�d0imm�j����B      l��&�ƍ�v��o     ���T0immb	     ��j&��7nt��7     @7��`2nܸ?��|B�e]ڳ$�c�*��/      tJM��[�,ۣ��]�;���|     �s�>��;�����[���m�3-�ɟ     tN���P(\����tu�yY���P�|     ��Uu0;vlyfɟl����+�bP���f�_     @���`R(.��1^}s�N	&�-����      �_��1c�����m]Nk�̷㸃����r�Z�<�Y�6     ��W��������Ka[Ǚ�tu��֒8h�n�#=>��      jC����k��~57أ_
;f�Iy�r�     jCU�Q�F���1�5ޛ�WƓ���<$��uŘ����&     @m��`��ܼO�Ow����sc���ư-�=���*ˀ     ��*�ICC���=fG1����o�ғ�A}�c{x����̜     @m��`R2x{�r��_���u��>�o��[,�,��j�w     �E�L�ۺY�hr���3>�w|r�A�e۶��5�⟞����4     ��T���[�/�PyFȿ<7;^�ݢ8���c��ty���b��o�#/��a     ��U��$��i�4s���~�˕幎�w`����^=6�̼��*���ߘKV�     ��Ue0��f�[Z9
YC���=���~}zF�r<�#V�]����/ZKV�     P_��)�y%��      �	     �<�     H�`     $O0     �'�      �L     ��	&     @�      y�	     �<�     H�`     $O0     �'�      �L     ��	&     @�      y�	     �<�     H�`     $O0     �'�@�1cF��G?�ٳgGGG���m��b�رq�)��.��     �L��-X� Ə˖-��3o��fL�>=~���	'�g�qFz�    �*�j��O?ݥX�~k׮��~�r���q��Wf��g�     �D0�����-�̙3�2�䦛n�Q�FU��G�B!     �`5�S��T��~�����[�[�n]<���c���q�i�Ÿq�b���    P��qMMMq������_�%�%�=O�y�Nm��[o��7�\�P��c���:9��c���!     �`u�w��q���w��E��C=<�@��������b1�z�ʱ��Gkkke��=��3     �`	*G�/|����^��N�4iR�Y�f�ϖc˄	*ǁX	'cƌ�^�z    @��R0imm=��2&˲cK��y>��~� jV9z��K.�${���O3f��Գ��R>n���=zt�u�Y1|��     �5[&W^yeaڴig�y~y�eG��Z�� �CKKK�y晕�Y'�'O�U�Vm���˗�}��W9ޛur��'Gsss     Ԃ��SO=��iӦ�Rz{�8�xo�ɟ�ٟţ�>?�p���K�z��Y'��'�tRe��C=4     �ه������y�_�9�d���g����_��I�#�<+V���+W�\?����/�8�9�     �FŐQ�F5���ܖe��]��\q��Y'�?�x%���⋝z�7��M����y|��ߏ�;.     �͆�$kii��X|�^�zEkkk�={v%����?�e˖m��<�+�M    �} ��7�/K/_�-(�������3×544    @5ZLƎ{D��;���͋|0~�����o����
�B�s�9    P�*���+�,�����ށMhoo�)S�T��z��g+�K��C������     ըH~��_}&˲�>s�έ�$)�Q��;�t�ٖ��=zt�u�Y1|��     �f�`���eP���V�MRޠ��瞫l��Y�e�;��q�	'DϞ=    �4�;v����$m֬Y���W��Z�ti��0`@�3&�<��2dH     ԚƆ��1]�/ȁ��r������J(�:uj��}o6I9�|�ӟ�ҟ%    P��<?6�����kq�����ɓcժU]zv�Сq�i�Ÿq���    P����,��],�	&Ĝ9s�X,n�����W��^�z�����~z�1"     �My�w@[�bE\x�1o޼n����&9��c�]v	    �z՘e���6eʔn�%�0r�'V�&9��     ��@�ʳI�8�8�S�w��    ��j�ȑ#cРA[5�d��w����ʲ[���    R%�@�+/�u�wtz�������L�c�=6�1     �oJ�0 ��o     [G0     �'�      �L     ��	&     @�      y�	     �<�     H�`     $O0     �'�      �L     ��	&�-\�0�y�X�x�V=?p��9rd���'     ��`l�����K.��˗o�8C��;�#���     �F06�n��XR��oƝw��^zi     T�ج9s�t�X3g�    �j$� ���y��U,    �	&     @���ƍ�]v�f������_    �Z � ]֣G��u�]7{Oc�?^    ���o4    ��	&     @�      y�	     �<�     H�`     $O0     �'�      �L     ��	&     @�      y�	ԉU�VŒ%Kb�=��,�    ��L��u�]q�7ƺu�b�}��뮻.�     t�`5�׿�u�p���y��Y�fŵ�^7�|s     �9�	Ը�^zi},y��	&t��k׮��ܜ9s�����s,    �Z!�@�kkk���]�˴i�*    @�L     ��	&P㚛��V��w    �"�@�;�â��1��ۣ�s�1    P��qÆ��|�;q����;�ըW�^q�y�Ÿq�    �	&PN:�ʱ|����<�M�>}���!     ��`u���%     �:�     H�`     $O0     �'�      �L     ��	&     @�      y�	     �<�     H�`     $O062��X�hQ�}Ϟ=c�������     �W�	��ڵk�+��������5�\#F�    �z$� ��y�Œ�ķ����4i��&    @]L��^|���V^�k�ܹ1lذ     �7�	�^[[�6]    �U�	     �<�     H�`     $O0     �'�      �L     ��	&     @�      y�	     �<�     H�`     $O0     �'�      �L     ��	&     P�����+ؾ�\0    �jU��#�`{+&      �	     �<�     H�`     $O0�khhئ�     �J0�>|xL�:u�ך��c�С    P�`�/~�`2cƌ��ݻw\y����     �H0��u�]c	1}��X�hQ�\Ϟ=�������    @�L��ѣG�1"     R"�      �L     ��	&     @�      y�	     �<�     H�`     $O0     �'�      �L     ��	&     @��y�ǓO>��̜93֬Yө��o߾��~��ȑ#c�����а~�_����#��+����N���wjܦ���s�=㤓N���??z��     �J0�:���W]uU%ll�r�={v����[o�5����e�]���b���[5f[[[̚5+n���ʸ?��c��    P��7�t�Vǒ͝;7.���ѣG,_��[�,�x��+��n�B�     �F0��p�¸뮻�u��r^�]ҫ�^~��xꩧbԨQ    Pm�qS�N���";��O?-�     UI0�W�a��,����|��/���k��/������k���?���f�1eʔ��ۂ    �	&P���cC�`r�%�ti���;����M^;�s��_�z444tz�9s�lL6�]    ��`T�w�yq��V6}�]w�5.��.�    �Z#� ������C�F�=    ��	&�z奼6T(    ��	&     @�      y�	 Uo���Wf��>�>�ڶ�X���y   v�<L ��mKz�)����b��پ�-֬�{  �'���У���Y� �OG���I�Ʀ����y   v�����<`us�9��Ӿ��j���}��  `�$     �`      �      &�z�{o��n�^�    ��	&�zGydL�<��:�     �w�	�^kkk̝;7��(�1v��8���    ��	&�zY��W��ո��+?
�     H�`lD(    R#�      �L������s��[�l{�G��    T�j�'?��J Y�x��s��zj�l\pA<���f͚�����q�y�    @5L�ƕg���?�c�v�m�p��J@9��sw�׊�Ç�]w��&M������    �j$�@:th\}��Qm��k���    P�      y�	     �<�     H�`     $O0     �'�      �L     ��	&     @�      y�	     �<�     H�`     $O0     �'�      �L     ��	&     @�      y�	     �<�     H�`     ժP�B����v��	     T�����M�;�     H�`     $O0     �'�      �L     ��	&     @�      y�	     �<�     H�`     $O0     �'�      �L     ��	&     @�      y�	     �<�     H�`     $O0     �'�      �L     ��	&     @�      y�	     �<�     H�`     $O0     �'�      �L     ��	&     @��˖-���;�~��8��c���Q/^�<�H���ǉ'��
    �j$�@�[�zu\x�������>�gώ/}�K;�{-Z�(>���Ƃ*?�~��q�wİa�    ��&P�L��>����;.�(
�B�,�/�Œ�+VT���W_     �F0�7���έZ���LW�~�bg�;wn��    T�j\��Q+j�    iL     ��	&     @�      y�	     �<�     H�`     $O0     �'�      �L��eY������3�Z�j�s    P��q}�����'�|2�>����,Y/���F�w�}�     �F�	Ը�~���<����ҥK�s��\���s�}�Y�f�UW]��&���    �	&P�>��QG�>��Η���[��.�(N;��$ּy����o����g��ѱ�����hmm    �j$�@��W��?��&�-�?~\s�5q�]wU����?����l�TB�<�֭����=��hii	    �j$�@8蠃����v\}��zϜ9s���f|���}-?��m��e˖ń	�{�5k�l��}�K_
    �j%�@�8��Sc���q�7nr��{^}�ո�����D%�>�K��r����\9�﷤<�����F�=    �Z	&PG.���1bD\w�u���/o��g�y�����'��Ǐ���o���,��'Vf��7�ߒ���8��+q�W�^    P��3���{�L�2%n�馘9s��[,cҤI��c��g>�8��bȐ!�����C=����.���766Vf��7�8p`     ����ȑ#��c��ɓ'�-��o��և�[ެ�'?�Ie?����/�@���G[[�?�P(�)��R٫d��    P��c�1f̘8�����[o�u��D�<�3fT��ʲ�f��Tb    @-L �e��<��J<)�")�CR^jk[q�q饗�     �L0������=�β^����3�	��.� !���� fť�d-��(-�h圥�ǶDT��Cת�T��9�Ğ��p"��B�.nB�T@��p5W��o߽KN���f������{��;1����<����>���Ї>T�k�ܹ�v��m���������#�    �V �@�����s���:����?���)9ꨣ꟫�    Z�`�c�=��/�s�=7n���뮻b�����K/E___�=:&O�\�d���1eʔ     hE�	�Ǐ��|�#�     G�	     �=�     Ȟ`     dO0     �'�      �L     ��	&     @�      {�	     �=�     Ȟ`     dO0��v�����Q�FE�R	    �V'� �lٲX�pa,^�8{�X�~}�x-���q��������P    ��$�@�-Z�^{m,]�t���j<�������7&M�g�yf�v�i1lذ     h�	d��&ɕW^��w�6}���~����r�Yg�駟.�     -��(�WSJ��Z(��7�<����g�����1w���'�	    ���SJ.��hIEQ�w����w��ܩ�^�r�p    ��ڐ\O�`-�6�ȭ��W_}u<��#�LWWW�|����އ���W��U���7�1�\w�uq�9�Dwww���    h�!��O)@K��Q�p���%˗/�gj�����SN9e�7Dj�M����ƽ�����Y�bE\z��9Nj��9s�p    4�Z0�=�tf M��&ȗ�����;t�ĉ�2lT*�8餓�ˢE�⪫�z���k��K.�����/})�8B�    [{[[ۂj�ڟRj�i�b��g��>��[^[%�3t�q�W_~�����������׆�:��bΜ9��W     U{oo����*�O�)�_�>.�����%���?������~���__~��_���<��������_\�4�vX     4��Z��!�@Ӻ�k��~��{�w=�����P(��	'�P_js���Ƀ>��������.����!�     M=�̟?��������Tjo�\��[=7a�%��v�N%�{�{�S_���ַ���x�裏��V���    �h^?y�g���mJiT Mc�ҥ�z��-�|��q�W��ѣ�{9���o�\~����I6W�K0    �?����?:s��O����4�|�ɭ?���5�lTr볟�l�r�-�r��M��&�    hD��$,X���f͚�R�@S�ɵ5x`�Z4�=�`�f͚     hD������ݽ���o�hJ�rΒ�ho��?/QE     4����?�WgΜ�XJ�;�{ M窫��h�|��     h�otb��?>�S�loo�FJ�_��M��lm�u     ����N�t�M,Wg̘1�J���)�Y�     ��p�7��\�5{��O�[�nZJ�r�Т(&�ۣv��5��     `�P0�h޼y����ז]�����r�_     `lS0��ĉ#���zhժU�aÆ     h�	���s�FWWא=���D,Y�$     ��`     dO0�&W�T���`��p`C9D    ��L�����[�s�=cԨQ1���o���8    Јhr'�pBL�6-n���~ggg\t�E1�>�������>�l}̘1q��    @#L��Ն���׾�/�U�VőG���P[��^{ŏ~�����[�Z��{���7n\     4"�Z@mn�c�=6MWWW|��    �F'�      �L     ��	&     @�      {�	     �=�     Ȟ`     dO0     �'�      �L     ��	&     @�      {�	     �=�     Ȟ`     dO0     �'�      �L     ��	&     @�      {������{��{�1v��lo��j56�Uc�Kk�����g^.��     h����J��=���IcG�����W�?��Z��x�O/     ��2�EQM)��g��>��	1���bܨ����G�}|}y왗�ǋ�Ǌ�     м2���������=����W��gʞ]��ǂ�=�<��z     h>L���˕Je��{��w�ON?�Mv�J%E��o��cG��_?U�     �NC�����v�����5�c��������-���â	     4��&EQ<���9bX{|�}��X��a����G���x      ͣ!���G��ҥK�/7��{��ĸ�4כ���I�Њ⑕/     �2�̙3������r�C;�~O�~�1R��>vJ|e���     M�!��k�N
&3��7�^��G0!�z�      _���������.O)ۑ�L�0:�?*۴C&
&     �$6���'?yn֬Y?+7Oۑ����
���Ǝ��^X     @ck�`RS�T�Q���'����wL     �	4t0�������r����|�n�b���*�'t�_W     ��:��T��RJw�K۶~vϮ�1����-     �����d���̚5�r����Q�;b(��    ��i�`R�aÆ�>�������am�J��C�|     ``�"�,\�pMww��)7�ˈ�~.UR�����     ��4E0��?��===�U��)�a     ��4M0�����yOO���j�{)%�      ;ES����������V���R      ;��IM�M�3f���v}���      �MLjn����Ϟ=��u��}��=/�T	     ��д��f޼y��էzzz�)�����     ���:�l��ۻ�\����sR�Z��r�T��     ��d��������rʄ���٣�w|��?2      �DK��n��g�����u���m�|�}X���h�{վ�����e[����(�6v���Α��3     �-Lv��c9!*����bՒ��+/��*���7\����E���	     �4�������[��s��1qڙ����ņ�V     �:�׌�x�ƒ�R{G�ylO���E�?     �� ��f�w3���G���o{g�~��      Z�`RJ�J��_?|�~�	     ���T6""�_�6|d      �C0�نX�]�     M0     �'�      �L     ��	&     @���T��X�z�����cĈ�:::֗�@&:��    ��`���(b͚5[���l�`2u�ԗ�Շ �}��    v�     Ȟ`     dO0     �'�      �L6�R�O𾹎��      Z�`��J��ƍ      �	     �=�     Ȟ`     dO0     �'����r     ��	&��+���u     ���T���+/��ac����{*     ��!����G��SO}���7��5O�>     ��!�����7FL:(F�3�/*�Xu�Ϣ��      Z�`�QQ�3��1��=����69ݿ~M���X��      Z�`�:��LjQ�ewǈIFǨ�Q��^x:�>�HT�^	     ��&[�꟟��z.  xs�   h	�	  ۭ��-=�   �f'� ��*������_�����L��t������_�{�h����˗   �`@�K�����fAqw,�ߋM�����ѿ��tt�]@(8�#�  � L �����bI���_.��D���o���Ԙ    l� �L��%����q��������k.
    L0�&��և�:�ܜ)Fmv���ܨ��dP#   ��L �I���Œ�Qn�P.]���O�=�^񩔢    �)� �X�w���(��rw�f�ϋ%1��-�]�V��   �7����-R1���aP ���Q��X�J�S��Ǧ'��ƨh/��Yij�    lUK�"�u����SZ 0�1���8)����G��MOƿ.(�,n��iZ�    �������K��{~�x. `������]1-��r�m���Y1:���M����u   �&Z:�D%-��g2�� �tl,+�ɑ�r��ӧFG�/�ķ���_.w�#��    hQ-L��q��]يib�� Y:&���r�M��dL/�Nߦ����/K�45�   ������I�aI��'G�0 `�c��bI�\n�~��7�1Q�_�[�   @j�`RI麢(=�E<>��/��� �������Ҙո��}�N�后sIf*��Qm;#  Z��#>y�:�j������Y�����˃A���d������| R���6�#��K �ڼ#Ž1=6���D*�m��_$���W��y �V�x�%��(��ɱS>��#�����$͙S}�G�]Z��/�E�����oۄ� �����ruj�$��\���E_��L���   ТZ>��L9�?\>�+�>EL��L꙳6 �����P�z(    �B��64ֲ������W[��KVĵ����    @�"��t�E\>�YEQܒ"���(����vç     h*���f�G�]zZ��?FJ�w潋��E��'�3g}      M%�`R��s�c�.}Oq}��Νs�����#/8h��     @��.��L��7�>���~��ξ��R|�<4l;o�hJ�?N����     д�&5�|�sk�Յ�\w���T��*���m���jW�����S�;��      �Z��d�?���,W,���??~��'Eqr��H�ۋH��s���K�,E������>���     h���^{S��-     @F      {�	     �=�     Ȟ`     dO0     �'�      �L     ��	&     @�      {�	     �=�     Ȟ`     dO0     �'�      �L     ��	&     @�      {�	     �=�     Ȟ`     dO0     �'�      �L     ��	&     @�      {�	     �=�     Ȟ`     dO0     �'�      �L     ��	&     @�      {�	     �=�     Ȟ`     dO0     �'�      �L     ��	&     @�      {�	     �=�     Ȟ`     dO0     �'�      �L     ��	&     @�      {�	     �=�     Ȟ`     dO0     �'�      �L     ��	&     @�      {�	     �=�     Ȟ`     dO0     �'�      �L     ��	&     @�      {�	     �=�     Ȟ`     dO0     �'�      �L     ��	&     @�      {�	     �=�     Ȟ`     dO0     �'�      �L     ��	&     @�      {�	     �=�     Ȟ`     dO0     �'�      �L     ��	&     @�      {�	     �=�     Ȟ`     dO0     �'�      �L     ��	&     @�      {�	     �=�     Ȟ`     dO0     �'�      �L     ��	&     @�      {�	     �=�     Ȟ`     dO0     �'�      �L     ��	&     @�      {�	     �=�     Ȟ`     dO0     �'�      �L     ��	&     @�      {�	     �=�     Ȟ`     dO0     �'�      �L     ��	&     @�      {�	     �=�     Ȟ`     dO0     �'�      �L     ��	&     @�      {�	     �=�     Ȟ`     dO0     �'�      �L     ��	&     @�      {�	     �=�     Ȟ`    �PQ�SJ��x* ����}�
Y�    IEND�B`�PK
     �k�[e���  �  /   images/6c1978d3-8c4d-4ea9-a1ba-37ab4b096c5d.png�PNG

   IHDR   d   0   ��ߵ   	pHYs  \F  \F�CA  �IDATx��{LGǿ��w��AN+Py\0!���hB������jL�6��h������Ķ�i�O����i+MK�6��FKm5)6& ����X�x���3{�	��=�N:������w�7��E'dnݺ5��9���T߾@�I��ڕ������D����	�\���`pA.H��I0��\�����O�&p.� 3�`,(Z'��Duz �v����%HFk0��G�s
49�&�6O�����LJ{f�낈4w�C٠iڛ�o��nĈ�	������W
����,���������x^^.T5�����;&Ռ6�",H�&����$�y��f
rV�oP<��b�D���^�Iϫ��?5��������)�#G��X��.UB�%�~�+�S/�Xh´��R�>��Ȳ��E���"�H%Z潷D7b���3#��P�A�[��}�w���L��R�$�:��ϜGEަ�����9^Mo�#�{ox��*!�Z��l�BOk��p���\HNIa"%@GD�#���6�(P����@��59�꼼�:1�K7�����Y|
oF�&�-��]��J�G��Oh�մxz)#b��>�������������ے	�]��wpbd����F�����?H,����?zoch܁��Q�>c)I�.��(��μ�}u[�}�����T�yj%�C{?/^��f������L�#�ʩ�YF�DBK|p�"��斖���������b�	�Z$����|jkk������!�.$k7L&�����ގ��.444$`o��#"A�ks:����@__233��א��$���鍺�n�#|�7pZ)�Q/kԙ(gϞEii)o�ç�Z5�����!����v���.N�|@�����a�?::�'N�b������N�yͅ�Ҩi����>W�~�F+U"�!�E#++K_�ĺ��,����	�j��(�`Â���F�c������E�����t�jCX&���\��{Y��.56��F}��K?����7�����ڵk��ƍ�	=�ߩ������l�cǐ����%|>+z���^��� V�^=o��:L���~ϡ�$����Ass�>u��ۋ]�v�� �}�-��(ӒN�4Ҭ�X�V466"99Y�h�b��ˢ�,X�������dJ���|}{��ˉ� .��gKs�?U�C�]B�c��]��hL�px�^4�N�<�Ʌ��e;��G�r���C}�1�F��hLVp�Ejmm��-������%w��(/\�����@]k,"�)�:+�Nё�i��#Q/��s�9,'`x�^C�|��:�C3)=g��&-�[6c̻�4j*-a"C� �9�/f�
Ց�Y!��<f�@_�D��2�&���^J��!�����P���]�� D�P4U?��<9QN�p�(nTVV"xߊY/�_��!l)�p\��['��̾�7������7m�2`0!�P�{&G3�(²W[��]m�)�#}l��wLL�®_���To=MK�iĘ�����>�����9BުU�<)�twq�`|�7�4o�k�9�:��a�FR��:�F�.�}k��oDF�3�L}�N�I��Ĥ��Yw#��N�q��V�V��T"� K�9��$\���`pA.HdL���{��X��aT��Z�    IEND�B`�PK
     �k�[�{�, �, /   images/f87b1235-301d-4eff-8a86-0c2fbb955692.png�PNG

   IHDR  �  "   �?��   sBIT|d�   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<    IDATx���k�^�}��9�}� ��%	� �II�(-���K�c���H�5�Ԯ[93Q:cw���I���4�v���4�$��:�ә�M��I\UR�Ē%R�����`����
)��������3�`���|p�g����?�����3X.����qD<�#b8"��6�.!          p��+���ZD|/˲�6�s�oFD=aF�P��;y�dyaa���F�Y��OEDq73           m�jD�qD�a�e055�/�b<=lW
�x"˲�F�OF��n          �(�G�ߏ������_O�4ZVp�'J.\��,���f�y�U�          �οȲ�oNMM����L�ݳ���'O����~&˲/G��;�>          �3��e�955��FD=uZoG��PD�7q�N�          ���l6�t�?H��ڑ����ľB��_E���          ���J�/����R�5�]p߿�G�<���߁<           �2?{����%uv^a�7?x��dY�[ѿS�           n�/"~bhh���#G�����f�@�;��gϞ�r���#���          �%�f��*�J?z�̙��Y��]p���Y__���t�           ܎��y��s���y� l�m����7Q,�ID<ܢ<           ��|�Px��ٳ�K���r�����c�F�#�D�           ܉��<���s�R���[yѱc�*�F㫡�          ������������p�Rp�VWW���x��a           ��D�e?"
��pg�����_���d�           lK�e�CCCť���:�/������T��_���.�          خf�e������A�=�Xp����/
�oD<��y           v¥b�x�̙3󩃰u�;}�P(�z(�          �i�^��Z�ܞ�Np߿��<Ͽ�]�          �SY�=;55�G���57�������          @g˛��WR�`��Vp?x��"�Y           v�{<���!ؚ�Mp�k��          �E�,��3�5ٛq���ӍF��LR*
122���Q(R� �������󱺺�:
   �MU�������Q  ��4��r�J���G�^O�h6��]�p��I��[{K��СC���l~$Uhy����`������`dY��	  ����F,..���\�����   �%�R)FGGcll,��r�8  ����j�����b;=/˲�qjj�3�spk7������������;��b�###166�j5u  ��f3�\�sssq���h6��#   ܱZ����122�b1u  �Y�;Z����?==}5u�ٍ�޳,�K��oQ��cff&fff���/&&&bpp0u,  h�f��ϟ�������L   `G������j\�x1���������  t�����p�AV������_���I�w�_�I�e?�2�����XXXH  Zfcc#fgg��  ���h4baa��J  ����R,--)��-�`(8m,�����8%�m��.  ���]   �� @7s�[���c�*�C���b����A����E�^O  Zbyy9u   ���z�j�  �2�waKj����M�w�GD4���S�N�l6�   е�\��:   @�]�z5�F�  ��VWWccc#u�Y��N��w������A�S,,,��   ;nmm-�]��:   @�5�XZZJ  v���b��Ioc���ă1�:t�+W����z�  �����SG    �5����#  ��j4177�:t�S����b�x"u�4333�#  �����9    =��ի����:  �������c@'�w�=�����q��i���  �5fff��h��   ��� �[4�M�pVWW�K���˛ͦ�M�F#._��:  l��Ɔ�]   @OZXX0� ��077׮]K:N�e����<"�N:���l�����  �r����  ��u��  `[��z\�t)u�HY�M�����1�:t�f�gϞ�f��:
  ܑ+W����B�    �,//�� ��v����c@Gj6���3psyD��juu5���S�  ��V���ܹs�c    $w���X__O  n���b��ϧ��L��M)��6]�t)���S�  ��r��Y�    "��h�����h4��  ��������T���t��T��!��5��x���ccc#u  ؒK�.���R�    mcmm-Ο?�:  lI�ш3g�h��l6�Sg����R��NW��Mu  �#,..ƥK�R�    h;sss1==�:  ��s�����J����<סnSy� �-VWW���_�f��:
  ����r�={6u   ��u�XXXH  ��ŋ��]O�v���R�;w.u  x��d�u   ��Ξ=W�\I  �fzz:._��:@�)�����7 ��������Z����Q    �^�ٌ�_]� ��2==.\H`W(�C\/�7���Q  �q����ꫯ*�   ܆f�gΜQr �-\�tI��)���[���G�^�#G�D�PH ����gϞ�F���k������   p'�����ի;�f�ш�_=<���;�6  lE�ٌ������l�( �J�Zhii)^{����bѧ  �gvv6Ο?ߒ]�j�Z���    wjxx8677cuuuG�m6�155�z=&&&vtm  ��F�aW!�g�@�[YY��|�;����:
  =���������K�R������    �5::�r�%k_�t)�������fK� �7[__�W_}U��Y
���z|�{ߋ����Q  �b��}/fffZ�~��166Y��d}   ��Ȳ,���#�[s�ʕ+���~7�]�֒�  "bii)�����
�4w�%�f3Ν;gϞ5� �w�ʕ��?��^��b�ز�   �+��o��׮]��~�����вc  Л��f\�x1^{���� $�� �l~~>�^�G������q  �p�F#.^�ز��׍��D�Ri�1    vB�\���ј��o�����q�̙X\\�C�  ������ٳgcyy9u���;mH`cc#^}��ػwoLLLD�e�# ЁVVV��ٳ-�����Ù   @G��������cee%��h�q  �n���q�h4�� �wH��l��˗caa!>�  [�h4����1==�f���*��122��c    ����p�����>�jtt48`�;  [���SSS����:
@���5$����  [v�ʕ���������P(���xˏ   �
Y����X\�|9677[z����XZZ�������XK� @gk6�1==�.]j�0�������F�ѷ�����	���&�_�:x�	�  ����z�?>�\��+�˲,���#��]9   @+�y���133�F��Ǫ��q�ܹX\\��F�Ri��  �<KKKq�����2�f�N�ŗ^y0
ygf����W�k߾z�@�+~9"|gm��h���b,--E�R�r��:  �5�����3g����ڮwll�MX   �+
�(�����+�[__������؈��>  ����8w�\\�x��]���'�j��}�x��D<u0��w��#��,˾������9x;whC1??kkk����B!u$  X\\����q�ʕ]ٞ����ص�   �Z�T��7�E�euu5���""���/�,۵c �677���˻>̪Z*į��c11\{���+��C��C���W��Z}�rA�Qpo_
��Ʈ]�sss�h4�Z���  �#����̙3��u��T*122�+   �u*�JlllD��{�f�W�^����(�JQ�Vw��  ��h4bff&Μ9KKK�z�,���+'㑣c�|ݡ���ȣ�����gS���Ł[�.�ۗ�;��f����1;;�F#j���; @�Z^^�s����˗w�F�u�b1����|   �Z�j5�]���C677cqq1�X,*� t�f����7vi���Έ�{����SG���B��CGF�����������M��v��޾ܡC\/����G��4� ��,//���T\�xqW��~�,�b�޽Q(�   `7dY�J%VWW��`Be�^����XZZ�b���[�  ��z����_����$����G���/~���os���Z)>x�@T���.D�a�;�A��})�C�i4q��՘���F��� ��ڡ�~��ؘ�   @O��<��b���&˰�����y�G�Z��6KH  ��.����}���՟x<j�;h�eY?4�ܿ/�ݹŘ_N{�v��{�Rp�u}����\lnnF�Z5m �C,..ƹs�����ɋ����100�:   ��)�Jɯ�����r�J\�rE� ��lnn���L�9s&y�="�T��o��G��h߶��+Ǐ<t �V7��/.�@:h_
��K�:\�ٌ�����������T*7.� �>��f,,,ę3gbvv6666RG���J�###n�   =�R����F����Qnݯ��\���� І���czz:Ξ=KKKɋ����GNē��ٱ�
yO�F�����f��ckC;Qpo_�����l6cqq1���?���CCC�c ��z�sss133�7K߬P(��ؘr;   гFGG���˱���:JD�q-�ҥK133����gϞ(�˩c ����՘������h6۫��ɧ�ď<t�%k�pr�_�����ZK�p3&�C��؈���X\\��! @"���q�ҥ���p]�e1>>Ţ�  �ޕeYT*�XYYI�-~x�r�lg ����cjj*.\�kk�W�~��H��'NF��n��@%�;1zv!�^k�q �ۗ�;t��[���G�e��  �`ee%���bjj*VVV�n��u���Q�VS�    H�P(D�Ph��RDĵk�bnn.VVV�T*�� �b�f3��ٳ1==���#�Ԟ�J��O>}������q���x}�jL͵�á�
��K�z@�ш�������z��j5
�B�X  ]���/Ƶk�=����?S�    h�R)��fۖ�"��1p~~�.�  -�h4bvv6Μ9���Q��SGzG�<�_��#qמ�];f����O��ҵx��ҮZI��}ًv@�V�r����������f������l���ľ}��R�| ���>�azz�m'|��r�###�c    �����X__o�{D���Z�={6.]�{�쉱����<u, ��U��cvv6fffbss3u�-�_�/<�����<�_�ȉ��w�ՙ]?>�;�a���j���ED���F����,�f3���c~~>cbb"���R� ��F#���bzz:666R�ٲ<�ctt4u   ��566�/_�F��:ʻZ__������˗c||<��ǣXT  ت�����������8��������Oܕ��Y�/��B���_O��n���m�T*7��###����Q%����XZZ����ػwo�� ж�Oo���m�-	���訛�    �P(bll,fgg��l���%�z=.]����7vq.�˩c ����՘�������9���X_��GN���=},�f��i�;��4�����,�n�/˲����z�/"byy9����Z�ƾ}�bxx�-6 �^v�ڵ��������;ϻ�ȑ#q�ȑ�1    :�ٳg���;k��]���cxx8����Z-u, �����333����:���
����C�Wi���_~�XYߌ��S�� ]�}��A)�166v�x�X�������K�l�����̙3Q,cϞ=166f�' г���bff&���RGٖ�Ƌ/��F   �-���������^M�5��XXX��������rm �I���1??333����:ζ|��qt�@�o�e_|�XZ݈�}�r�8@)~9"*��@�Ȳ,���s��w�T�F���lg5��z�j������J�y�JŅ/ ��mll���l�={6fgg;�BW����Q*�RG   �Y�ŏ�>��_'�V�Rǹc��뱸�sss����R�p+ �'���ƥK��ܹsq�ʕ���Li[^y�p|����1n*˲x�}{�[����ҵ�q�dY����������e����@�سgOT*[{&dzz��QoV,���?���bhh(
�B�H  ;b}}=�\�����%��dY��Gcbb"u   ����X��_����6���j�CCC188�����  �f�+++������=���`(~����R!O喖V7�~�Objn%uز,�~gjj�S���Lp��044}}}[~}�Z����h6�-L�{�F\�v-�\��������F#J���; �Q��f,//���LLMMťK�bii��.tED<���199�:   @G:���#1<�����:Ύ��뱼����1;;׮�1e�T*�� �(�z=����155�������F#u�3X-ů��c1T+���*�B<:9��O/F}�{��n&��/{��U�����
�B������lהܯk4���KKK155uc�{�j����s h�������N߆���}��q�ĉ�1    :ާN?��s�}�[���z�sss177Y�E�R���������/R �c}}=���cuu�Ə�,ϲ��O����Z�([v�x|��Ư��oE���]��[��y������T*100KKK;���\"rqq1"�(�_/�W�ըT*Q�T"��{� �󭯯ǵk��ڵk7.n������������g�M   �k|�>�څx��t�(-�l6cmm-���bnn."ޘ�~}�U�R�j��� �\�ټq�omm-VVVbuu5��z�h��ǟ��'�O㶽ﾽ�c�=���_O�`
�����*f�(Z����͸z�j\�z�-�/��7.~U*�(�JQ.��T*)� [�l6�^����Flllܸ�u���'���<�����Q*�RG   ��J)�����㿏����qv���F,,,�����y~c����R�t��.� �V4������[[[�k׮���z4{|��ɻF�/����1��g��7��م�wS��� J�����@T��m�3::���=_�Z__�����N�/
o��U,�P(�x{��<�B���O  �f��F#677�^����捷���؈z����Q��{��֭��}���Λ�    ���9�7���p�������$�h4buu5VWWo��b��r�Əy�G�X�b����
�x ��F�����������zm����>~2�sϓ
y_�������/c�k��)��-��ڑ�
�B������쎬׍��̮��m���yY����ͥw� �=lnn�(�7���f��������8~�x�    ]��?��Ι��?�ש���;)�]����{��j ���׻~������Y�{0�m kj�Gj�W>t����ߦ�t �	�-����hA�Z����@\�zu���u�O��� �^������S�    �z�3���T��4�:J�p� ��x�x�}{S��1/�:��;��GߙN�0���zST*�_whh(��� @���<^xᅖ��   �V�j9��/��(�iga  خc���/�p_�;�/���Y���Qp����<���Z�v�e166��m�  `;�x�طo_�    =�����_L �.Q+�~�d�,u�7�_�Ϟ>�:�a4l�&���ZZ@/
122Ҳ� ���S�N��   �s~�CO��?u  ��_:���R�h��=�h��Y�;)��)�J������Z����-?  ݫV�ų�>Y�}�    �]�e�}��|8u  :�K��N�O���,�z ���J�~���Ю�FFF�T*�ʱ  �.Y����?�+g   ps�}����d
n� p���鏟����聃C����c �w��&�r9���sl���    IDATl,�ܧ"  ��G����   ����H|��ϥ� @�)����8�R!u�]���������|��7��c���m!  [�o߾x��GS�    �>����Ǐ�� @��������V⣏J� 
���r9*�J�c���%;6  �%��x��g�   �F�,����W�\*�� @x��H��ho���ɨ�{gj=pg4"��dd$�,K� ����C���H�    ��C�F�?���1  hs�<�����ѫU��r|��éc mN�"�X,F�ZM�a`���� ���#�<�:    ��3{&&�I �6�c�;G������'�:żG���(�CD�ˇ���X�m!  7���O;_   hc�B!~�'?�:  mj�P5��3w�����@9�p�@Sp��eY�Z-u�ڥl @{ٳgO�u�]�c    �.�:yO<r���1  hC�~z2�E�͈�}���qށ����Z�y�>�
����r �6�=�X�    l�g_y6u  ��h9>�Ё�1��ѽ�q��h�@�j�V/$��ߟ:�ۘ� �������   �A�s�x�>�s  ��>��d�Lo��Q�n�WKzZ�X�r��:�����G�PH �6�裏��    �m�鏽?u  ���@%^~�P�m���1X-���!wzZ___���w  ""FFF��ѣ�c    p��~�X�d�  ��O>yW�Mo�R1���HhC�b��j�Z�隷�/�ܧ( @�;q�D�    ܡ}���  H�T��CH�m=wB�x;�YzV�T�b��:�;���  �^�T�{�7u    �Ї�w*���� �e�?8�}��1�փ�Gb�P5u��(�ӳ�����b�  $t�ر(�]�   �T�R1>���S�   ��>~8u���e�<�/u��(�ӳ:a:z�T�J��:  �?~<u    ��G_|2�,K ��?0�J����=�# mF�����y���1��w ��t���M   �m:�w4��н�c  ��Ǟ0�}+N��J!u��(�ӓ*�Jd2%�V�E��T �5���    쐏=�H�  첾J1�}`_���g�����1�6�5KO�T*�#ܖ����  �E�r9�=�:    ;������ �������[��=c�# mD���T.�SG�-�Z-u  v���d���1    �!�B!~�=�� �.z��#t��w��� �wzN�eW*��� �;w�ر�    �ay�é#  �K&�kq����8<��}�5�hwzN�\�,�RǸm����#  �c����c    ��N�}0�9�7u  v�����%�eJh
���R��:���jY� ����   н^~�w �n�eY|�To�jF�zy�&�?4�ck�M���S,SG�#�B!*�J�  �ؽ�ޛ:    -��OEn� @W;u��?җ:Ʈ�V���Hl�Gwd�ɽ;�����9�r9u�;V�VSG  �����chȶ{    �j��`�:v8u  Z���<�ro���U�DD�#'wd=w�:wzN�PH��j��  h�����    h��<�:  -�eY<���(Tzc�{��F!}�6���K�{���W��~�s��)y�G�w��y��� ������    h���`�Y�:  -�бñol�g
���7~���wp��eYġ��m�t��m�������)� t����J   ��S��� @|�7v�ɋ��Iv��	�ת�vd͉a�8@����Z��:  -099�:    ��'O��  �˲,��xDD��/�7�R4��__��P�}D?Pp��tC�=�sS� ���wߝ:    ����<y��� �z����7�Ǝ�Y��8M��o-�o��,n���X�Pp���yw�'�� �]���chh(u    v���@�:v8u  v������dYw��n�Qx�����ȶ��/�������_E�M���^�yJ ����   �{^x�Ļ� ���eY<���7��;zj����^D�(o{ݡZi�k �����d]��_�禸 t�����    �e/<u"�.�	 ��:v8���֎ͭ��>ԧ�(��c���
�  ]b||<��z�b    {G�Աéc  �>�T��γ���྾��
;=��
�Z���<  ����N   �D^x���P  �&˲x���c�F^~�����hf�m�[)��
���n*��y���O  �,����#    ��O�����a �����}c��cs�p��Z����.J
�@(��c�����w  :���x���.    ްwd0N;�:  �Ы��l*7}�8��u�y]V�;t�Z��u�} �^bz;    ����B @7Ȳ,N?q<u�$���&�Gԋ��Z7�"
:q��ܡ��y���O  hG�M   �Ğ{�~C�  :����o�7wlndś����p~(�C��V��#  p���bdd$u    ;�g$�ݵ/u  ���?u�d����;PpPp�W��RG  �LNN��    @�x�RG  �<�����y�	�}���F
���
�B�J��1  �MG�M   �6���[� �T�'�b����1�i�7�m����Y���]�w �����{����.    ������о��1  ��{�!�f�G3�y�����0��&w�
�  ��ȑ#�eY�    ��<z�  ܆���{��,��R�[)�C(�Q,��� ��q����    h3���P �N�gd N�} u�dy��+�ۤ�]�Z���  ��J�8p�w/v   ps������1  ؂<�@O����o=��^�ۥ$@�Rp�.Q��RG  `�9y�[1    �*ϲx��R�  `�{���jd�.�ok�G��D�\�B��:  ���ѣ�#    Ц����R  ���V��O��=�f^����Z��Qp�.R�z� ���y�J   �6�䉻��VI �[x������H�[��Mp�K��H���7 �vv�С(�n=�    ��U*⽧�M �[x�1��4�]
�E=6`{ܡ�T*��s��  �����ު   �w���
S  �T,�{Nݝ:Fr����F��]�t�b� �4::������B�KKK����/_����G���(ݥR����j�  ��,��ȑ#�c    ��y�X���بo�� �yϩ{��ZI#����fd�,T"ۼ�K��n�U�b�O=�T��=�'N����-_�ʕ�����'��+++��Z�V�)� ������V��c    �����x���㏾���Q  �!�=f����ƻLp���̫�+�w�+
�����O}*^x�������z*�z����>_����_�j�;w��i����jdYfw �6399�:    ��'�+� ��B!�<v�m����f�X����.��QG���r���+�c?�c��׷��*�J|���ӧO�?�g�,~��;���w()�,ˢR����Z�(  ��ѣGSG    �C<������cs��:
  ?�ĉ��^O�k�[��^��5p���1�6u�=��W����g>��r���y�O�����ߌg�}v�օ�T��RG  �M&&&���?u    :��@-{�� �vr���#��F���FA��sYp�W��������-;F___|�K_�/|�Q(��ch'
�  �err2u    :�O�H �(�y<���c���
�&���Q�,��g~�g���|��]9��/���˿�0LGɲ,�U'  ���QӶ    �=�=v򎺥 е����c�
�@�u�w�y������ǧ>��]?��?��+�}}}�~l�S
�  �aϞ=100�:    flx ��p�  D�i��Ec�F��I�n�1��~����/$;�<_��T*%� ��V�E�e�c  ����;u    :��'���  ���,��w^��
;p�:����O~2>�񏧎�N��/~�c���y�r9u ��799�:    ���'� H�ԱñgĎ�o���w�5�ε}��ĉ��|&u�N�>/��R��%�Z-u ��6>>����c    С����{�� ����v�0�h��.�����/��/F���_w��?��8z�h��ժ�  	��   �v�~R�
  �,��o&�Ng3ˣ�w!Ѝں����}.��ۗ:�۔J����������(
Q.��  w    ����� H���bb|8u���̶6��w�N�mC�ĉ��/���������?�:��j��: @O��a�    ؞{F⁣�S�  �I/<y"u����b��QPp�L[��<�����k����~*Rǀ[��j�#  �$��   �)�?q<u ���<���-����[�VmYp��;�������Sǀ[*
Q.;Q  �m��=    ��&� ���C{GS�hK��w��ڮ��eY|�ӟNc�^y����On�w ��522��.v   �3O���G��� �S>�ԃ�#��FV���Lp�P����8z�h�[���/��R�pK}}}�eY�  =��{�M   �.����J �gdY/�G��沈-Np�Tp�P��_~��_syy9��� ��կ��˗w|�}�C��m�W	7�y岓 ��r�=���    @����NE�}i �]���G�����1�R3�#bk�V�Jk� ]��:���ݻ7��]���f|�+_���ň��{����>��-��߿?~����7��ck�N���k׮�� ��&&&bpp0u    �̞��x������z�(  ]��9﬙���F��ܙ�z���g���I����7�W�Wo��#"666�~���~��v�8�=�܎�;�Z�F�m��9  �ܽ�ޛ:    ]��O?�: @�+
���S�h[͸��{���$@7k����O?�ckMOO�o��oD�^�����������;v���z*
���ݖ�yT���1  �Z�e199�:    ]�O��J��6j �:�<r,�j�c��f��ک	���j�����h�w�};�����;������F#����[����#���'O��Z�*}}}�#  t����C�    �L�O?|,u ������s+�|�\6�R� ݬm
�=�P������׿_�����u/^�����ߑcFD<���;��B�Zݱ�3  ���17   h���q_ �U��k��#���J�6j�
���j���NN?���l������;r�|pGցV��l� �
�J%�9�:    ]�量���@�  ]��O��ri��{�mLpc�{ֺ,@�j���N��_}����?��-�~qq1�����ȱ�;��'�ho.v �±c��   @�y|���� ��+�>�:B�k�Va=�FA��}mѾ(��q������;���=��nt7@7@�k7A�Z���LI�(�ڭՊ��J�{���$e{�Tj�Nnn���I����8�br�x���)�(7�c�d˱e)�,٤�$ApAb�F��i��^N�/�OK���?��F����#k��?��9?�я���󩽽ݑ��B���R86  ����q�      P!��vY�0  �4�ӦؖM�c?�7����� (gEQp���tl��[o���s��}-//;�ww�#� ��y�f�   �JKK�L�      @���Ԩ�❦c   ����bz{&�&�Ki�	� �W4w'�={V'O���ykkk:z��#:::Y(����|�q   p
��     ����a:  @���t�C�c�;��i�CO@�����FY'���G}�H���fG�
�������t  �����xo      ��=��`�t  ��p�A����*#w �W���&G֙�������ӎdp�c
mh�+  ��Ÿ;      \W����n7  �,<{h��%æ��EQpohhpd���ٜ�;33�H�>���y�f�1   J޶m�LG      @�z�;���i  ��uk�S�z�L�(�����(	�rV?����8�ιs�r~���H�`0��:�MG   (i[�lQ}}��      �P�M�:p{�t  ����{MG()�Ǜ����d�(
�~�3W�,--�����EG28�� nزe�B���   %khh�t      T���c:  @�jm�ׁ\0��l'��=�d�(
�>�3/`���9?7�Nkmm-��@ �5 �X��w  �544h��ͦc      ����ڥ��6�1   Jҳ��Q��(j�%ö��|Qp���xe�z��e�F��t^�O$yg���r�������  ��l߾�t      @���}�MG   (9�j��k���'˂���(�rV�b����1�����3�   Kuuu���3      �$=�o��[L�   ()�ڣ��~ٲee�����U ٣�~
�T��r��~��  �Ԏ;����      ����ы�0  �d�������Q���� {42�B�����khh�t  �����     ���Н�hKk��   %�WܫH��t��dgY;�=Lp�=
�WI$��C��hhh��]  �0�      �����Ǚ�  p3u5=����ey�4�*P �V�U�*����R����k���c   �p8���^�1      �u=�o�zۛM�   (j�{�N�j�M�(YLp�
�WY]]ud�`�T����t  ���w�^Y�e:      �.�e���g:  @�jn��w��Q�lew�Ԗ%ۢ�
 ;�j\��;*]UU���N�1   �Rww�:;;M�       n�S��tp׀�   E�+���j����#��:S�d���U�*���~G�L���Pww��   E���k�޽�c       �ʯ=���[   W���~ݽs�����; Pp�
܁K���υ   Wٵk�jkkM�       2�T_��?u�t  ��QS�����e!�	�i�� I �3
�Wa�;pI0Ԯ]�L�   (
������      (-Oݷ[��m�c   �/>sP�!�1������U���Ҷm����m:  �Q~�_��s�,�2      Ȋǲ�_zF�uA�Q   ��󶘞�o��e�Ρv��0�@v(�_%�H8�w��(��  `�eY:x� �      P�Z���?��'�a�  �P�-���x��V����2mQp�
�Wa�;p-�߯|P555��   �n�޽���0      �˝����6  �u�P���/Vu5���d[9Lp�� KܯB���p8�|P� �.  �c׮]4      pēw��O4  �5�P���W?��M�����
�������Qp�J"�pd����:@�hllԣ�>�P(d:
  @��ݻW��v��      ��^|����ǲLG  (�h�N�ۿ���V�Qʒ�C�	� �E��*Lp6���c�����t  ���x<���{544d:
      POݻK���'��R   �ksT����ߩ���t���ɥ��w ��֫Ppn,�GQ[[��(   ������Ç���c:
      PP������ϩ�.h:
  ��vm�֟�ދ��To:JY�e���a�;��Pp��Sw����:@1
:|��n��V�Q   ��ب�\�7o6      p��m�����7����V  �<|��N�.�s�-+��x�� ;ܯ�w 3�ei��ݺ��{����  ����>=��c
�B��       �ji����tx�-��   �,���?��~��="��:�+<ެ����� ;�j\��;����E�Q��G?�ɓ'M�  Ș��Ӟ={400`:
      `L�ߧ��7>��v����w���l:  @�{���ç����t�
������*���qw�;    IDAT
�@�B��~�a���?�[o��t:m:  ����鮻�Rmm��(      @Q�w�6�����_��~����8   7��z��c�����0��m����ۖ� I �3
�W���nhhHz�7t��	�q   >!j��݊�b��       E���N��o~F�����?��܅ӑ   >a��.}�W����t�ʕ�E��[�  ���Pp�S__�Ç�رcz�74??o:  �<���v���{u      �,��Cwޢ{v�[�����%�R�c  (�ӗ�=����˲,�q*ZN�=TUd�W��$	ٶ��7@J3�t���jkkӑ#G��hyy�t$  P�,�RWW�v�ܩH$b:      P2�������{����?ԫo�Bi�6  T�pmP�rx�>��^>�q IVw��*���q�t:���5�|�}#��H^�W۷o����>��#}��ZZZ2  T���N�ܹSMMM��       %kKk�����K�ߥ������P�t�t,  Pj�z��]z�O���>^Ѱ<��G&����Y]]ͻ���x����L&J����*i۶m�|���ϛ�  ʐ��Qoo�n��544��      ����xB�������]����ZXZ5  ����=q�}��N�j�M��ulY9?϶<�l.��
��Y]]U]]]����~
��U<������߯'N��ѣ:v��Lx   y
��ںu���8wS      
���A_z�>��G?��}�}����j��ӱ  @��z<�c{���w����/��[��g���ƶ��d���uVW���<hqqё��r��ޮ��v���jllL���:{���X  ��������_��ͦ�       �6��ޡ��CM��~�3��O��9G  2�߹I�V=�wHM����<9?��TIi����8Yppc�@@������?�cǎ����m�t<  Pd��������ӣ��vy<�<      ���]���ժ��WЇ���/���|���s�� �"�,ŻZu�m1ݷg�z�dUr��N]@�xŸw����:h``@���:y��_sss��  �~�6mڤ��6�������t$       �X�n�u��X����}��9��1���N꽏�uqq�tD  `@{K�vtk�@�vo�V#��K\����u0�rG��:����������-IZZZҙ3gt���+�L$fC  GY��H$�h4���f577���QV        ���֬��f={��m['���'���������Ri�1 ��j���ժm=m�m�P_��B�c�A���]�=�Ud�W��8U���8���F]]]����{���:��.\����9]�xQZ\\T:́0  �U P(R]]�����D���z�b      (G�R_G��:Z���;$Ik���N����Y�?��?�̙9͜�Ӆ�%É �F���!�E#joiP��&��7��5���zX�9;��Z�Ud�W��0�(������UGG�5��N��������+�VWW��syyY�dR�//hI��Z[[s�c  ��Y�%��'I��������Quu��������T[[{�9       *[��{��~��k�lieUg�47��˚[X�����0����%]�_V2��Z*���K��VI%�R&>  JV0�W��#Y�ꂗ�n��Շ�jը��V�uժ�(RW��p���:U1����~����@�(�_��;P�<����TWWg:
         ��T��5�-�M��   �*�����iQp���_mʔSw����:               ��3��y� 2G��:Lp              ��E��;(�_'�H8�w              P>r����u0�rG��:Lp              ���w .��~�
�~�ߑu               ̣��ܯ�w              ���1�=my��Qp�w              �k�yTNm�	� 2G��:�              �e��\&����$	G֡�              ʅe�Q9�0�@�(�_�	�               �J����Lp�.���Sw����:   (�`0�h4j:F�Ο?����1����&��Ԙ������R)�1P�������l:FI[[[��߿d2�T*����u�        �V��t>��T
��a�;  @�صk�v��e:F֎9��}�{�c �=��"���Y{�W4>>n:JPKK��z�)�1�^:�V2���ʊ������-//k~~^��>��c%�I�Q       @Y�c���� sܯC�  �r���������>y�^&�����,�KR<��1�ǣ@ �@ �����������kvvV333���Q"�p1)        (+�La�PW�9^1�C�  �2lڴ醥�b������E���b1�r���+����g����թ��N����$۶u��9MNNjxxXgΜ1�        �;�	����T
�ס�  PJuz�e�X��{�+�1�ϧ��n������A�e)�*�j��ݚ���ѣG��_�B����       �bg�^pO[^� (w\s�d2�t:��:�  �[)��%���O^/ �U4UCC��y)�	� 2�D�o�>���Kz��K�u        Z�S�d���:�D�k�|>y<|z  �QKK�"���y�<aũ�������|�c p���Ѷm���/衇R04	        !;�	�,ɢS	 3�Z�cuu5�5,˒��w    �V�cI���#`�~� ��E===�c p�eYںu�^|�Em߾�t        Ptr/�KR��*��j�'
�Y   �*��$���0a�555����tGpP���:��{��3        ����.I�x����Qp_�Sw&�  ���E"�1������m:�SN����n~�*X__�>�Ϩ���t        P�v~wۢ� 3���w  ����LGpT9���E��!@��^����L� `P4�s�=W6�       �<�9�=M�@�(����;  @�*��$�����󙎁�F���h:���� ���zꩧMG        F�Wp���;��Pp_w  �����Rvh�^�z{{M���)�($�����m (����ˁg        *�m�W9��y ���
�   �\'Q���U�������Q__�� �@[[�<h:        0��o��mQp�
���  P��q��$uww�����Q񚚚���h:FA��q� ��۷����t        `D~�4w �ྎD"��:�  �Gss�"�����z��]��
I���T04@���{��r        �Jc�Yp��� 2C�}Lp  (?�X�t��*�����s���E ��D"ڹs��        �mV~w�	� 2D�}N��~�#�    �<][����T]]m:F�jllTcc���E ��g�.�       ��Pp�
��H$��É^  ���F���`:FAy<�����Q�*����٩`0h:�"����}�v�1        ��l+��iZ�d���:��  P^*�|,I[�n5�bU�טeYe' ٹ��[e�y+R        PB�=/�� 3���T��	�   šRJ�L�6 �����tW��q� �p8����1        �k�+��y>@��
�   �#�����tWx<�����Qq*ir~{{�jkkM� PDMG         .ɷ�n[TVd�W�uPp  (�X�tW1a�}�r� I�,��>^ 7�e�y��N       ���oA����T�P�(�  ��J+�vtt���V�����T�H$�h4j:������}�1 	�ϧ��vMOO���
PWW���W�J$���~��^�*����ޕ�&''u��YW�      �;;�<�d�
��H$��S]]��:妵�UPSS�B��B�������u��MMM�ȑ#��ʊ��  �DE�Q566�{yyY������qu_˲���W�,����?55���&��չ���͛UWW���W�P����(���pX��ԧ\�kaa���O���ە�VVV(�      � �	�iQp�
��`��󚛛u�}����SKK�M��IR*�қo��W_}U�����t�� �2�Ō�=::��G��^p�.��+����_c����l٢�;w���eY��bz��w]�@�����믿n:        (0[V~�ϳ �rPp_�Sw����:����Y��k��ȓ��E�^���߯����̙3�ַ������ @F�����=22��'Ojaa��	�mmm�����⢫�V�H$�h4jd���U;vL����ܥKQPppYCC�|>��ɤ�(        ���+��	� 2D�}�Du*����������'����sd���f��o���x�	}��_���#� ���F���hd���e?~\�mkttT��~���_����{ﹺo������S:�������
�\�ӦM
�B���wu_�F�������t��y<�+?7[��`0x�WMM�����������lX����f��̘�        
��w��ס pR(�W��ռ�9w���O�āD �u95�=8�N����З��e���d���}�k_�w����_�5�� ��LNo�mے.Mrw��.���b����GFF�����v������e)����vu_�FVWWu��i�1
&j˖-��b�����.i��F)�       �+��N�x<F���#
��n�{��Ǐ;�����:(��nϞ=��W��������z����+��������R��  @�)���ɓ'������:W3l޼�	��D�F�콺��cǎ]�owI��-//룏>�G}���Z�߿_������S��        �=��;/�V��������t�l��E(����������݂�ۯ�s�N�������]�  ���&566�{uu����m���ؘ�9,�2Z�/w&?����J�RW�{ff�ȅ---�Y\\����}���ˎ��Wss��        ����cY^�� (w�בJ������:�Tp����������z����߯�����jkk]�  ���~c{���)�N_�{WOtw��1�����BR��b(�������%	�Q
�LG         ��wۢ�
 3�Zl��	h^��H��m;w����E��E߲e�~��~O>��X  P<L�n�+����hqq��,���L�.�p8llRq2�����'~��E�QLL�Lj��ӧ�ꫯ��������        @���}>w ��bNM?+�)�[�l�o��oE�hhH_�җL�   �566�����ޫ��������۶ml�6Sܝg��=>>�T*���?y�\��F������ �5<<���7Y�����        @aYy�)���pb��T�w�ϧ/�˪��6�{�W4  d��=>>�t:�����
��3�9�hR�m�u9�%Lq��O�S�T[[k:        (�|'�SY�)^-6@���^z�%uww���	_�����j:  0�d��F㙙-..��撖�&l;(�������dRSSS��F��B�����}���F30�        ܈myMG P"(�o������wd�b����C������j}�_0  ��Р��F#{߬|l۶���]L�KLqw��2��Ą���6��'Ojaa��D�466�{�Z���\F�       ��f����V~�P9(�o�	��x<���(��x�|n��v�۷�t  �2��㱱1�R�>fxxإ4ע������!@�t��ؘKi��w�8LOOݿ�����        ��,+�� �d�xʆQp�������k:�M����z�� @%)��$�8qB���.��V4e¶�ᰚ����L&599y�Ǎ��>�:�n�jd_ �:}�����       ��f�@�y ��W�Pp_����3�<c:FFZ[[u�=���  \�D���dd�d2�����>ζ팊�������qY�n�799�d2y�����hqqхD׊D"�F����Z���ZXX0�?w        .1tZ��}`6�U ��b��w��w����t��=��s�x�2 ��� =11�����kj�v<7�o9)�;H�.�+p���5�.ۛ�;        ��v޳΋S��}��(ߒ<��@�w���裏������V�ܹ�t��S�o�  �������Le?~������f}���L��C8Vss���S��&&&2~���p�l��;L3u��b���dl着*c{       PL�t�t��p�ufsN@(�o �H8�N9����/�-,,��_��~��]��;����z���%���Î�Y�(� �M$1V�N&�������&'l��@^�b������䤒�dƏ������b����^---���Z&�Lp       �;�����b����w �1^)6��O����]ovvV_��W�����:��FFF���}M���7�g�Νjhhpt�R�J�LG  �Q&'Gg[>�������1&l�����z�m[���Jsc\D����$'��t        �J�93`��x
f10��Qp� �ky<�ݻױ������:}��'��;���^y����x<ڷo�c���� (&K����Y?�رcZ^^.@��D"jnnv}�R
��i�&#{�R)MLLd���������[���d�.��dɜ��       �$�,�~�ܩ�� �p� ���YǴ��E"����?�S���n�����d����;�V9XYY1  �D"E�Q#{�Z>�m[cccHtsLq�^,3V����T"��t�'N��"
�����}��ɒ9�       �$�X2� lہ5,j� n�W�0��Z�w�vl���zK?��On��T*�?��?s�����jjjY�,-��( @e2Y؞��T2��鹦&l��v_�L~�r�¶��.��� �LN�_[[3�7        �$�Z��,�CPp�	^)6�˔������۷;��m���7���c�����o8��������#k����՜�x  �e�|�8s��q#����i�&��-Uuuu�>_�tZ���9?��;"e���{ RUU���MN�/6�@��������5�B��'�k(�R��zy��5_�r>    �|��5�V�?�
'�Qp�sg=�����Z�������;�hjj*�ǿ��˺��;�{ppP��ӎ�U.^����&�1  �K$Q45�w*����D�Ϸm[���r0Uf��N�:����(�+�LMM��s��(�����n.
i��͚��qu_ ��,���w˲
��D�U[[������(*���)���ʱϿm�J$Z[[��ښ�ɤVVV������e---ieeEKKK�p����� ��x�^544(
)���V�`���|����x.�x��w:��2`#�Jiee�ʯ���k�{~~^sss�x�"K�ϧ��V555)
]s�VUU�|>ߺ�K�RJ$Z\\ԅt��E���ivvVgΜ��Ľ�    (bk�����_'~���� �7�T����ڑuL�����ud�W_}5�Ǐ��hjjJ]]]y�=00����{�r177G� P��񸱽����.����)��b1�����[�L�!`tt4��۶���1��Ɣ�X,F�0�	��RKK�6m�t�W8�R�t�eYW��fjyyY.\����u�ԩ+%�t:]���Ҟ={�~�Sǧ2QSS��^zɵ�����~W��������?��o555���؝wީݻw��_>&''��k����5˲��ܬ��&566���AMMM���/����װL��l���.\��.��?���N�:U��c~�aE"�����|7��4::���G9�_UU���.������]�h4���D�    IDAT�^��ʅ�_��H$t��)���룏>r��f�e��_t�L:��_��_jeeŕ�
)���g�um����y��    �,���c90}�f�;�Pp߀S�r�%gww�#묮��w���y?��)�wvv�F99w����L�   /�\>����i����~Q��	�'O�tu�RSWW�M�6�;�Nkll,�uFFF����2�0�d�}ii��޹
�B���UOO�:::\-P;�r����U۶m�t颃3g��رc+�;�TWW����t��x<E��j7*���aW�깸��[
��sy���������]���N�.��
����q��S��N�:����<yR'N�p���[]��X��#���u�-������_'~�_��������w߭��i���{����{m۶533s������u��Q��+�͛7�zGb�G    (kvZ�2.��NK�J�X< �Pp� �ɩb�|�������g?�ټ���FO��˷//��0  �)��RXO:����x��ض���q:�*;�X��7��
2�2ǎs�g�cǎiyy���Xmm����t��	W� ��E''����U<׭�ު��V�q
������U���ڳg����5>>��G�jvv�t< ��֦���������tGx�^������Mҥ�����5::�����UN��dV����վ}����\�D7fY������ե��Y��'?���t^k����Zp���)���[��洸���~    ��Ҝ�Ԛ����|+&��m�8uP�͉������:~�aNϛ����Ғ#ӑ����>�_�l���ӧ��� @)19�}jjʱ"�������^�u&l�@<7���Ȉ#�ض���1#S���8w� ���}�{ �Ν;u�-��̤h��B!�v�m���4;;�w�yG���� J\uu��o߮[n�E�p�t���z�WJ�w�}�FGG��{����Ӧ�������h4�C�Յ^���zꩧt����?��g��?��un���K�e������������    &$�ϙ�PX�� �7�Ta��c7559����XN�K�Ӛ��rd����~���
� ��e�|<::��Z���ZYYq��?���ڼy�fff\ݷT���iӦMF��<��)###F
�XL���Z�=�R
���J��v�eYҝw�Y��������G�ŋ��o�ȑ#�#�RMM���٣�۷W�+}>��mۦm۶ijjJo��FEߡ�fw˲�o�>�޽[Oq�H޶m�:::�w�w9���|�5������{U0T}}�k�Qp   P��TB���M�(,'
�*�� ��p��^�Y'����ޖ��J=ѳ����kaa�t  �V__�h4jd�t:���	��s�̜�	�X,&ˁ�3�8v옖���v�L�A.�\��zU[[kd����������I���gu��!����z������;v@ay�^�߿_/���n��v�y����.}�3���Ç�}?4�F�]����~�i�q�E[n�,
�駟VWWWN�w��L������Ӝ��o�(�   (g+�OʶӦc�#��� �Rl�	�G��&�I]�p!��9s&�ҥ�>�����  d�d1���㎗�GFF]/S�x�X���������.�@���L�D"�
k�ϟ7������3������MG)	������>g� 2�e������;8ֹ˲400�^xA[�n5�uMp����s�=WR��|>=��9�ǧ���H$
�j}===��U�7ovm�������    ��N%�:w�t80���;��J��D"���R���T�����>�N�(/��4&���0� Prb����QF���r��l�A�'�����ZWO�_�PetSQ�b1ރ.2Y�v��t��۷O�<�H�p[UU�:�C�q�Pd<�8�'�|R������@ ��zH<���^��8�Y��^[[��{�$����xt��a555e��T*���n���A�Hĵ�������^Lo   P�VΟ��N��Qx'
�s�@�hl��mG&|����>!�ԉ�������T�r�'���	 @.�ᰱ�m�+ȺL�.�X��{�'Nhii��u����~O��@ ���N��*�ɿo�O�6�����n�ݻ���ǘ�}�v=��G�Duu��~�i�ڵ�׶,ꩧ�*�A4�J&������ӓO>�p8l(Q��~��x≬��}�o�Nq�z��c��   �\��Z��5���@���*��JqN��=OI�*֩��XϖS����fgg�� (&�Ǐ���rA�65a�����H�)�;H\D��P�e�e-���ǁ�={�hǎ�c����>>|� �*��+��P(���;/塽�]O?�tE�ܯ��~��!E�QCi��u�����399��y�l�j�}ӦM��倂;   �r�|z�2��;Ţ�
��x��������`0��:�N��mۑX�m���/~a:  1Y>.��SSS����F0TGG������Zm޼��ޅ�C�e�.����s�0T����B!#{���Z\\4���zzz��~�1�J<םw�i:P������3�(���R�ZZZ��O���ҫ݃��ںu��4�R[[[ƏO�R���(`�k����习l>�����+���    ���9%>6�=N0��1 Π�~�/���	��t
�?^��Ӧc  pC�pX---F��m��'��鴱	��Tz�W,36Uvff��'������4�@@[�lq}_���r�-�����2��e�`P<� ��`׮]���5�8~�_O=�����MG)���z��M�(��܃����n�i�eY��뮬�3::Z�4���xJ��7/�fz;   �rd�״tz�t��>�� ��H$��S��b��wkii�t  6�Ǎ�}�ĉ�O35a���_?H�>��|Q�4n���J�iӦ�~�����;��kY���￟�/�"˲�������t����u�m���Q0���ԧJ���FZ[[��ٙ��'&&��j_h===���
�    ���SJ�9�1,��0�@h�� ܥ��G�a�{iH�R���eێ� �q&K�n�����{�&l_RSS���ٯf۶+_c����c=����z9P�������olr��433cd����ڸ�����`�Ss�n׮]���6�l8p@�c��ښ"��MG)�ݻwg�ص�5MNN.�u���K�n2�H���(�   (7+�g��?k:��,ˁʩk ({�R� w���ڑu(������룏>2 �O��jnn6��[��T*��������E,3VF8y�
���Ԕ��(|>����\�(w�e�СC�F��2���?7��e���/�2Y�PKK��@�kii����M�(kUUU���{M�(�d2�ݻw������N�B����҂��������sss�+    �)�4��3Ӧc���T��*��Jq��3������c�S�;(�����)MOW�0 @����N���̸v"֍"�z���*~�v��!@�t�Q 塪�J=���m�f,C2���~�3c�K��YF3T
˲�o�>�1��fY���^y<�/���N���������2��,��֭[3~��Ą��d]����f����    �I:��œ#r��]j�9_o[�}^@f8R~Lp��^Ɏ=��g+�6: ��U	�c�҅fN]h���_��kjj\=�5��p������+��gdo�ܴ���W�W�_8�����+��n��V��W���n��כ�����!�����Q1�H���=��ښ��\zzz\�+_nN���   �\����9*;�f:��V����ܶ����*��w
�̶m����ڽ{7'� ƅ�a577�۶m�����_*����DV��ǍM�6-�+��:uJ����7==���U�N��|���6V�J]UU�zzzt�m�����t-,,��7�4�!���T*��g�jaaAKKKZZZ��ʊ��.��H$��K� ,˺r׿��*UWW+(+�����ʗ�ei�������Q����zu�w��QQ�������FUSS�����?22������$�*
��3^.��\��ĉ��    ��^Kh��ϕN���bN�ǫϞ={���d���Pp����Yge��������5���[ڱc����L� T0�����Y�OL)�������*�J���i&��v�&�Ji||\۶msu_���
��J���,K�pX�HD�6mRkk�:::��.����'&�����W^��ۘ���irrR:}��Ν;w����ǣ��f������M===ƿ�����oT�����o߮P(d:FŹ���yZ�,�RGG����3z����R��k�zzz����̕�r������繹9-,,��    ��Jh��/*��.I��g�d2����mQpps�o��;�q� ������oW45 P�L��GGG]�sjjJ�D��TW���~uww�:���A���������訑�{oo�|>��R,�Sss�y��1���x������T]]}��S�w?�����^��$��$	���;z��;~��t:�S�N�ԩSz�����z��ݭ;v����חq���Y���o��t�k��i-..^�#E:�V2�T*�����5��������������TWW�P(d��������Ԥs�Ι�R���t��E���kuuU����m[�eɲ,�A�B!544��*��{2����k�J��~�Լ;~��k{   @!��V5O�]�d�Pp_YYQ"��{ ����\��R.����8���v��~뭷jӦM��  *L(RKK���M��S��&&&�Lq���EQZt��;�:uJ/^t}_SQx�^���P�DA���� �R�<yR�����W&��055�������{�R)���illL:t�"���9����z-_\\��ӧ�~���w��M��:{��+{9�F�Ϝ9�����z׎k��ϗ���.8�fWW���˗��i�<yRǎ�ٳgu��ق|�W���Sss�ZZZ�e�m޼��{���A����F�6-�LjllL��Ӛ������3z�eY�F����նm�T___ट��q걱1�
�Ea/w    ����g>R:U�?�)��7����<�g� Ń��85���҈����Yge�+�J]:��{ｧ���%0 @���ƾ����)K��Ȉ��{OOOџ�wZ��!@2w�4�9sF������(jjj22P��?�?��?˶m���������o}K<����˺���z��#Gt�ȑ����ѡg�y&��3����o�ۮ�Uh/��rN�{�������p��������]٫�����z��4::������-,,hbbB?��OU[[��۷kǎ������V\��ܹsz��5<<|�d6b۶Μ9�3g���7���А��nW��755ɲ���'���)�J�r� �׫��N���|�\X��� �'N��    8)1VK�c�m��ċE.GƓɤ��֔L&�;��� ��܀S�R����t����&���Ą�}�݊*� ����7����$MNN�~�����������A������ט��ywwwI_T���Y}���-���M�]lbb�h��%�I�����FFF\ݷ��F�h��=�r��z]�����y���+�����#G��q���E���?՟����~G�H$���FW�4euuU�����o|CG�ɩ�~=۶�������H��כ՝�������Z===�항���.F���s��    �ak��O�Pn���&�K�n��U 7�+�Ppw�ྴ���:(gΜ�o�al�- �r���)�]f�||y¶	�x�Ⱦ&����C��ӧ577gdoI���R"�p}_�׫��>����#G�����c�I������~�DB�������~�m���������|�������թ�Ǐ�7�񍢝,������ۿտ�뿺����0;;��������8��^~�e������yp\W�6��R�Z�%˖,y�%Y^eI����@�0)��d(2�LM2�� C��	��P���!2���pHbgqbku��l˲d�ڬ}�Eju���?/�խ>��{��_55�t�W[/�>�=���?�P_����{ff��ZgΜ�V������H����-���4�y-����ȋrf��NDA`��*D�=p<��uH?\.���p��q]OODD�)//Oi�x||\I�9����Y�v�Ԑ�J*��*7P j7Q���*�KD�����޽{���K�#���"����z����,���+���P�"���zzz�k�.%�Cu��;vLZ==��E������{8�NM����N�JLL��O�<)dj}0�-[&�V�V�X!�VO!DDDDDd���8݄Y���Vt+��	�sעFGG�g��EܯB�d���X!�`���^#0���~?:;;Q]]���Q��QR�U.�PWW��	��0��n�K��)�w@����ի��(�=zO?�4ZZZT�3/��ggg���,��b������WZ���4i��"��d�����v��W_����ߖv]9333b_�����W^���?|�0�n��Z			!}����ԉ�z�8���!��DDDDDd~�4&ϴ�5p�q����������'�2�ND�`��*D܍za�l6	�OOOs�w�s:�hhh@kk+�^��v��(B$$$`������!|<;;���.%��a�vNN�f5o����t�A���K��7�ٌ���u���� :;;��s���^���r�Ʉ��di�����]#�Zcc��Z���Qs��V��Ҥ];�����Ԕ�Z�x<<xPJ-�Ʉ��t)�d�����ݻ���2;;��ǏK��w �z�ˍ㉉����-���&'9��������+���=t]�1�R{��a�x�z ��D__��B�"�Hŀ�UD�w��S�OJ�5���
���ƾ}�p��q�_ODDƓ��'��b��=������5k�Q3Xyyy�j�a �|>tvv*����ODs:�8t��~�i����P��U����b�H����-�V�����M�5�L��N&YS��n�!N��Okk���)*7Xke���J66�>}ZJ�Ŝ@{��Ii�S���p8RjK�)f2���&���ALt�g�� �/�����w:����9(ODщ����	�v�]�:���%}�I���8uꔡ�=&""}Q9A���]Y�Kuvv*��m�Xt9mN�ݎ��,e���;����+W
{�AD����Dss3v�څ'�|���n6w-D�����~���133#����Ti��"����';���v�ԩSRj-[�LJY�����Ң������{�x<�6��L&�]�VJ�`effJ����#�Q���L�:g�	�ggT�c<�@H>�5�S�N��	�Dܯ�w1aNp�N3338z�(��ߏ�'Obf�/
��(x			J���)|<;;���.%�Un2�ZNN�f5o����122���|�����V3����ɑ^�(�uww�駟�SO=�7�x�N�B �Ҫ�>)ottTj�pɜ��	�D�4���A�%+�i���ze��.������Y�k�k֬�V+2'�3�NDDDDD��cz| ]�1�s�i�ꎌ+�����v��?d��;D��W��;�>�ǃ��v�۷MMMW�@nn.L��%�]�MU�~��Ջ:��������
@�&
�?�h�����7b�ƍ���0�5���i�<���T�144$�VBB��ZD��f�!99Y�:�@ }}}��ђ��lrr�!����z�ol�qx�?����yo�kaժU�X,Rj-�j�Jۜ666&e���|^x��`��!�N�7�[�B�J�SO�`|V�0"2yw�w1w��#d26�ߏ��^���"99���X�|yĆ戈(<*C��C �������j�Z�l6cݺuhmm�ZWkv�YYY��wtt(�}%'N�P�w������M�D���������022���n�������®�hE�w#�F&scy||��ZD�&55Uʦޱ�1�mԹ���0����/�Ʉ��4���jZG�'N(���\�O�[�\n�===X�r���.g�Z����S�Ni^k!�N��nN    IDAT2;s挔:DDDDDD�	��u�bzb^�(`�L�/��3W
��ԏ/����1�لND�À�U����w�U�R���Ǳcǐ�����,_�ܰ+DD$VBB�/_����s�sss����ˋ��{NN������:Y7X�6Q�L&�_�MMMR��_ͅ����PXX�@ ���n=z���W������*=~��9-�w��KII�RgxxXJ-�|>LLLH�x���w=��e�g2z{{���; �]�V?�+VH�%��"""""�s�uObfb3S#��w]�(B@������&}VԌ��*�,�&nD ��1�~^�>�/��#��p�1���)`tt���8z�(�������%K�`ɒ%�9�������͕2�p>ccc�����+	��Z�*�&l�_�^Y��Ǐ+�}5�7Q0�N�&�	�V�ªU���| ���8t��)�����O�S)��~�M��yFԵ#�h$+�.sӋ���ǥ�#��g�x���'N��n�r�aݺux��5��܉����(������0���=�P�$��_������(Mdȝ�.À�fff¾Yg�Za6�wST�MJ��#d�l�@ cccp���\�=))				�GD%Tl��5|���������f�u�b�٤M�O{{���Q��"++�N�Szm"�:�ݎ��rl۶���hjjB@ǹ��~LOO�nC�|>���6�͐׼�����z�	w�˥���W��&J8w�ۍ��dgg�h~���HKKS���d2I;-oll,b{�����H'~��]��v��q����y4%B�(���i;��-CE� �&^k&��b�}���B�ޱ���z�
�GҴO�������>'&&			HLL����n��fC\\�aOJ "��%$$ ##CY}=��gggq��)%�����#&����V"���RR;*7Q�_����R�Q��v;n�����cϞ=�7&�~MOOKy<7�L���R͒%K��1�5�+��8���(��������N�8!%����2����*��N """""c����?;���|�i�gܘ�8�q�>:�t!��C^��Di�R�pCD�0� Q����w3�f�	Y�wevv��)�2�͈����f��b��j��dBL̹����KDD�v�u���[��è��VR;X			X�j���K�.��� ��ǥ��n��̌����պ>%  >�m۶I�����^xAz]�l6+�#�-]�w�u�y晈���&&&+�Vww��0e ���v�u������qi�������~���I���<y2"��YYYغu��ubbb4�~MMMI����yff���~�?��������R6A/]�T�ϥ��J�czCC�.~�D)K�@�,O&"""!�~?~� �Y��l�a�=�r��w�2�?���	�""�`�s"�F�	�d$~���pI���b��{����o����N%����ߏ��KZ`�B8|����"9�\�R����ݻu�;���c�ƍ��feeajj
����k�XIII���H�ٌO}�S��/�W_}Uu;tN����Rj���I���p8�=�x<�?okmbbB����ٳQ�����0��R�����˓��r88u����.�K��Sgg�.~������>�/쯵���:����LcbB���o�]���[o�����Dϙ���P��>�L!}x �M� ��L�i��׬A��ΐ� �ȡ�X
�c�=|Q0RSS�����~mm����r��hllTR���RI]���ʔ��288����B�{�=a�Ba2�PVV&�.-��lƽ�ދ�n�Mu+t����jY�Vi��"��I� "f㙬ǵ��a��U���[F��\WW'���l���ۥԚO~~��:}}}�E�P��/v���gŵ�]���7n��f[�:Ddl�/���q�;���Bʱ��1�����j%u��󑚚���(*C���Նxx<n� ��}�3����=y�jTm#22�w��Z��qG��G2�W����F��Iqq��:�JNN���˥�jmm�R�������	q�����\rr2�����O~��r6oތ��t^�&��K_@4�E�|r�\B�!""��V^^��vMM�!�� p��A��� 66Vj]�ٌ��
�޽[j]Q6mڤ��N�S]]���R�usss������~鵉hq�f3����������U�]�܉�-99YZ�po"��I��CZ--D��\������K�p^XX����


��b�������(xK]�=x�ٌ��ldgg�����)x<�������T������bbbTr�5]�������&�{<!�Q�Z�d	����7R�xn���;�׮��4l����L�N���attt(���R��8�sz饗��%�ŋ��×��%|��_g�NGd�,8)�(t��:�����Di���	���p���(((@SS��.$�k�À;Q�m���צ��� d�@ ���Qtww���cccB�%�����y�{||��u�n��u���(rUTT�l6+�m��1pn⼊�{nn.���188(�v�***��6�	����*7Q0�N��t:�x~!�͆��8X�V����n�+{~źu�p����WGdZ9��(t2����E��\����s�=0�x��bEl����CCCRj�*��w6�u
�Ʉ��T���b۶m8{�,��ݭ�5��ƀ��9�n�ل�À;-���\Ym������^�Wz��d2���/���Ժ�r8ؼy���555�j/��M�֭CFF�����&��������nC8�Պ�K�"==���X�~=���l�2խ]�o��o�w�^8�Nխh�f�!>>����+mFp������x<������2�뎅�EQ�E�)Ӽe~�&����Ǐ�o~�Mk�zNƉ'���+d��)))���k��̉���ڵk����v"""""���;q��.�l�2�|��BMM�!�E�033#d���X!��Ā;ɐ��"���K1|��xp��a%d#�KKK�������ە���M��)�/�����Dz��z��ׇ��>9r����Z�
����Ї>$u�8�ܹ�>���V-&&YYY���FZZ��Ұt�R,Y�III���G||<,KXu|>���1<<���1add��������Ԕ�����J��;wF�棥K�J�e�^tvv���SuA����p�����+��۫y- ��ɑ�~�w"""""��g
q��Q�s�.]��o�G�E}}�nE���EL����6	Qd����w�F@]]������둙����>��'�N�&
܉�s��i�>}�v�­�ފO|�ʯ=�v�m����ǣ��`eggc������ǪU����vx=���Q�����CGG�����Ѐ��Q�{""�D	��7�,�V����[ jjj�O}J��$�����2
0�NDDDDDB|�l�;p�ӂ�,_�o��&&&&T�D5p_@��-��i�����DEDDDک��PVۨ�c ���W6a����v�^w1�nݪ�~]]���᪭�Up_�z5������#�6������_FCC|�Adee)��n����o������b�`�����֭[������yeff"33�\s��^;v������0;;��="�h׊��Oc����ɓ���ѼVqq1���?i^ ���������А�ZDDDDDD�N �&�_(55w�q��ك�gϪn�(*��i ��F�(.j��Q���)))R��]���c�ۍ#G�(�]YY���b���H;��Rccc8v옒�"�m�P�H�cDz��ׇ�z]]]J��馛�֟ϪU�p����?�9|�A\{��_�l6��� ��?�x�	�|��R����p�7��Ijkk��ٰa��uL&��k.��NDDDDDD�
�6w%qqq�Ї>�e˖�n�(*0ྀh��/d��-d"""�L0�ռ$5z�87�^��k�*�
�A隚CO%�x<hllTR���JI]"����ģ�>���)e=���!--MY�����+_�
������[oERR���������������׫n���`�k���h�jH���j)u,
5����)���DDDDDDt)#�'��Պ}�CX�d��V�"�������nZ��v!�0�NDDDWSQQ������ p��Ae���˕������-[��7�	sdM0�TVVV�\��6W�MY��g��g�Q�CQQ������x����#�`ǎ0�B;2Uﲳ����㮻��(Z0@�o��D��gϢ��SJ-��d��ǀ;Q�������_��j�M7���HDc�}�:��f�	Y���Y����"OJJ�ԛ�������DSS���*7'���V�UI���q���)�-��M*���[o����ne�Uܯ��:<��c�x�
��b��wߍ��111��!���Vߌv-�Ē�ɷ���E�������ahhHJ-""""""R+�QC�>�())��Ri��p�{x\.��u���(򔗗�lV�r4R�ǀ�#�/�z�jdgg+�,��ƺ����J�r/-���Ǟ={��/((��o�X��}��w��V��k��<�y@���R�>���j�,郬��			���ӴƆ4]N�\_!""""""�"�^�B֮]�իW�n�(b�J��u�{||��u�n��u���(����G��bvvVIm=Oǵ��غu������ɠjEff&֬Y��6Q$x�w�����v8��ȐV/>>_���p�-�H��';v��g?�Y�mQL���r&�p�n���8}���ZZ�z�p8������jmm�R���������V�Op�SVV��4��5�n�ل�À;�'99Y�$�����(�-��	��\s����(--UL������*7QTVV*�K�-J��t:q��qe�sss�Ա�lx衇�m�6)���[n���2]��.�oH��k��Ś����/���)u������H�Pn�D����$$$ ??_uD���
����
YGQw��#d"""�,����n�^*��ǀ����+�j�*%�R^^��v}}����Zp:�8r䈒ڕ���pJA���嚛���^�r��5�f3���/b�����2�/|�HOOW���Y�Ɵ�:�j�ʕ��z#��z?�����"""""""��ymٲEY��(��j�p��������E���
e�#-|���TMخ��RR�jl6��I��tB����Z%u�/_�u��)�M�MJ���٩�vff��5>��Ocǎ��1
�͆O}�S�� � �f����C������Rk��횬+�ԼH @DDDDDDa�}>���Gdd�R� Q���8!��"j�����E���d(��*��%�өlJoee���WSZZ
�ժ������*7Q��Cdt�O�VV[�i�s


��X�FTYY�o�Q��"���Ɵ�6._�b� ''G������DDDDDD$���W݂T<m�H<^�]@���v��uD}����(r���)8�N���(��5US�322t7a���\Y�:eAp-��Dq�5���q�D�W����. /_�\���V+���/0�x�����իW�n��Ȱ��B���v2lܸQ���9k׮�vO*R����p�.�&�@vv6,��6�"
��.���\.!�Q�P9�;R�ǀگMO�m6�mۦ�~$�0G�&���4N<��Dۅ�`��~���)�'��¥>�я"++K����d���UF�͕�;	���G�:V�[�n�f~~�������CCCRj�>�r/&ڮ���f����n�(�Ĩn@��~?�^/�VkX�Dk���vY����"CRR


��߱c6mڤ���T1*++����V����b���*����>�OY}-���(���hooWV���a�����"55UI픔��l6n��6�k���n#'�Ӝ��|�cӼNqq1��녭'+����*��'�_�ҥKU�@Qp���L�a�ł���ܼp�x<B�!""��PVV�4,������De�#ղeː���'N�nUUUJ��6*++���Q7�B�J�!�d��HIIA__��5?��򹜈��Y�ƀ;͑p/))��l�~'//O�:a�������(������$''�n�(�0����i8��׉�����;'�х*++U�@���Tp���ضm��H������G[[��V����*�m�ل�g6��|D�DD*�<񧧧G�f'#W����ӧ��Ӄ��,M�$%%aݺuB�S���#--M@Wkii�R��������#��z4�9��H,܃ �@ll,�N����&�&����_RR


T�A�����BEQQbcc��'mUTT0�N�333�j�{ޥ���uwR������0���188���	���`zzn����bcc/z�r8p8�����HOOGVV���d}9D$��Si�qtvvJ�Gi���p�]wi^���HH�=??_@7�����А�ZDDDDDD�#��'�G��̼WM$�Ap������&�{<!��񕕕�b��n�4������<;vLY<! �UTT�W��UT^��D�$�`�����[^^.t���z�8t�q��Q���k>%?!!�������֭[�e���H.��M!�t$�����J	����{Y���V)u������H_B���mx�H,܃�����n!���UTT�n�4VQQ�,�n��QXX��6ɑ���������n��P"%�n2�PVV&l�PMMMᥗ^�޽{155%�v{{;��۱{�n$$$��k��Ν;���&�"C�=��,�Q$���D__2335��v�Z���axx8�up'""""""-�2J!��G$�n������Jo��~$%%a�ƍ�� �UVV*��ȷ(�)�D��z��Ո�T�j�*ea���j�w�}صk��p�|�����+���_�"��y����H��L9��(|uuu��0�L(**
k�ݎU�V	���񘈈���(J�p���2Q�pB��cbb�p���;�����reeeܭ�,Y"mZܥxB@t(//�c	Q�D��_,����ak����c�=�ө��������^����-]�GDW&��KNp'
_mm��:��sss��_�����А�u������HBI27HD���� D[�]��v�\�����8J��PUU%�f\\�m�&�.ɗ���M�6�n��PT�E���~�zak���3~���K����6<��üCd 2�^p'
_GG4��u�ְ�#��p���*��Q��p'�p��vDmw��%d"""26R�KEE��	���Ű�lRk�:����[ 2�S�C%2T);���Ӄ����Rk��ĉxꩧT�ADA�"㩫�ӼFlllX�Op'""""""���Ϸ�M�/��	��A2��%"""�*--�x&u���PPP���fi5yB@t)//�/~���Ϊn�����^�W�:f����B�
�SO=%�Y�z�-|���-[T�B!��o��tj���X�V�'K\jff&����M9��H���Z�ܹS�:���8t�Pȟg6�����AG�kii�R��������'�w"��� D[�=>>^�:�DDDDD ��Ѩ��RZ�=..۷o�R����p`���8|���VHgL2���4e�EmDIJJ�:��ԩShjj�VO�?����O~�a�)^��t�3���&k�?�A|����l�g�}/��bP+3��$�Hr��	"==]�:�����/~r ;;[ؽ�������А�u������H�B�����냈�ǷAT�]�	A"����	�DDD����͛7�n�$+++�6����H�	DdUUU�[ 2�%K�(�=33#d�!�w�}װ�eZZZ��ӣ��	��kE��G(닺��W�hPWW�y���4�Z�*�����נ�˵��J�CDDDDDD��%6^�$�p1�Q7d�2�]T@��r	Y��������TZЙ�#))	�6m�R���BJҗ;vp)Q�EMp_�t��u�����K�'���U�@!иzM�    IDAT�&o ]LO���	;��D����J�SRR��0�NDDDDDD2�4]"��� p���x<!��qUVV�n��1a;..۷o׼����֭[U�A:� ��rrr��50 55U�:�p�����VOMMM�[�0�.���cccvr1܉�9~�8���5�S\\��lذA�N.���"��OQ�p����Q&��
���n!��1%&&J��M�SVV���Mk	;}���h�R�r�5k�(���z��#󱾷����Ϝ9��"]�S�}ttT�N.ƀ;�8�@ uuu�����Arrr������˗k��9���Ҽ�W �ߋ1��v"R�� 0�8��NDD�JKKa�XT�A�Ș�]^^����o����9%�����˩>�`rrR�:V�U�:����VK+###:` ��9�~��	�D�U[[�y���ie������J�CDDDDDD���'�(\�!��&��f*Qt�te��w ...��yl6
U�A�[���ظq��D8enfq�\�ji%��t�n����M���Y�֦��|��?��r	��܉�:v�FFF4�STT�����k��_1�NDDDDDDDD2Ũn��-�.��DDD���p(Ցz����Z��z���޾}����ȸ*++Q__��"]���DL���>���B֑p����xM� ����{ll˗/ר��JIIѼ�YYY���(����(y�)��x�~?���q뭷jZ���0��Ӳ&����H�CDDDDDD�!����À{fff��c�����o�E���2�:R�n�����׮���&OII	l6[�R)<<���f3v�ܩ����a��e���bS�
�&CS��|���\��ݍ��H	�gddh^C���$�[�NJ���)uȸjkk5���v�ȑ#W�8�Պ5k�h� ���chhH�:DDDDDD�s&s���6D��q�X�Mp��lB��M4""��UYY���	-~�VkHǵS䊋�����U�A:a2�T��7�x#233�� jz; ���
[k!fsd\*�9�^&�dl�0�Lp8���5M�7�,��5D�Zy%�����ը�����G��c��ֹI���ֆ��Q���w����Z�����ڪy""""""�,�Q�"㮝Ƣ-�.j���ImDDDd,��6mR��Dqq��]QQ��M�d|��Osx�����t�s�=����𰰵D���H������VKFX�n�k��tE��Kd��%&&j�~�אϜ9�Q'3��X�r��ZZ���w!��;dL~�_���.URR������k���;�ǀ{D܍2=K�4�po��1���EL8��g�ۅO[g��.TRR�AN�P9|��_��߄���I����J�IժDZ�:!!A���=]Q��o-�����p�`�$�d�)�����X�|9�����1yyy��0�NDDDDDD���!&"�p1y�h��.��po��1���)���{�addDizTUU�,�VQQ!���jEqq���������VV_��m<�Z�(**��'ҋe˖�+_�
V�^�� b��^�W�ZINN�VK+�C� �*���EӐwRR�fk���xX�/��-cb���!}�̀{AA^}�Ui���|�ri�dn�"�jii��Ą��%%%������L&)X088�y""""""�,�Q�pB��EMz�w""���p8�u�Ve��^/�q����b��7ި�vqq1�v���Kaa���G����se���l6c�ƍʂ�UUU�S�2�͸��k��|FW�f��M��t�,Y"��VdN9�M�Dq����rh9M����hX�/����4{@ۿ�����a��n)�n!..���m�S��~�����QWW��o�Y�:EEEx饗��o��sa~""""""�sLA$�D.������������Q�&{�z,/_ii)bb��<|�0�W�2���۷Y���R�:�USS���^��~aS����P�	��v�4>>7�t~������tn���nak�;�:+V����z=��M�i�Z��W�\���ccca}����Z�ccc5�����|�8}���ͦ��peddH��>44$����@6l@bb������R�]�� !��bccq�T�DL��'�q"""҇��
�������׳��f��KUUU����jU���|8x��z�r��jŎ;��'���p��� w�y'����������A�	Ћ199���a�[k!���X�t��zZؼy��4355%���'�h��
��P��;%%E��

`�X4[��붶6��\�Ν;qmz>"�K���ٳR�q���hz�pm۶���dmjc���������8���$R7^�`����~�L&�����(X��*�f��ZDDD������-[���z�x�����;�ߏ��j�v�mJ�o߾v�=�I��������
Mcc#�N���zw��Q"==]I���
�۷OIm҇%K�(�h*��~�{�$$$ 11���HJJBBB���4ڊ���"t���A��-d�ƍ�}<Q�zLk�^�V�UJ��+Wj@NKK�ڵk5Y{N����IA�,,;;[����$9::���kmmŝw�)�����䠬�L�;�a�Xp��7K�)�y��kn�7ިi���b�߿���p��)��{�DLp���8]���ㅬ#�c"""҇;v &F���Ç�5�TܭV+JJJ���.z��U�pu�@ 555عs������HHH�>ݗ�c͚5x��T�A �����7::
�ϧ���6�~���#..Nu����Djj��Z�W��l�n�	f�v�k�|���P�|NMMM��y<..�^{��u/��ۻ��kkk�����w�B����Ǐ=eCk��G���&�&'�S(jkk5�o߾�>����9�X�BӺ����DDDDDDDDD��s�<�
���&�����E��㚚����رcJ'�UVV.�s�V��7����� ��`�X�c�e��诎9"t=��/5�YRR���$i�D��l�6�$3t�i�&M�MJJ?�aM֞300 ���2'����;��C���tww/���n7:;;wse��ɸ���u�zNvv6>�OH����144$�&ۑ#G4nr8��˻�����l�immռG ��?6��͇� EK��f�	Y���Y�������p`�֭��{�^�����.*,,v��b466r2x:::��ק�~UU���Dt�����������%|�+�Z���;�����6�\���i����PPP tM�Ʉ�}�s�\_H��țn�I��k֬��w�)|�K�9sfџ+{:rAA���o�~#OZZ��oH����ׇ��Y�5��|><�y�K7|���k^`�����������a�=H��B�ъ�	�.�K�:DDDd%%%���QV����|�$�������,�s���w��(��y�f݇��"�V�'Nh���q�X�n�Ԛᨪ��m�ݦ�)d������`�X��e2���OZ��p�s���t�m۶	=�'##_��W5������ӳ��W��|���x��Gu�9pӦMx�G���&�����2�/��(=��������Ȥ�"�"�)Z&�����v���CDDD�PYY��~mm���Fr��ɰ8�ZL��j�.:/���|�b����j[,���*�OD�[o��ɺ��횬{%������$\�뮻��wL�踱��	W����/}�Ka�������H;���3�5|>Ξ=+���}�K_25������w������u�eGG���穩��������������j��å���q�}��?��?�������Ǐ+�K�����өi���ldff8�:E�F<�'L]HݘM�������¹�CDDD��p8�e�e��^/��!�����?�q%��n݊��DLNN�9۶m�s1�9���)e������O�ƪU��ԯ���޽{��&�v�O��ɓ'5Y�ĉ���0���jX�l���o����D_�ݎ��;j&�����^����W����?���zx�ޠ?7##�^{-n��va''.������M�Z�����2��v|���믿�ݻw����j�b�֭��;�i�&���� �;＃��[@7�۰a6l؀��	:t���hii��А�����ؼy3��˱y�f����ijjRZ��inS�u�]�i���"�޽k׮����ڪy""""""�\�@@uDdp�)Z�.�r�;Q�())Q:��.�KY}#:p�����܄�7�x#��)//װ���8n>�8p@Y�}ӦMHNN������D�lϞ=���v���с��\�j�gٲex�������#FGG�֟��f�M7݄�;w"55Uu;�uuu!H�X�b�
����x<hmmEWW����r��r�0==���X�l6���b�ʕX�v-V�^-�O �����Ą��N�<��۷Y+Xf���z+n��V�:u
'N�@?�N'����OIv8���Gff&V�Z���|%�"����^��w��'?�I�'1$%%������_ p:����Eoo/155���ILLL������;;;{�ڹ�f��b9���b��nG\\�V+�,Y����X�+W�DRR����JΞ=�dE���:��۷o��ݻ����i�9��eB�~ŀ;��� 1��̈���GEE������J�QOON�:�$p���	6�n�XPRR�qGW�����Р��Q8p@YH�l6���������D���r��w�մFMM��;p���n�-�܂Ç��������Cjj*


PZZ��۷K��G���Ê+�Է�l(**BQQ����9��رc��Z�իW+{��@  d���� ����u�V]��p8�����qW���z�-��>|n�[���M�6�f�!//O�s���!""""""""��A����N��=��u���H��v�����,<�����߿_YXh˖-HJJ
j��m��p8$t5���&LMM)�oT8qℲ@TUU�D��ڵ��Te�����ӟ���	�����(.. ����̙3����������SSS��������=�����篗�M5�c�Z������$&&"))	K�,AVV������&��չ�G�*�Acc����?����,l�H���)�Ԙ�_~YW�h��~�-��y�^���{��k4����B)�El�!"""""���TvNp'�p1�$Np�DDDѡ��V�UY���F��t�j����ۿ�[����ٳ��VVVJ���jjj��7���je�6 55###J�E������+��B{{�����HIIAJJ
6oެ�����ֆo�Qu�466&t����Dww�������;�[������Q51]ON�:����m�����hp�{�G�Ʒ��V�kQdS5���"G���C�r���CDDD�V^^��>�ǋ744�'N(�_UU����M�U����08p ~�_Im�٬��(�<��s�,��^�R����������Хw�y>�O蚵��B׋>�O���_��W�l�ȫ����� ��������5]�DDDDDD.^�"�p1�$Q7jccc�����&d��-d"""�/�͆m۶)���q�8��vAARSS��1۶mCBB���.��҂��	e��nttmmm��WTT(�MM������oK�w�����I�gT����C�z�t:q���m�Ҿ}�����5����������ǹ�W������)zy�^:tHua����6������H�8���db�=H��z��/d����z����Z���766��t*�	TO�.++��Ǩ(WWW+�	T����M7$�VSSS��(�����ᥗ^�VϨ~��_E��U>O_���	�O��n__:;;��kt��5Y��'��&K�~���;��(N�hiiQ�E Np'�p1�$Np'�E���r��j
��ؘn'l[,���H��b>���G������*�m2��DAD����CCC�k�۷===������;＃��$խh���###��Еg�}V��w�ޭ��Ft�������~���tvv��7�T�E�C�~ P�o�#""""""""c`�=H�2��n�Y��r	Y������f����PY}�χ��{OY�H�r����t��y��֭[��� ���jnn��L�����Ԥ�~ee���D��w�����@���x�'�����׻�{���v#11Qu+��z�x��U��hoo�l�w�}}}}��o4����4]�����UH�������'$���4��}�m��w""""""""�܃Ā{h�>������nǎ�Z���766bjjJY�HR]]��	�W��.C$+�*7Q���"##CY}�H������_T�C{{;��󘜜Į]�`2��������ٳ�S�q��3�<�i�ߏ?����0�}��i��`γ�>���:��D�g�}�۠d���T�E �PHD�b�=H����vY���������t:q��e�盰m�X�c�ݜ���Q__��~������̌��W�DAD������^P� ��^@[[��6t巿�-&''�Ţ�������'���%������۫y�w�y��S��u��Y<��Rj��~<���hll�R/�TWWs�i���vOI����-���T7@DQ�� 1�Np'""�\6�۶mSV��󡡡AY�HT]]��vnn.���/��-[� !!AQG@ss3&&&�Տ4�Gin�MD:�ۍ��G�	��������=tvv�nE��o @TLo�s���ݻWu�444`Ϟ=Rj���?�ړ�|>�q��=�^/����|knnƏ~����Cڙ��6����V�-`�=h�p7�L��la������ztDDDDzTRR���Xe�����6T���M&�e'����s��e�׭[���e��"Aww7��o`߾}�[��������=����nE������p���~���ې���������5GFF������R�������Ǐ�^�����î]���СC������פ����-,
�DDDDDDt5�:ED21�$Q�=�ccca6��+!s�ɧz�Qo�����C��տ�w�b����DY/~�uuu��G��*}���q�Ȩfff��/����ӧU�sE�����׿���&խ(188��|�;p�\��-))IaG�y<<���8y��V�9y�$����*y~}�����c����I���\���w�Q��o~�<��<i(���
����[��^�.4�F����n�������"�5Q�pR4Lp���B�a����(r��vl۶MY}�χ��e�#Yuu���999��� l޼Yi(�����!x�^<xPY}܉B���QSS����>��!�Y�����w��W_}Uu+R���⡇����E�mw p�\��w����6խh����Ƿ��m8�Ne=���������Qփ��?��nN�hhh���˿`����A���<����/53H=�ǃÇ�n#$---�[ """""""":�� EC��f�	Y�aDDDY�����~ss3&''�Տd�'l��� ***�� �� -8p@Y�իW#++KY}"��x<سg����?��7������'��7��M�9sFu;�����׿�u_�ߒ��t�������o��矇��Wݎp>��?�<y����9555x��q��)խh���_��n�����q|���ѣGU��k~������~��׫n����NkmmU��y1�0
Qw�������Y'�'7E3�S��.�$^����k�ԯ����'�رCI}�\ ���>|���HLLTR���/�����Dz��ގ�{����&"Nekii�W���q���;�����%�FGG�����U=�����/����V�s�=X�n�ꖄhkkï�kttt�n�"������w|�����.l��J�/��2v�ڥ�,�?��z���    IDAT�6mwމ��B�L&�m���Cuu5^~�etuu�n��X}}=�^/�V��V�;�	�A��|��|�X,a���	�v�]�:�p3����.g��QXX���������ՏPp_�f���:$%%)������+��|>�����~PI���*܉�?�ۍ��V���{8t�м�������_�+���n�����������8�N���kصkׂ�^T>��EKK��կ������{�GWW�}�Y:tHu+W4==��{���:>�������5�+�z�x�����/bbbBu;AkiiAKK�/_�믿�]w���U�����8�~�m��/���62�ۍ#G����Xu+:{���N�!""""""�B�4섈��!���{�yLL,|>����u�w""��TTT��4���CM����Q��[n�EI�9<!@{�����YYYX�r%�����'R��񠳳]]]�����nM
�ǃ���/x�װq�F������K�,Q�Z�:;;���o��7��Լ��d��2�@ �������Ǎ7ވ��
aC��r�P]]�}���رc��4::������3�<�k��7�prssU������۷�������vm`` �=��{�9�[����شirrr3=z1P__���;v,j���8jkkpoiiQ��Ep���;p.H�r�t$���`����(RUTT(����TO�^�v��� �����Р�~�hii���RSS�ԯ���s�=��6�h.�N����u:����1<<��g�btt�0�X-��~477���O=�֯_���lذ����6w�������MMMhhh@OOO�k0�~�cǎ�رc������<lݺ[�lANNbb�^"������Fss3ZZZ��؈���=���vcϞ=سg�,Yr�{�y�f����nN����hmm��Çq���-	w��I�<y `�Z������|���c������s!�׋��N������ٳgU�EtU���U�\�܉�����(��@D2�����LOOYG�wQӫp'""�LO<�~�(���R���K�d�Y���TwW�����&	v�E w���� !�`�$@Y�B?P6\l@�	EH��"!)B!�����?v���;3�k�LOwW�:u9�����=Uuޮ˩�G�d�T=��n�fb�z����.>��,��,ˢ�������ώ���u��4��$~��~/Z�����x=��3�;��;˾F���7�;�e�V6�d2�g�}6�}������Ȳ,~�~ ���w�{��x���?��?���9s�����7o�yCµk����K/��/�\�������la!�͛7rN*��8�y�x�g���bkk+Ξ=�}�{���|0|��8s�L���L��z4���~\�x1^}�ոp�B�?>^x���s}�ƍ�җ�_�җ""�ĉ����7z�x衇��w���w�#Μ9��죣���ۋ.ī���ϟ�W^y%Ο?�Q�'��o}+���o���<��]�zW�={������wũS��ԩSq������Z�=��������ߏ���;���.]�󿽽����}�\�'�]�|y!�0������G?:��>��O�{��c���=���;  ��`�P��}�6'���&��Z��I�� ����m3���K9���p)�X^K��,KQk����|�r\�|9��7����N�w�}��v#���t:��v#˲���z˅��$z�ޝ7Q���(�2��~ܸq�X����;��M3��q��~bP�ۍ'N���w:�;���j��{�ޝ ���(�����5���ӿ���Ν����y�������״,�(�"�֭[q�֭�oi��(⥗^��^z�-��t���S�NE�ۍv�}��v�N�������w}��`0x�k�h4��`�^/������~m��i4�8>����w�ka�]�r%�^����    `���ྊlp   x��p{{{�����|�˂����ߏ���e_����x���7��<����ԫs��-�,   �\�� �d9���R��(�Y}�Ʃy	�     f��?��=O�   �*�Ϡ��k�\��     `v�ܟ~�酞  �:�~�{UU�x`�g�*p���M2'�T�{QI�      l���Y�Y�/_��W�.�<   6��HA�>����n7ɜ^��d     ��h����~�ܹ��    ��Ϡ�{��I2���'�     �)y����^�yO=����  `�Y�,��}M��<O2�(�$s      6ŏ�؏-�<�   XU��e�dΪ�6�     ,�"��/����v   �/˦{\e�;���}Mܻ�n�9w     ��Z�x��߿��zꩅ�    ���`0$��n���I-��$s��H2     `<��#q��酝'p  �dӮzx��
�Wq�{�eI�5c4%�     �f�ٟ�م�UUU<���;  ����#p�AY�I�bྻ��V����~��      l�����[�Y�ϟ��7o.�<    ���}�6����$sR�t:I��     �����?���|�Ʌ�  @�L��=�lz��� Uྊ��<O2�(�$s      6�?������'�xbag   �<�3hr��j�{��K2     `��/����*�2�~�酝  @sT����K�>�&��n7ɜ~��d     @ӽ��zha�;w.ʲ\�y   l�j��.�3hr���y�9EQ$�     �t��k������  �f���K�>�&�N'��     ��}�{_��O���Ϋ�*{책�    ���@�~ow     ���eY��o��B7ڽ��������   h�Y�/��@]���(�$s      ����p��O��B�����    ��Ϡ,˨����&�6�     ���g���>�����_��_?    �!p��d2��hT{N��Np���<O2G�     pwy���?���v�=��_�.,�L   f���Y��=�� p��`0�=��j���N�ۤc�;     ��i����������o�g�_\��   l���������R����I�"p     8��w_���Q|�X�٣�(}�х�  @�L���Ե���������a�Y)�     �{�������<��R�������u��R�   �y�g���y�'�#p     �8{�l|���~��K�\�/��/K;  ��d�;P��}FMܻ�n�9EQ$�     �
���c4M��S�N�����ć?����>�V�o��^~��8w��R�   @3Tղo l�����w:�$slp     ��~�������q�ʕ�y�fFY���yt�ݸ����G�|p��}���^�    `f��e�dΪ�y�'�#p     ���ɓq���x�G�}������W��e_  ��ȲY;Ã�b�����Rmpo��I椒j�{QI�      0��~��1�}    ���}F��U���j��ܧ,���	n     ��.^�_���}    ���}FM�ྻ���#A��~��      P�����[J  @bղ/ l������=��$s�      �����W���e_  ��b�.���3*�2ɜU
ܻ�n�9w     ��������˾   Md�;�@�5q�{��I2G�     �<����cooo��    �Z�3J����$sR��<ɜ�(��     `6������o���k    @m�����z�^�9      L綾^��������y�   �,��3<�.�3jb���v�̱�     `�n޼���'�w    C�>�&�y�'������     ��n޼��{{{˾
   �SÀE�^��MY�I�R���t���     ,�իW�O��O��ŋ˾
   �A�e�2P��}FM��.p     X/��b|����ׯ/�*   �&��u	�g�*po��I� p     X}UU��?����g>��p��  ��ʲl�W ֜�}FM����y�9EQ$�     �ݸq#����:��o,�*    p��3jb��j�{��K2     ����~���k|�s��i�   ,�,;�mp��Ϩ��{��M2ǿT     H����������>˾   L���e_Xs�51p��<ɜT_     �M4�L��g�������/��QŲ�   �k�h�w�.�����aL&�h�Z��R���t�̱�     `6{{{q�ܹx���'�����e_	   j�u	��P�e��;;;�j�b2�$���R�^/�     �U�裏��������q�̙�������ӧO�ɓ'��QUUܸq#._�W�\�K�.�ŋ��矏˗/�_    ����A��=˲h��+�ђ��U�k     H�g��g�y�?���'O��n��N'���"��'���(�2ʲ�^�U5�G�  �:���K�>��`�d����JD�uc��ۛGV�     `Q��q���������    ��Z��Q����n'�SG��Jr��`��$��         �U2�'����%p�C��˖�y�_L��~��          �L��%p�C��N��dNQI�          �K��%p�����lp        �f�%Z�u	�� p�^��d         ���@]�9��,��         X1U5�C�@]�9�e�dN��~��d         ���@]�9���f�^/�          `s	��*po��I�ԑ*p/�"�         `�TS?�w�.��ʲL2�I���~�9         ���u	��Ф�y�'�#p        �f�b�h]��%p�C���w          ����A��fw         h�*���jIS�z���A��fw          ˲e_Xs�94)p��<��;          P��}M
�Smp/�"�         `�TS?�w�.��ʲL2g�n��d��         ���K�>�&�y�'�#p        �f�b�h��ڼ4����p��潊$0���         M����p8\��Q6�U$�T�{��N2��n�[{�d2I��         X_Y6�����CZ�94e����V���Ԟ3b2�$�         �r���M��~xx��+@�lޫHM	��<O2�(�$s          �ͭ[��}h����q�F��s��w��$sz�^�9         �z���׮][��Q6�U$�[ܷ��bkk+�m���t�����I�          �-˲e_a�\���+@���T�e�9����y�9)b         `5eQM��M��~��U%$�Y�"	�z1Zf��j�{��K2         Xo������_��q�sjB���v�����I�          ���lp���h/��ⲯ��9�"��
���v�9���<��;         4�,K�7i������d=)�=�95a�{��I2�(�$s         �4��M	�G�Q|��\�5���s�O��K2         X=6���O<���c"p�S�<ϓ����I�          �g���j5?M�~�z<��S˾4V�_E�I�T܋�H2         XE��M܇�a����{L&�e_�ٯ"�H��=6�        @se�<6���륪������˾
4��}NeY&�#p         VZe�{D�c�=���w�}h�澊3ܿ�(�$s         ��3}�~;po���{,Ν;��k�F�^�֕��c�;         4W6S��eYT3l}_e��0���/��$p�S���v;ɜy�y�dN��K2         X�V+&�ɲ�Qۍ7�_�B���/�*�Q�sJ�7a�{QI�          �'���[[[1���.�0���'��o|���a���Ԅ��~��d         �z�����V�nr���q|��ߎo~�qtt����������&�I�e��6         �jjv�~�ڵx���_��V��}N��ooo��v�oQ3�3         XY����U�'�I��q�֭�u�V\�z5.^��^o��^G�>�u�Slo��T        ���qn��}<Ǖ+W�ҥKq�ƍ��ߏ^���(��q�s��!p����6�;         �zu������s��+��"d�#p�SY�I�,+p��<��;         4�b6�gQ��ϿO|����?�`�	���ܻ�n�9EQ$�         ������w���S���{�+1Of~>��9�{���t�̱�         �-�f{�,�{+���7��:�f>h&���R��v;ɜY�y�dN��K2         XMՌܷ���Sw[����W⁝4M&��9�eUUEV��B���(�$s         �f�f�{wk�x�J��.�F�:��3 x����,��s��v�H~��~��d         ��f�wvv�����(~��eq;pW�����j���B~�         �t�������?��U�3W��֨��א"p�����M2gy�'�#p         ^����<}�m���n�5�s���v��)�"�         `EUi6�?����C�!���5�e�w-#p�t:I���         ͖e�=~{{��?��CE�l�<�y�5���<ϓ̱�         n�&�n��~(���#�&�.4����u�Smp��zI�          ����p��ڊ�uk���v<����;�w��	�kH����$sf��v�����I�          �)��C���,{C�~���;�ew��	�kX���,�"�         `U�����7˲x����xf�;p��9p�t:I���         7G��Z�~�̙��٩7�(��9p�v�I��z�$s         �U5��ӧO�(�;���5�s���y���8��a��          M�Z�~�ԩ��h6��"p��,�$s�������V�9EQ$�         �ʲl�������z�B���v`
�Rmp�]J���v����zI�          ���#Lo�ۑ�yd���I�[M%p�a]7�w:�$slp        ��c�{���ޥ����7�{�6�/:p��}�!p         ��鼩����l�{����������         V؜a�;��7�y�	܁{��P�e�9�v;ɜiu��$s��~�9         ��ʲ��w�ĉ7�@5����5���T�E�d         ���97��C�^ú�N'��        `�	�3܁)�k������%�         ��,� �;0�{��E�d         �ª4��!p�A�.p        �����p�lp� p�a��^��d         ��Rmp�	������,��Yt���y�9�~?�         `��
����	�k�1�k�i��	n3�n��dNQI�          ͗	܁)�kJ��}gg'Z��}+:�N�96�        @�
���4�5�$svww�̙F��I��z�$sVQU�E         nK��U�4s�F�״��{��EQ$�         ��TKc���5mr������YE6�        �mي��M�^����&�        ��R-��|�7�{M��gYy�מ3�b4%��j�        ���҄�Y���M�^Ӻ��v;Z����&oo��        ��$ڼ^���M�^SY�I�,*p�t:I�E�dΪ�L&Q%z�         �5܁�הj�{��N2�^�<O2���%����c�        9��    IDAT�Tܳ��&p�)Uྨ��n7ɜ�op��        @DD�j����5�e�d΢6�w:�$s��~�9�L�         �%�����5���T�lB�>��}         X	U�8=�,��M�^Ӻ��n7��;         l�ܳ�L�N�^Ӻ�N'ɜM�#D�         p[�8=K�h>�{M���y�d��         6H�`�z5�?h<�{MeY&��n��̹�T܋�H2g���e_         �ab�;po���m�{��M2gS6��         "���[!p�M�^S��
��<O2gS��;         DU?p�j\�x���m�{��I2�(�$s�A�71         ������4����M�{�^�9�@�        ��K�g6�S�ה*po��I��K�����'������h��k         �z�L�}`�kZ��=��$s��H2g]��        �&���qz+���	�kJ����&�s/6��'��         ��xR՞QU�7�N�^Ӻ��n7ɜ^��dκ��*��Ჯ         K1׏ӳ[����^��ݺ�y�'�SE�9�,����Y�5         `�n1y�~��������o��o,�s9s�L��_�ղ�o p�i2��p8�>/"pϲ,�9��0�;���`0�n�Y�-�*         �0�Ɖ�?���{D������0��m)1����4AY��glmm�����n�Z����~?�m�S���         ���I\�qU��ӛ���H=��N��d�&�EQ,�
         �0�c<�"&U�YY5Np#���	�
���v�9o%U�ɑ�d2��p��k         �B|�����Q�������	l��^��dκ���        ��q�f/���Ka�q���4�	lZ������YW��0F�Ѳ�         ��K�w���&���4��=�u	��<O2�s_         �m�Gi���d!p�M�����6��S�eL&~�        ��^�t�?PU5'V�՞l�{����         @�ꕱw�x�֌�o��w���	�e�dκ�EQ��A`0��        @�i{{DTu��Wz;`:�lp�\b         ��7�国��L���Z�6��=����        �&y��q�e�57�g���#pO U��n���y+y�'�#p����|=         h���A\�~tן��z�zV�����'P�e�96����`㱏N        `�={�Ʊ����'�.��ǧ��-�
         0��7{�wP���WUU� �;0%�{�������y�9�7�1�}         �YU�{{{5��g!p�#pO`]�n��d����lq        `�r�V�Z�Zo�{f�;0%�{��w:�$s��?�d����d/         �"�Ɠx����?��@#�X��=��$slpk�~?��޻�         `Q^�t3�)���l�lp�%pO�,�$slp_���          X�2^�|k��V5u�;0-�{����j%�_�e��>&��E��h��         ��TUO}�ZL�-f�Zw`:��!p��<�,�=�v��-�
         �se?�{��O����w`J�R��v;ɜ���<���t�㱯         +�_���Wo�������=�S�'�ܻ�n�9��������˾         ��S/_��d�`���ԳJOLG���:�6�/���Ѳ�          w\�;��[��ϫjn`��w`:�˾@�ØL&�j�{�@��8g/+p�t�R|�s��=g?�m�7��(�c��        �4��8�}���Ϟm����.p�#pO���(˲vļ��Y�EU��E�.:�N�9�
�ϟ?����k�y�;�y���������Nlmm-�\         x�o�|-�ќ���f�>�{>�1���`P{F�e�n���ͺ�n�9�
�����ᱼq         ������?X���lp�$pO�,�$s�k�x���)�"ɜM3����-�         l��� ��F�U�@]�LK��H����w:�$slp��`0H�F         ��xRœ/^�I��u7������=�;�8::���/�         ,�S/_�������n�6�`3�I����$s���}5TU˾         �����x�(ɬ�����q�{ �'pOd�7��y�dNQI�l��x�^o��         ����x�����g5�l�{"�����.�N�(�d�         �땣q<���O�d3�I��=lp�#pOd��n��dN��O2������F˾         2��x�ūq4HۧUU�X~���#pOd��<ϓ�)�"�n;88�I�w�        �k�~e/�G�W/poUZ9`:�DʲL2��N��d��=�������;�         �x/]ޏ���evUs�kV��h:�{"���=U�������{��q�o(         ��n���7��z�\������N��Л         ��aO�x%�z�۪&��l2Jt�����n����~)����Ǩ(
__         f�����_�������[�g1It��
܏c�{��J���L�s�z�^���         h��p_�Re���Ө�z�`V��f�'���Slo�����I�������,�e_        �V�����]��`����'w`:�DVy�{���(�$s����C�;         w5O���]���pq�N����U�����C���*�y�'�c��b�p���|         ��F�I|��Kq���%�u6�ga{;0=�{"����������az"w         ""b2��^����#"�j��1���'�	�{QI�0��        �'���/����|�d���U	܁�	��s\������(�ſ�        ���'����GDD������=�T��*�^/��sxx��         ����׾u1n-��j�1���^���w���(&�I��)         ��?��?)�r���6���'�	�{��O2�z��~L&�8q�Ĳ�        �1ٻՏ�_����ayZ�ߣw`z�DR��v;ɜ��7�`0��x�N��,˖}         z��A<�ݽ:Kӓ�&���k�;0�ֲ/���8���/�Ǳ�=��$s�e4���~�F�e_        �&UO�|-�~e��������O����	��⾽�[[[	n�=6�7�d2�[�nEY�˾
         5�(��[����e_宪�}VY�
Lo{�h��`�n��������z	nt������nǉ'"˲e_        �\�ًs/_�r4���c7���]��jz����S7n<RwΙ��v�Rh;�,"NDD7":����L��P����<ϓ�)�"��GY�1���ɓ���m        �U7�T�����+˾�=UU���'�	�h]��vz��œ	F�d��/lBeY&�����d�klp���$nݺ�N'��        ��n���{qT�}���	�[����}m��I�@��=���S�v�I���G�ߏ�,�ĉ��        ��ɤ��/ތ�.�GU-�63�q�l2JxRJՆ�<�b	:ܦ|M(U���],y�'�#p_/��8nݺ�����v���?         ������Q��Ѽ�̿�=��j2�DY����N���ܸq#���d�e_�IV5p�t:I����`0��7oFQ˾
        �F�?�׾u1�|��Z�����^��_�f���O2�G�G���{B�����$s^�"p�:��������	ݫ��\        ��t�/���W�u1n�i��������W_M2�'�'���{B��omm���N�9�� &5~qb5L&���z���/t        8&{����?9}�ոt����Q�7���.$��}(�����b�m/�M���{���EQ$��jx-t��z����������         `^�h��+W�.�:�UQc�{%p_e�ϟO2������~0��$���R�&�����k�;�x��`�� Z�V���h��bw        �)��Q\��ǥGq�����|�U���V�ބ�Ν;�l֯����W����}ϙ��5�&��~?�V�d2��(�l���ى�����ڊ���h�Z�eْo	        �xUQG�+�qX�V���E����L^U56�O�Ϋ���n�����ӧk�z�{���+���O���fl*�{BeY&��2p��<ɜעg6�p8������e��     �������^���
 ��O&1W1�4x5��j���&��F�uTUU|�ߌ}�CI�������'���_~9�<6��=�T���v�96��^UUQ5�st       "�Q�"  xM5�����W�׾��d����n���A���aܼy3�L6Kk�h�U����v���        ��j��}�=��cqtt�l�ٳg���������f�9�	����2p��4�'p        ��5���z^VM"�*�mHm8ƣ�>�t�������?��x�ᇓΥ��	�
���v�9�N'ɜ�(��         �PUE���޾>>���GU�}3�ٳg�/��/�W�Wckk+�l�K���*npO��z�$s         ��TM&3?'����w����׿�|n�ݎ�}�c����K��KBw�I���*�y�'������         �S5������9,�g?��c������?���ԧ>��ۿ?��?��������^��d�T܋�H2         XO�lpo	���s�=_����~���ӧO�G>���G>�����(�"F��m�?q�įd���Z���	59p��         6�\�'��I�S��T��O�T�y����<_�Y��,�n.�`ޞw$������ػ������s�oݪ��~���8��q�$L�	�a� �jY��h5Lf��V��,�#�$`�A$+%Z+��lL2�LL�`X�y���q'�;v����]��ު{�9��q�~��Suν���ZJW��;���e��_����         L�<���I>ڃ%�W_}5z衲g0�����*�*�E��         �d���L�>�>��OƩS�ʞ���h�op��         L�<����x��ײ,�x .]�T�f���@[[[�����)2p�t:�����9         �Lnp�-�.]����ߋ4��?w��{��,��h�_�[�Vk^377W�9�ᰐs         �ɴ��=���>����Ї>T��p��������Z-��fk"��n!��B�         &S�e�~O-�O�G}4>��=�"p/X�{DD��.�N���3�,�����          +�~��d�=�~{����hd;�&�.�{���7��h4�>g8��         0��,��{j�ܧŧ?�������H���� �C�^�*�E��1
9         �\�w7�O�G}4>�����J�S�b��U)p�v�,�         ���~��}�<�������O�=�)%p/���V!��         ��,o�=�|���VVV��`<���1˞Ô��J7�����$|�         "�l�oI2���J�4����,~��>{챲�0E�+*po�Z�>������         @D�m?p�e�=XB�����[��[�˿��q������IL�F��M�np�t:,������         L�<K���$w���x��g�����;�ɟ����^�W�,&���`U
܋��}8r         0���'yI��[ߙlgΜ����я~4����������,{B�^�*�sss,���         L�<Ϸ��$��&�h4��'O�ɓ'#I���;���;�#�?Ǐ��F��,{*#p/���V!��w:���        ��,o��w^��y�9s&Μ9�?�����tb~~>�$ٷM����q������J7��        ��d�^^˷�3��4����������&I���j����Z��MQ�{����sss,�         y�m���lk�� �L�^�*����vX19         �\y���}�GK�i&p/��V1�mTD���t
X"p         "b�7�܁��lop�����         L�,o������{��t����\K"�A!�          �+��m����N�V��Vk�gt:��D��B�         &W���z}�si00[�+*p/��n�[�7�         ��k���>�{��1p�����         L�<˶��Z6ڣ%�4������j���N���3�4��ȿ`         `��w`�	�V�ܛ�f���]���>         �|Y�n��w`'�+*p����sss����         L������l4E��/�W�l6w��V���w         �5�6opO��=ZL3�������f�I����E�E�H         L�l�{�܁��"�Z����;~����7D�        ������_�d[��k~�Y&p������T�{�W��/�         `�e��knovH�.\�P�9��zk)��^E}.         �d����ؙF��ѥK�
9�-oyK<��c;~o��\         �ɖm#Z�e�{����}����}��w{Ή�}��/�El�q���	����s�
9��o��ޗ$I��mo+dCQ�         0������Z���K�����\([=je/�F���w9�ĉ��t����o�=���
�P��         L�<��kk�܁���3g�rN�ٌw��]�~�����4M���/�,         `�eY����	܁��g���V1?Z���Ƿ��Z����y�ٳgc4r         0��<�4���ֲb:J`����x<�o~󛅜�����q���~�������y��O>Y�9         �tH��8��
܁���ӧOrN�V���韾��~�(��}         ���n��ts�� �J�G������������������ﾻ�g�i�N�*�,         `:d���^W�����}�<���q���B�J�$~�~!�����cǎ�������no_[[+�<         `�e��k�܁���<��_�Ba�;v,~�W5Z�֛�lii)~�����v=��c��         L�<���=�;#p�C�>�h�������߈cǎ]�؉'�7�7����=g4�ɓ';         �Yz��=��H�t� ӨQ��i���O�3�<o}�[;�ĉ�}(�z�h��q�=�D�$�����>���
=         �|��nov��{�3��L�g���������{�-<n��x�G
?         �|7�gw`��{�/��/����eϸa�O��o|�e�          *(ˮ�׳�}XL+��������=��ɟ�I�         ���ƣ뾦����9��>���>/��r�3��_�j�>}��         @E�Yz�����}XL+��>�F�|���4��c�X�3         �
������9��>y�����+{�U=���q��ٲg          �g�뾦�
�-��3    IDAT���|�#q�ҥ�g�ɷ���x衇ʞ         T\���}M}<؇%����������Ȳ��)��x��b<��wT         �-����z�w`�����������=#""�4����߉_|��)         ��n���܁]���S��T|�S�*uC������կ~��         �����k� O��]��w�������Gy��g�y����/��/Jy>         0���ځ{#��`Z	�K�eY|���������4M����ӟ���>         �|yz���.pv�Q��Y��O|".^�?�s?�nwO�u���x������{�         `:e��^����
x��G�W~�W�駟޳g|�_�_��_�         ;�������`�� �����K/ů�گ�����������馛
9��^�?��?��'Or         0���ځ{#s�;�;�
ɲ,N�<_���G�G�'~�'�����9�N���~����c�E�e{�         �5�ht�?������V�
��ڊGy$y䑸뮻���~w�w�}q�ĉ��zW|ϥK�⩧����z*���/�+���ϫ�K�$eO         ����׾��>Zߧ%���Wܳ�>�>�����z�X\\�D������������'         `o�G�����xc�� �J�>a666bcc#^|�Ų�L57�        ��Yd�8j�+$�y���<���� U$p        �+��[W�xc���������V�W         �䪁�xc�� �H�W p        �+KG�W�x]�@�W p        �+�ǣ+~����y	0�T�pI�D�$e�         �ʹ����>/�����^��=         *g�u��c�;�{w��F�Q�         ��|k���%y��Z	k�i#p���        ��5c���5F���Y	k�i#p��h6�eO         �����7}���\�`	��*�$�z�^�         ���ƛ��h��%�4��5��         �^�Q��f���76��C���j�ʞ          �q����e�o�xs��@1�p�F#�$){         T�M碑"��oq����_!z�	�;\G��.{         ��ըő�H�q�ӿ�;�s%����������_��         �����%IDD���?��R�$`
	ܙ);	���z4�=X         ��#��wc�I�E��Ra��v���E��L�I���t
^         ���B'��˿o�_�;��Q˶
yF��fw�uw��V+j5]         �Mwݼ��߷�"��X\~��g����3c�,��{��        �,��6��b�ko���~&��3�!pg��&po�ۑ$I�k         �����?^�}�p�z0��̔��I�D�۽�        `J,t�q��޾<ku��/��M��L�M���t�V��        ��p�K�$����hT�R�������%sss,        �j;|�7-�_3�:�wf�x<���V+��fk         ��jI��o?��ϼ������I��Lɲ,�<��9nq        `��ul1z�������>�&�;3��[���zt���         @��:͸���}����}&P=wfN�{DD�ۍF�Q�Y         PI��Z-��g���w@���F�����
;         ���c���k��s�,�����ܙAE��z]�        �TX���[����1g�<��;3���="��nG��*�L         �O�z-���7E-IJy�s��Ky.P=wfN����i�g�z���녞	         �!I"��֣�m5J���9�;��;3iss���$����HJ��5         ة�.ő�R7<uv����!pg&mmm~f�V������        ��r���x�͋�nH�<���j����3��"p��h6�"w         &����Gw.{F|����e� *B��L�F1����V��^oO�        �"��]w��$){J��' "pgfmnn����v;�����|         ة�n3�}��Q���GD|��W˞ T����5���N��nwO�         ��k7�=��f�	ikO��R��B���	J0#˲=}F�ۍN����         ��k7�'n�V�^��˞x�b����@�ܙi{}�{D���\�����s         �j��x�[�]��="��^-{P1wf�`0ؗ�t:���z��,         �^�:���G�,���se� *�Q� (�p8�4M�^��i����j���y�ǩ         ���-��;�r4j���)o��g^��fZ��b����������f��$��         �˝7-�;ﺩ�q{D�_}���' $pg��g��h4����rk<         ���D����q�퇣����F�O�Z����̼�x������z��v����        `�uZ�x�[⎣eO��ϝz)FiV���e�*X[[���<I���z�h4bccc_�        ��9�؍w�u4��j����ċe� *J������(���?��nG�ш���H�tߟ        �dK������o9IR����ڳ��.����ߢ�h}}��g���8p����"        �d�k7�=��{�OF��/~��	@����N�ߏ���h4��k�$I�z�h�Z���Y���        ��K��ێ,��n;�ڄ������x��Ųg &p�ﱾ�,uC�ٌ���1K�        @��w��}w��^��)�����"��^T���G�ߏ����nq]�$177w�6�4MK�        @�jI�[n^�{��Z29���������o�+{Pqw�y����j:t��)�h4bqq1��a��}�        �L:�4�޺�v��);����g#���!p�`0���f�����-�N'��v���Bw        �q�׎�-��|��)��V�O���>�;\���J=z4�
��$I���F�Ӊ~����eO        `��:͸���8��+{ʮ�y�G����nW�F��
F�Q�������I�D�׋N���P�        0E�͸��bܲ4��uW�������e� &���bee%:�N�����\Q�^�^��n7677c8F���         &��|;�:�7-Ε=�P�Q��wʞL�;\E�籲��*{�5�j��v�o��4-{         �QK"�-����|�Y��=�����xuuX�`����A��v�eO�!�v;��v�����܌��-��        TH�D���^_�E�Y/{Ҟ��K��<_�`���:�����jE�>9��h4��hD���        T�|��������kO��fy��z*�L�l����]ʲ,.]�G�){ʎ������h4��x��(�4-{        ��j�kqh��:qd��v��I�����g��s�e� &��n���f������|�Sv,I�h�Z�j�"""���F��w�;        ��5�X����ע��v$I٫������_8S�`B	������!�tW
��4��+˲˿�<�<�cb        �ٕ$�F-��zt���k�ݯN3t[�iI2#"և�����dd���_M��y/^��G�F�^/{N�$�F���տ,����     �v���[�m�ze�  �dIѨ�"�ڹ�,���������)���6�i.\��G�F2�?;���y?w      fK���m�  �����?_�΅�g η�6�F��x�[�        ��|�;�?�\�3�) p�����Z�         (�s���?u*2���������F�3         �4׷������L˞L	�;�����        ����9���O���˞L�;����r����g         ��������x��z�S�)#p���        ��,���x��岧 S�Q� �y�ǥK�"˲���/{         ��Q���S�g.�=�Rw(���J�yeO        �B���?��'�3�ʞL1�;luu5��q,--�=         
�6������V˞L9�;�~�Y�šC�"I���         ����<�������~�S�P+{ L��p�Ν��hT�         ؑo�����_�����q�?>������=         n����K������� 3D�{,��x�b�z�X\\�$Iʞ         W�fy|�����gʞ� �;쓍����܌C�E��,{         ���˃��O��o��Z�`F	�a���8w�\8p ʞ         ���7�Ň>�T��eOf��J����� �����        @�����g���Wʞ p���F�8�|���Ł�V��=	        ��7�8��7cyc��) !p�R�y���caa!ʞ        �x�� >�oŗ��j�S �@���y���F�ߏ�������$Iʞ        �������~7����b�fe�x�;T�x<������؈D��){         S`�����g�O>��7˞pUw���h.\�F��^/z���        ض,���7��������A�s �K�6�cee%��֢�����\4��        pm�Q�>�r<����ً��� �0�,L�,�bmm-��֢�n���\t:���jeO        �Bέ�'�����X�ʞ�mw�0������I�D�Ӊn��N'�$){         %gy����#���x�ً��yٓ vL�*��1""��nG�Ӊv��f��u         �,��/���y.������Vٓ 
!p�)�����Z-Z���_�f3j�Z�        ؍��(������3�+�\�����>w�BY��p8��px�c�z=��~�������w        �
���O�]�'_X��^X�o��Y��=`O	�aF�ii�^�����j��.I���      ���usD�ʞ ��X�o�++�x�� �;�Ͼ�Ͻ�����f�)#p"�[߳,+{      T�}>^��/{  S`csy1J�����9���(V[�6�++�l�e���;       �����eO   ��T+{            D�          ��;           � p          ��           T��          �J�          P	w           *A�          @%�          ��;           � p          ��           T��          �J�          P	w           *A�          @%�          ��;           � p          ��           T��          �J�          P	w           *A�          @%�          ��;           � p          ��           T��          �J�          P	w           *A�          @%�          ��;           � p          ��           T��          �J�          P	w           *A�          @%�          ��;           � p          ��           T��          �J�          P	w           *A�          @%�          ��;           � p          ��           T��          �J�          P	w           *�Q� �e�Z�f�j�h�k�i�#I��g 0V���Ҳg      ����<�<���,���{ &���H�$ql�o�i!nY���t��N�o�|���z�Z�г ����~1�rf��      ���<�,�"M�H�4�,��x��(��q���� �L�9�4��y(��`�yd.n?ԉ^�^�,        ���$I����ׯ�o�y[[[1�bkk+677#˲}^	���a�{�xϽ7ǻ�z8�~|!�7˞        �u$I�v;���句i��0677� %��6�|�?r����{�=7�"I�^        �n�����z���""bss3�A�;�>��u�w[���y[��o�)�y.j�v        �����o���</{����U�����u[���K�n�ʞ        �>K�$:�Nt:�X\\�~��~?F�Q�� ����G-I⟼�x��=W�         *�V����|������V����p8,{���CD4����sW�����82�,{         �j�����1�bmm-�Aٓ �����VK���w����7h�=        �	�l6�СC1�cuuU�P �;3�}o�%���;nYl�=        �	�h4�СC������1�ʞ0��̜;o:?��N�;�8P�         �H�Պ�G�F�ߏ���Ȳ��I�5��O��񍍍�ݞs�ԩ�s�΍��4�Z��33�Z|�����[�Y��=        �)�$I�z�����������({p_���N=������	ܙ	��y$~��}[ܺ�.{
         3 I�8x�`t:�XYY����� 7B��T�ג�W�����?p[�kI�s         �1�N'Z�V������ܙZ�^��S�(W�         fX�V��F�ݎ���Ȳ��I �%pg*���n��忹':�Z�S          ""��n�Z��x�blmm�=���L�Z-����x�mQK���         ����8r�H,//G��/{@�ܙ�N3�����n[({
   �?{�#�}��wN]�t�m.�s�ep��=�cǗ� ��$�1!�Y��c%҂�V�� /@$�Y=R����U^��P���R$ �DH�^;���%3��g�R�]g_8N|�t���_u��F�t����]�/��+      .�(�ػwot:�8w�\�u�;��Pp������o�k���         Wd~~>��v<���J� �W� ��������?�Tn        `�TU+++�j�rG
�L�������{zތ         ����tbyyY� ܙ`���`����s]?�        �l�v�&w�PpgB�����?}STmG        �fh�Z����v;w�l���8o�������DtZE�(         �T�Պ��e�܁����D��������[��8�         4��;0ͼ���������*����Վ�ݍ�3e{&���⟢�(��[Q���� ���[D,_�     �1���u]�ŋ�����܌�`[[[���kkk����~?wԩ�n�c߾}q��ɨ�:w��Qpg",�f�����X��m����h��E{f.ZU/�N��B;  y-�cys6w      &���V������z�;w.Ν;gϞ�����ѦJ�ۍ}�����?��Lw�^�U����qh��;ʔ+�=;�ޞh�.Dkf.���        h�V����1??���?�������'O��s��)^Yعu�    IDATUU���gΜ�`$�S{��n���rǘJe��No):s{��[����        �lff&VVVbee%������؈�'O�����f477�~?VWWsG:mU����X�����/$��Չ����..G�Z�        c333q���8z�h�x���㩧���{.�A�x��gϞ��܌~��;
�P)�3�����_��c*E��}�]X���RD�#        �,�X^^����x�b|��ߍ��z*^x����(�ػwo<��sQ�u�8�+KKKq�ȑX\\���bff&���G�aϞ='>��ύ�1�2
n���M�i)ZS���̞C1��`�N�8        @Ct:����k��k���g���?�>��b�.���طo_�:u*w�bUU�M7�7�|s��-o����:���rǊ���[>��ϝ˝��Rpg,�ҽo��{gr�h��SE��P�,�(��q        �[ZZ�[n�%VWW����'�|R�}���^�������%u�ݸ뮻�=�yO�r�-�j�rGb�(�3v~����_n\�����L�._݅�a;>        0:�^/N�8ǎStߥ�����؈����Q�VVV�C�P�}�����r�aB)�3V�N������uREيj���        �ꥢ�5�\=�P�:u*w��S�e�ٳ�׎�q�������=�yO������X���8��:�c4H3{�����h��        �c~~>��x��������ܑ&JUU���buu5w�X�Պ{�7>�DUU���
[�[��oܟ;Fc��*�^�م�Q         .���ñ�������'����sG�KKK����� w������W~�W��ѣ���0
VY����7GY��4�����]�6���;
        �e���x�[�+++�����_��,cqq1Μ9�;
S�(���>?��?�*2�9U����X\�6w��W��1w��h��rG        ض}��Ż�����7��>�l�8���Ņ��ŋ��0���_��_�;�3w�� f����:w��מ]��koVn        &Z�Ӊ[o�5n��(K5��)�"����������'?����y�'����X����n�,���ND���        ��UW]w�ygt�zQ�333UU�A��ݻ7~�w~'n����Q�
�d�w��{�v0w�	V���5�;���·3        �,{��w��177�;��[XX�����z��O~2�����Q��du��_U�1ܑ����ǣ�w4w        ����z�w�#��ݛ;�X�v����\�ۍO|�q�ر�Q�"��d�w���ߴ�;�d*��?r<:s�r'        �n�w�qG,//�2�lq'�_��_�o�1w���;��/�8]�۷�(b��r;        0]ʲ�[o��&�7��v����AC�s�=�c?�c�c0���ɢ�n�O�|0w�	�������        ��i�Zq�m����R�(c�wR8v�X|����)��N?��kbq��;���\ks;        0���v�~��ܗPUU���y�\Y������trGaJ)���=��a�t�cf��        @�Ӊ�n�-��n�(cinn.w&�=��Ǐ��)�%:�����ď,��1QZ�\�|S�         c���x���_��ע���q�J�׋�g���Z\\��|�##y�����c�=�<�L���#y̗۳g��GG��\��;#��ۯ�a��v��!���         /��������G�e��e�������;
�~꧆� gϞ�������|�+��c��`0�c]NQ�V����Rpg�Ze�:�?w���[9e���         ��뮻.Ξ=�=�\�(cennN��m��z�?��C�}������Cy�C�����n<s�V���[���J�         c�n�3g�D���el���DY�Y7d3Y��ޡlo��W����g�̙3�g�Le� L�w�p w��Qe��.w        ����v����c�������(�"����%����>>��O+��-
�L�U�m���11�嫢�T�c         L����:��ݛ;�X�*4��7��J:����_�B�u�t.ͧ����z�JTG�J��NT{�        0QN�8e�������(��1� �y�{�����<�@ҙL���oZ�ab��;Q��        ؎���8z�h�ceff&w&��ߞl�7����?��d�>���m?�_�D�j�����1         &ұc�l-���rG`�>|8���,1������~6�A�yL'wFbei6/yؕ����l�        0�z�^:t(w��a�;�s��7'����3�<�l�I��������#L���J�         �뮳�����v�Z��1cǏO2��ŋ��$��tSpg$N\�7w��О]����r         �1??����clt���cG�M2������ٳIf1����Y�a"t�sG         h�Ç�06�y#G�I2�����w��Uq�^[�/���W        �p���(K5Ɉ�N��;c������b�Y���7����ݏZ�Nk�Gm�݋��CCH4�ڳ�Q��J         �N�����c,(�s)sssI�>}:Ξ=�d(�3to:��W�����]qz߭����l�W@        ��0ʲ�V��;c���%����&���h�kW�}�Fu0�3/�rnPv�\Lk촫��         �4�������V�������Y[[K2g��8r�Ȯ��'O��V��_M�i�1����FD'"
�ݡ=�۾gu����=������Sk&ͫ�         xQUU���buU��w^O��I2gss3ɜQ��7�y[��V�; �w`qf[���^��ma����l^e���}�         �������B�m'20����ߜ����ޛ��ԑ�΋��"w        �ƙ�o���+��L
w���cnf{ok�Q����[��܋V���         ���_�jm�����;C�w~���J����jͦ�3�ʖW�        ����{lMTE� WD����3Wm���ݥW�}К�_.
ߊ         �PU��5QY����C���n���(c�����m�ۛ1�
�8         E���a,(��³C՛��/��Ũ_��|0w         �C����܁I����괷��A�����ZݨS        `�(u�PQ�# \�gm���������:-�n��         ���Lw��]n��f���#"�L�8         0�܁I���P����.���������          �N��1R�V������Έ�           ������j��������=�4          ��)�366/��="�.�         �����K~nPtF�          �A�����w�         ���o���.mp         ��Spgl�Q�}`�;          4��;cc�ݻ��lp         ��Spg<eޠ�>Pp         ��Spg,l�f�~���EkdY          �<�[e���6�         @�)�3�Z�o|Ai�;          4��;caо�wG          Ok����z�{���          �Qpg,l�f���u�Q           w���6�
G          �Nk��0h���(ʨG          �D���p��ED�I           w��#b����u��;          4��;�ZUDq��X��;          4��;�Z���Q
�          �d
�d7hUWt]]*�         @�)��ݠ�^�u6�         @�)��ݠ5se*�         @�)���Vye�A�         @�i�ݠ�^�u��          �h
�d7h]Y�=�         ����nК����         ����n���;          4��;��+��
�          �h
�d7h]Y�}��          ���NVuъ�
��u�         @�i�Օno���         ����jP^y�}��          ���NV[e��/.��          d��NVu��7�ׅ�
          M�1LV�mlpDk�I          ����jPv���R�          �L����mlp�w          h2w�l���         @�i�ՠ�^��
�          �h�d���+          4��0Ym��^1	          ���;Y��_\��          �N���lp          ^��NV�*��+          4��0��E+�h]�
�          �h�d������
          ��1L6u����bHI          �q��N6�b{܋�5�$          �8Pp'�A���{��         @S)���v�u��         @Si�M���{(�         @ci�͠ho��:�!$          Ɓ�;���
�6�         @ci�͠�l�&w          h,ma���wG          K[�l�r�˦�"w           �n�+�!�        �ʲ�cǎ�7�7�pC:t(bqq1""Ν;/��B<��S���ǃ>���wb0dNͧ�N6[�N
�6�         ;����~���{�\�^���7���q��wGDĩS��o��o�����Qb�>
�dS��c�;         �=�����/����EY��������Ї>�w�G�O�N�Pp'�����{(�         W��j�}���Ї���&�Y�e�}��q�]w��?��x��b0$�(��Q]n��ա�         \���J�گ�Z�x�C�_UU����\�~����|�6wHD[�l�^_�÷         ��M7����g�Vn��o�9~��~/��?Lma�(ʨ�ֶo��         x#w�yg|򓟌����=�޽{�S��T�r�-#{Lh*ma��������H�         h�;�#~�7~#��������������F���$
�dQ�;+�G����         @���o��}�c�j��v�����?W]uU�0����w          ��{���?��*w�����������rG����Nu��ٍ�#         �PY��������;�:t(~�~)w�H��d1(w��]�         x�~��q�-����z׻����&��0Y���
�#         |���J����c\��������b�0Q��ɢ���:��I         �I�я~4�������p�0Q��b�ܣl�         L�n�!���w�qY�����ѣ�c��Pp'�A�����         @D���ߟ;�)�2~�g~&w�
�dQ�;��^8�         0�?��rK�W�����СC�c�D�&���kw         �z��{o���j�����0���b���Xi�          eaa!~�G4�����������������p���a���������7:�Nҙ�D
�����         ����~wҢ��ӧ�7�7�/��/ccc#����K_�R|������d����w�qG�y�T
�dQ+�         ;p�]w%�u����ԧ>���w^�Gy$~�w7�A��K��J��,���
�         0�����ĉ�����q|��߾�����ǟ�ٟ%{�;�#��yh"w����B�         ������(�4���<����������i�:u*�c�z�����̂�Rp'���mp        ��u�M7%����>��e���؈/~��7��H��,��ٍ�#         ��o}k�9�<�L�˿��_��/9.\���O�8�d4��0Y�t�{m�;         L����8t�P�Y_��h{�K��~|�+_I���_}�>$\��;Y����        `*]{��f��?��������$�]UU8p �,h"w�����        �4JUp����O>���{��ccc#I�k��&�h"ma2("vXp�mp        ��t���$s���o�辭��x�G�dH�o�&Rpg��N��GD(�        �4ڷo_�9�>���}�ǒdH�o�&Rpg��.�ud        `�*�?��;��?��?�dPp�K�f���         ��,,,$�s�ԩ�{���$�́&Rpg��r��	s          �cff&ɜӧO���3g�$���v�́&Rpg��b���pd        `u:�$s666���r����D��`%�:��I         �IQUU�9���;����'�`�;\��;�W�|�{](�        ��)�2���~���`W��`�;\��;#WGkw+�        ����*�Kr���vu���Ʈ3D(��Qpg��b�n7�         ���$sv[p�x��6��D�.M[��;��^��         Sgvv6ɜ��뺎~����n7�Fzh"wF�l��^O�         0uƥ������EQD����h"wF���wG         �OUUI欯��zF��333I�@�h3ru��cW��         S�i�#��R���l��nw         �6�^/�w
�\���l�;         L�������{��M2�F��������Vp        �i3;;�d�8�mp�ק������7��M����         $���C������.�V        �i���C������(Y         �6UU%������
�0\�\���z�0         0Rmp_]]���~�� ��;\��;#W��l�;         L�^��d��0�����h�rB�$         0��J2'E��w.wF�����Pp        �i2;;�d���ڮg�����v�́�Qpg�lp         �#U�}uuu�3R�mp�ק����e{wv�         �,�
���뻞a�;��0#W���Յ�         0MR��NRp�����a�;\��;#W��]NPp        �iQ�e�m�1��IA�^��;#V�n굂;         L���#"��֒�Qp��Rpg��"��K1         �UU%�����d��;��0#U���H�         �M����v�́�Qpg��lp�"�         `�*����&�c�;��;������$         L�T�T�tw�v� I�|�ӟ����$�r������җ��;�P�I^Sa�;         L�T����$s��~�9
���Ƣ�^�i6r�߿?ɜ����sG�4���        `Z�*����&�c�;W�f9\�$�B�         �E�����z�9��������9�n7AhwF�h�zD�          0R���֒̉H�Ž��D���^%4��;#UG���6�        ����*ɜq+�G���G����lp�B�         �ES7�GD���$�M���H�E�#��         �B����;����^'�         L�T����$s""��~�9
��Z
�T]�v=�H�         �UU%�����dN��;��0#U��g$�         L�q�ྱ*X�<    IDAT��d��;���;��`�{��K�         �d��zI欭�%���ä��H�	���         0=��J2g��n7�hwF�.��w         ����I�c��wx-wF*I�=�        `Z�(�����	Ҽ�wwF+A��nb���s'         ���j�����z���F��~8/�������E��         �VUU�9���I�$�6xwx-wF����uՃ��         )��nF���%�����d�Klp��Qpg�Rܛh�y1w        �FRp�l���I欭�%��wmcF�Nq��mpl�y�         ^iss3wv���$sR�_����u��$s�I����bH��epq#��*A        ��R��T�WWW��y��0<
�T]����,�G]�����)         g}]7k��z�$s��֒�y��;��;#���E������a         D\�p!wv���$sƵ���v�́&Qpg�R�js��         ����#����I���o�;��1#�b�{��ྐྵz.w        ��9wN7k��*����&��wwF��V�ck���~ڷ@        �fq��1؅����Y[K��Sp��Qpg��"���[��U����         �ԩS�#�K�6����'��w��6�O��o��d�         ����O��.�*����C����l_�#��1��q!�6�        �n��}�`\��~?���wx-wF*E��(�[p��X?��         ����O') �W�����z�9/�����9
��Z
�T���5y�{DD���\L��        `�<��e�M0��#"666v=�,��t:	�@s(�3Z	6�7_��?�;        ��:y�d�={6w��*ɜ���$s^.E�="���&�M�m�H�Ek�C�fop���8��\L�        `�<�裹#�H��K2g}}=ɜ�KUp���I2�B����lp������X;���S         L��'O��ӧs� �T���֒�y9wwF*E�=����N��~�        ؎o}�[�#�����g����	Ҽ��;��;#TD�rz�� c��G�l�        0�x�8{�l�$�n���n�z���z�u����;��;#�f{{D�h�$l�c��wr�         {�����#��AB)��GD���%��j���+��+MOS��Rܧi�{D�ƙg��3�c         �������Flmm�BB�^p���C��������3�Ġ?��         ��'��ӧO�AbUU%����E��I��=ٜ	Rom����Qom�        0VN�<?�p�A��K2g}}=ɜWKUp�v�I�@SL_S�l�D���N2f�l����3�DĔ~         ^�������=�i-�5���l�96��dQpgd����omm����7�E�*�Ĺx�L�>�h(�        Ӯ��ǿ���d��*ɜ���$s^���'�������蔯<n[[[q�̙m������q�9%w        `������W�:��2�!�����$s^�wwF�~�q��܌^xa������        L������W�����$U�}mm-ɜWKUp�v�I�@S�s`��,�����*��鎈K�u]����^�        h���5�ۧȴ�mp�WRpgd^��}mm-�������/��^.n����Q�:��         �����k_�ڎ�2���J2G�&��όN��b���j\�x1�m�d�k���\;����Z?�;
        �P<���O��O��S���%�3�s��á�����^�u�;w.�Alnnnk�����a�ُ�|0.�?�;
        @2u]�C=��o����ovv6ɜamp���I�(��+�s`z^Vpi{{ċO�N��6���z���p�,�ٕk�(}{        �k}}=����=N�>�;
�TU�d��0Y4`��ӟ����KE�mJ��6�>/�����3�7w        �m��w�=���e4I��I�Z��{��M2�B��z��^�u�<y���[t��~Y��~�ꡘ�s(f����        ��ϟ�|���!��ꫣ�A��'�LV�ގT�q���jS=4��+�S�q���W��nsss���j��3���NE�|u�,_;        `mnn��?�=�X��q�c�X9rdG�=��CH��R���֒�y5�a8��:���:�y�W||kkk�sꔱo�u1V�}46N?�������;        @DD�xꩧ�[��V����q3�6��{�}ff&�h
wF�(��g�}���np/l!ߑ��Z\x���}.��WE{v1w$  ����;����?����]�	IH��Bò$�a��Gb�7�4uR�iZ��'i�ę$�x2�q�:�t&M�ɴqj���9�IǍ-�!�2 s���������66Ǯ���~���|�0ia�~�-t�����        �Q������u�����J��A%uޏ�;`�Lx�!ǎ��狀�]��%�hpD�y��Z)��i��            �����رc��;U�C��X,&�hT�4�F%��ai�!�\��;,����JH,����pO�*���8 ����-�Oa�8�|I             ����9rDN�<)��sd����nq:�i�1���H$�v��v�a|n �iVXb��b
_>���w��U�G�%x���w�T�+�&���"���(            �ۂ�������������+�c�I���i��x<���@� ����
d���>11�Z�;�M�HH��Y��;+�K<SJ�]P*n_!aw             I	�r��I���Q�� ��|>%u������G�����T��U�3Vr�װ��~�	9%�#���0��+��H��"qz��            �M�����А����v(��V����
�{<%u�l@��p8�d��V�ɵ���p�VJ$��H48"!1�nq�
ę�/N�_�yS�p�            �v�hT���dllLΝ;'CCCt��,�j�{0TR�JTnppw(��zeŊ2s�̤^��%��aI��Z�y�+�J��Y�sg/���t�3�/��'��s��;OW�.��#��[             ��b1���q	���7��ؘ� /��߯�N(RR�J��p�Ruuu��ܜ�S�X,逻��w��Ǣ��G.�q8��p"C�S�!b|�  0S��1�c         �����b1I$��.�����=p���UR'+�s%��H�B���*Y�x�TTTL����xүM��=�$$�������Y   r���Y�=          L���;܁�C����x���V�͛'ӦMK�V*wa�;              Y���)��Թ�zܑ���),,���2������r1CI��$�             �j���pXI�+�D"J�p�E�=���~������b)**��'.�K�nwJu�^���nq8���p              �,S�lp�#��e


���N�̙#EEE��I�             ����`PI�+Qp�x<J� ـ�{�(--�n�AfϞ�{�II)�N�             ����z��	�BJ�\I$QR�����g8��/7�x�����%-��$�             �j~�_I�p8��Ε��P��{�;w��������=J�R	�o              ��|>%u���*��w�]�3�a�|�����^�X,��&&              ��z�J��A%u���;���r���[o���jݣ(�H%��`�;              �L��p8��Εp�#��A\.��q�R^^�{���xүe�;              �MU�=
)�s%��� 9�a�-�ܒ��v���a�;              ٌ�;���g�%K��̙3u�a�X,���ɷ             ���x�޴��b1���P0ѕE"%u��"��f̘!�_��1L�H$Rx���               �<�F�W����p�@���N�����Ñ�k�S	�K��/              �e>�OI+����J�p�E���-Z$��0]<O��!�             @��z�J��A%u�FU����(�d�6���'����ǰD*�S��              2���WR'+�s5lp�#�nc����v�u�a�T6��             �Z>�OI�P(����p�#�nS�C���u�a��6���             �l��z�Ա"���$��]��;�.�6UYY)����ǰL*w��[              �U&mpQ����t���T0��H
�TMM��,�J�              d�\��������MUVV��R�܉�             ���^��:܁�D�ݦ�N��{K���^�0m              �����pXI�k�D"J�p�#�nCG��S�             �l�����ɴ��GI �p�!�Ƚ��D"�{              `^�WI�L���8ϥ{ @$��9��    ��s����x�����xTg(�X,&�����	        �҅���^	����R��ήw    @�(//���:�>}�TTTHEE����KiiiR'�E�Q������Q���aٳg�:t���        ��
��A%u���Z�mȑ��S	�;$��?    ��PVV&.���Fijj���Ҵ��n)))���������^|�E�        ��T�C���:�B�P��;l!�'����     ؞��o�QV�Z%�/Nj3;        @6�z�J��a%u���;�wd��p    �>EEE�v�Z��[�m!        �lprw�F"�G2�u��    �������o��k�l        ��߯�N0TR�Z�jp�m��qq:��~a��Y     0CKK�<��#RXX�{         ��z�J��a%u�%�(�C�8��;2O2[�    ���-6l��|�#�G        �5�á$��F%�)���Tmp�x<J� ���;l#�Hn5{�/    ��O�.O<�TWW�        ������0���B!�$��Z�a����    �����o|CJJJt�        �|>��:V�Ump'��G���l��x;     ̙3G�|�I),,�=
        @�Pp��J�$CU����(�d:d�I�y    @���J��7�!����G        �(���`PI�d��P��= �2;�    �����o��o�        L���UR'
)���Z�a�x<�Wp    ؓa�/|AfΜ�{        ���j�{8VR'��lp���W"��=     iY�f�,Y�D�         KU���@�E�����`����    ����jY�n��1         2w ��     d2�0�/��/��v�         ��
���a%u��D��!��G������$��     k�z���Р{        ���w �a��    ���#����1         �B��Ud 	��pGr�     ����.)))�=        @V�z�J�XpO$�FӮ��x�� #	p�m��    �i����{��=        @����J�Xp9��=]�a���R0���,�m��q�#     ���Ò���{�K�9sF:$CCC%�����B),,���
����=&        �ee�w�����������)�d2��<�    ���)w�q��1$�IOO�������#����|��!�ǂ�         R��w����ܹsJj���;l#�H�    �����ȴiӴ������o���?/���)�m"�Pv�        @%�߯�N&܁\G���Hv3;Ax    ����~��	����/�6        �|>��:܁�E���w    @�������-�����瞓`0��?        ���^��:�pXI�dE"%u��a#�ܓ��    �IV�X��Id
mݺU����J,��7        �Tmp�:��w@C�       ���p�ʕ+-�g�y��g	�       ��e���w$���������QR�dܑyX�    �h޼yRQQaiϡ�!����'��        ����Ur�n(R0Mj���C�      ---���я~$��Ö�        ����UR��;���     �ছn��ߖ-[d����        ����+�C��l�a�D"�W��     �Q[[+������b�ӟ�Բ~         :e��H$��w��;l$��;     z477[��7ސ�'OZ�        @U�p8��N*���C���p$���<    @�%K�X�+�H�/~���        ������	�J�BU����(�d2�6�    쬰�Pjkk-�w�^9v�e�         t���J�B!%uR�w@��8��y    @�n�AúK)����-�        `^�WI�p8��N*"���:��6�    �lѢE���F��u�V��        ؁��SR��@f#��p8��͞��     P��p�-���[oi�,        �w�w��    vUUU%��Ŗ���견        �]p�x<J� ���;l��;    ��,X`i��۷[�        �T�u���w@��8��    Vkjj��ױc�d``��~         v��z��	�J꤂�;�w     ��p8���hY�={�X�        �N�~��:�PHI�Tp�!�     p3gΔ��"�����Y�        �NTmp��J꤂�;�w�F"��=     ���di���^K�        ؅��SRG��H$��w��;2�á{    @�2�>66&'O���        ��dr�=�J<O�w��;     ��!��Ϸ�����9�        �,U�p8��N����Ӯ�v��0��"�� �H�>��    �9s�Z�������        ��D"��w�ǣ�����6�P    ��X��СC��        ��0�����%�+�hr�U���SR�T�a�C�     \�����~���        �]���."
��ԙ�.� $���<    ��C,�
��ԩS��2��땼�<�z������pH^^������_����LLL��H4���qI$266&�Ν�v\m���˓��),,��+.��K�^�W�N���MLL\����$
I �P($�`�����0�2e��������)^��������_C��%�����crÐ��|����|m��Ͽ��F�Q�D"
�d||\��	L     �Uw��{	�jp     ����),,��ߡC������z���Ȓ^�HD���,�e��'���2}�t�������:u�Jaa�'�T%���������Ȉ�:uJN�8!200 gϞ�l;����3fHUU�TUUIuu����JAA���.�pXehhHeppP�9"G��cǯ��    IDAT�I,S���^�̞=����¯��)((Pr*f<�������3g�ȩS��ȑ#r��aQ�_���_���h�_'Ð��j�3g�TVVʴiӤ��\�M�&%%%�<(�B4���Q9{������?~\�;&ǎ���Q��py��	��9�}    ���7L܁�G����M|V�    ̷`�K�͟?_^|�Ŕ�&��?̦ciii�G}Ԓ^{��o}�[��Jה)Sd�ܹRWW'���2g�K I��햒�)))��k"���8qB���/��퓾�>9q℅S�Q^^.7�p�466JSS�L�:���^�W�������611!G��={��Ν;孷�ʚ�N�S,Xp�}]WWgz��0�:u��^GGG���Wv��-;w�w�y��yT[�h�|�_����ݻ婧�J��*++e�ҥ�p�B�?����p��RZZ*������ӧO˾}����W�z�-9r�e�e��-ӦM�����L���eʔ)���%??���}��%.����&��׾&����=FV���>'�Ї��>|��|�K_��;�TTT�~�m��������/�(/����޹d͚5�a�m�_{�5�я~��?  �2U�u�ZH�P��;lCŶ!     Till�=�5���˂dǎ�G>`֬Y���"���2{�l��(��xd֬Y2k�,���?,""��òo�>ٵk�tuue͖w��/˖-��+WJCC���ݹ\.������Z�뮻dbbBzzz�����twwg���뮻NV�Z%���{����P������YDD������k200�y:{Ie۹�瓛o�YV�\)uuu&N����2)++�+V��ȉ'd��Ͳi�&9x�����6m�ůA�gϖٳgKYY�� KmܸQ[�}֬Y2cƌ�{�*�,[�Lk��Ǐˌ3��noo'�n���V��7nܨ�?  �2Uw�1"���:ܑ���6���n�{i    �,�p8���A�Iimm%��(,,�;�CV�Z%���ǱDqq����Jkk�<��ò�~y��ץ��C떠�*((���On��v�x<��I��咥K��ҥKeddD~����/�K��'�n�����u�]�{������}��'��{��ݻW^|�Eٳg��ladd䚯����f�����%??߂�Ԫ���{�W��^y���׿������`I��^�����ҥK����0; �O���PV[[[ʧ_!5mmmZ����k��O~RK着*�={�:tHK�\PZZ����@ �ϯ  ؘ����k�lp� ��H:�    ��jjjl�A�Jn��&�����2�_ee��}�ݲjժ�	E���pH}}�����C=$���'���/�ĉ�G�&��-w�}��Y�F�~��q&���H֭['��v�������N���>���V>��Oʂt�2i�C������I�o�.����.G��=�VcccW�3��!+W��6Hqq��S����V}�Q��'>!/���m?�&��r�M7�$�Їd���t:u��J,�͛7��ի��_�bw���Kmm�������ꫯ�]w�%%%%Zfhoo'�n���v�'Dm޼Y&&&��  WG��]ܑ��#㐃    �-���`�����=
r���x@>��{��#�W��[o�U6n�(�?���:uJ�X�UVV&�?��̝;W�(��g>�Y�|�|�{ߓ�g��ID·�?�Ȇ��ʞ��/�����s�����]f2<<|���z���}N�-[f�D�())��|�3��X~������u�4ir�m���7ߜ1;�lܸQ[����R�̙#���Z�g;�߯6o�,�hT6o�,w�y���/_.?���r�g����j���٩�?  �:U�p8���dD"%ury� "b�      �n���t������# -Y�D�}�Y���	�_�aC��ׯ�ۭ{�K,[�L�}�٬
�������g������E����'���z(���8�Ny��������R�Ν����3�<�=,h���Zy��eݺuZ��NFAA�<������r�=�n��w�^��?�����֦���M�DDoyڴiR__��6+--���:m����޽[[  pmlpW�^c. �     ��aHCC��1R���B��q:���C�W��U)++�=N�p�ݲv�Z��w�#s���=����Z�J>��ϋ���=�������'����Fm3�|>��׿.K�,�6�U�����_������7����˷��-����4��Ðx@�x�	����ǹ&��)k׮����r�����-0Y�x\�l٢�����3�a�LP^^.��������ʞ={DDd߾}r��m����k����ڴ~�nٲE&&&��  �F��]ܑ���6�?⍋U     ����HAA��1RRXXh����~�G���G?�Qݣd���jy��e���Z�X�b���_��Fn\"��˓'�xB���:�{{�^��׿�uS��.\(�?�x�=|����o}+gZ�d�<��S����{�+�6m�<��S�~�ze7ρ\��ѡ�wii�̛7O[�le��q,����/lsס��=�~�����t�   ��jG6�=��:@�ʍ��lY     �ASS��&E�1��~n�[��կ��ŋu����n�<��#�a�-���ϟ/�W�3��|>�|�_�4��p8�������[��.�������=��FFFD�������p��gϖ'�|Җ�D477����������+gϞ��_wP6��w���7n�4���u� ��JKK�>�d׮]�� ����]lpG�˭;��d7���    �)S�---9V�uÐ�{L,X�{���f���g>ci�=??_{챜�FYVV&����-�w�wȍ7�hY?�����sfs}<�����;�E�i���Ν+_��l�3ʚ5k��_������"��a;����ɜ9s���ݻw_�{�ӧOk������}B�֭[ebbB[  ��l�G"%u�#���"     �f�aHCC��1&���(cg���]�V�6�l�z�j�ԧ>eY�Gy$�J�|��r�7�ާ��F��O���>v�t:�s������f9w���q),,�u����V�.]*w�u��1DD�{�6��*�7l� �:˖-�>޲e��b�K~/�Hh�kmm�ۭ����o���N�� @rT���ԙ6�jd�Ued�d/�$��    �����HAA��1&���U��B��͓��_�Y��;�իW��g����l�2��d�?��?1��C=D J�omii�=�����DD���8��/����TWWk�a͚59��	`���>����F����R�]g�=??ߒ#sAII�̝;W[�@  ;w���  $���"��\G��� �    Ь��I�iikkˉ-������~���t:u���>��OI]]��=֯_oj�L2w�\����M�?�|S�g�u��e�����Q�2e��Z�J�(��v���G��q�x�by�����]"��M�6i�����e
����u�]�� ��{�^������ĉO����vm��I[[�����dbbB[  �<�߯��΀;�5���22J�����_    @v��{qq�̛7O��"w�q�̜9S�9�B����Rɒ%2�|Sjg���۴ڟ��'L���fΜ),�=��FFF��[o5�s8���Iss��}KJJ��G�����ۋ-��?[,[�L���͛7_5|��!�o�Q�^����®'   �Q��w �p     �0���A�ikii�=������O�9���Zx�Sj���T.���B�u������j+V��=��-Z$�֭�=��}�c�4@i�<��c�|�xׁd``@[�e˖i�-��ڴ��V����âI>���ʒ%K���S�N���zm����ڵK[  ��ϧ�N6�Y��\G�     @Djjj���@�i�}�7�Ǉ>�!�|�����J�5��ʤ��Qi�l�t:My(��oV^3�������=�i�^/[��P[[+�/����ի��� �.tn�nnnV��E���RWW�� �={�\�5��cǎY4����k�����0�ES���$�j�  R��g�x<.�HD�4�C�P��;     ��455��#���訩=JJJd�ܹ��@�3Cn��v�c�$��%�ׯWZs�ʕZ%v��ڪ����f���|>����u���;,�������﷤ ���Nm����ذ��Io޼Y&&&��:�c�/���|m�3�ꟹS��c  ���t*Y�0>>.�x\�D�����\� .`�    @'+���������?lj���6���3��[cc��-�H^KK�̘1C�y�%�V�Z��N6�����)�XLI��K�~����F����=��9~��?~\FFFdllLFGGellL���%H"����X,&N��yyy�v���rIAA�L�2���N�:U���d����r���eʔ)r��9S��u�]R\\lj ����'Nh����]:::���t��K6|��oj{p��vKss�����Z�g���b�7o����PHv�ܩ�?  H���UR'+�3Y�5�q5���k�    ���!����핮�.��?�sS�nkk�������T���:�0��{���iת���a���z�2{�l9x�z�/VR'[����A�h4*;v쐮�.����Ǐ[����tJ]]�466J[[���֚��j��t�M��k��֣��P��������NY�v��ދ/���lSZZ*uuu��ٽ{wR�=v�=zTfΜi�T��|�r���֦�4�-[�H4��  ����+��ԙ,��a�^�g�;    @���)((0�O__��ѣG���ƴ>���r�u�ɁL���p8䦛n�=�%b���>}ZN�<)�N��3g�H(�h4*�@@�ѨD"��������%�G


.�� /--��x���6��O~"�P(�:V�Nq9�Ν���>9r䈜<yR���Aq:�������˔)S���J��뵆��͛�,���ب�N�>,���r��Q�P($�����~�_������V���h����N\.�LLLh���Ȉ��W�������@ `y�X,&������+/������ʺu뤹���YD�?Hef���oV��@�:::��].�477���-�3U[[��S��lْ�������,���B��?S���i�i�&�� @j|>��:�^SMW<�h4*n�;�:ܑ���6t^<    �6�����""���ej�]D�����;&���J���t�!���M�6��ݻ������L��v����V���.�r��]>�x<��ښvHk���&J�����7����ڵ+���Y�f��w�-+W���:�9s�ԙ6m�L�>]I�dy�W�7ސӧO'�v^�W�/_.�������8���n������~K��H$��W_�����ڷ����o�-�<󌴵��g?�Y��Ϸ�������t�����[n1�.��;r䈼��;2c�-��/_N�=E���Z�wvv�����y��L���N�����o�[-�3Qqq�̛7O[�p8,===�� �ԩzX=+���H$�v���t��@��;     �%�ӧO��ࠈ�tww���pٲe���I��\0�|m���lڴI���K�9bi�h4*}}}���'/�����7�,��v�TTTX:�+W�L;�e�<###��s�M:@r��a��~ �7o��<�?�P�=��m�o����'?��&�p8,���盧�S���/���_oW6}���	�G�Q��(�G����N9y�|��Tvx2<�̞=[��	�U__�-\@d�ƍ��,���"��?Ӕ���ܹs���k׮������r��a�5k�IS]����	�����U�)Y[�l�h4��?  H]�lpW�P //��;r�}��E�c�;    @�0�����>�����Lm���eeeʶ#�X��p9������O˳�>ky��J���+�����~�3-[�ڰ]\\,%%%
'��'N�W��%��n�*�����`��ںn���^xA���qR���
��|GN�8�h��X��^�x<.����mn����_�{�9����d{;��ƍ��6C��ڴ��4mmmZ��[�n�TPG��XCC����i�it>nڴIk  �:U��%ஂ��QR�D�aIo�c�    @���)((0�O__���;�����M���yd���F�{�9sF�x�	ٹs�彯%���/�,_������Ӗ�N7�5s�L��\^0������xB�
��,��]XX����_�uy�����B��LY�d�J����^�͛7�#i]]]�����t8r�7*� yǎ����e˴��4������9������vR�����~�EEE��9jю;��  ���z��ɦ�{^^��:@&"��`�;    @���&K��۷��۶m��Խ-�gʔ)�o$�����O[O�ѣG��'��|����_?鷵"���/���Ǖ�L$����^i�k)//O�������W�u�l�b��"��}mw'N���_~Y�){饗,Ξ=[y͙3gJqq�� RÆm��:u����k�&�p�ɓ'���V<Q���۵��$����O�F��� ����|J��8�����#��H6�N    ���p8��-�;v��q쩨�����ZS{ ���>���r��1��N��А|���Uvs"����>{����ꫦ�޵k�)u����0��/((��S�*���~�_H0T^7�˞={�׽+NM��^��@Ց#Gd�����3�{�������m��&���Mk����+��|���˙iҡ��p�'   �T�͸��*�@�\�      ��0K��޿��b�K~/
�[o���v�d���j�n��bu�}``����Y>,����)���'-����e�����ߟ��VWW�0ѻ^��|mS��ɓ2>>n��)S����UUU�&����	���hZ�#G�XB��������]����,��������+��l��U�E�Q����K~���K(�x<~�����IS���}LJKKu�M�СC��Ԑ���vy�W������Z�������C|�Am'�����K/���w&(,,��Z˕��a�����  L���UR'
)���@��    ��USScI�n߾}�����nӃXmmm���ϛ�����������^&x��W���e�����I���(�u�V�j��q9v�̙3Ǵ�n����D�$��o�>5���ÇM��~龯��+#��_�w�^K����)��3C�ϟ���b������޽{���O�y�9s�LF~L�m��F�=�utth�ϙ3G*++�ĉZ��]qq�̛7O[�@ ��i=gΜ��ܹsM��+Vp����Vq:���wuuI$��  L����pXI�tpҧ��1�}�}�>�0y    @�hjj��Ooo�e�����ޕ��RSSczd���2�z%	y��7-�R4�_��W��kll��ۙp�
ݧbxx����n躸�X�$��n�ZFFFL��^n�[��J;2���l��4p�2 ]QQaˏ������7y�G�������?���n9u�Tֆ����o굷�k�mwmmmb�b��ybJuu�̚5K[���d�+���t  �u��]o���#��\F�     �,+��x\8p�?��Ǐ�>����9��9r��P�j7n�,�8��~��ԛG�1��?�Z��ҽyf���C��Z�ܹs���l�1��~�#�%��Аe�����՚1c��Z*�B!��,_���׿����0 vt��)9x��˗/����t��;;;�����вe˴�����B�'��B!�����  �GU�=*��6��s� H+�    �3CL�s��ѫ�4����{�1u���vy�L�����-�u��2�ٳg���ג�Fii�x�ޔ��5;p}��	S�X�v�һTn���쇡���������	9}���1�644�t���x<e��p?t�|��ߕ��ݣ ZuvvJ]]�����ղ~�z[ln��0d޼y���Aٹs��Z������gɿ�/g�Q�jh    IDAT�U||]�̙3��tj���ݭl[*  ������py:���/;�"     \CMM��ާ������mz����JfΜ)G�5�2�ʠ�Xqz�����kI��0��������ߦ���ĉĒM�VS����3���7��n����r��i��dU�����;555�j��������������C6l� �CK��k�j�+ۺu�D�Qe�6nܨ-�^ZZ*>���޸��7�  �AU��"���f�5{�n� ${qK�50    @�ijj��ϵ�T�۷��U�}=2���O�<iY/�\��R�Ll�6~+6~OLL���t7�{�^E�|P,3�Xe�A�dFvޚ�z�YR9-"]*��TWW+�5Y�@@���on����Aٿ��1`#�6mRZ���3+.��PHv�ء{  �U��̾��6���Ϋ��H��7     r�]�X̒�---��@�2�>22bY/����ۖ�J5�i��+V������.u9�@@��i�ED���b1S{�W��o�����*X�p���;����jMֿ�˿�ٳgu��
۔qA8����5���e߾}Jk"suww[z
  PO��+޿6��#��H�&���r     9�0K�1����k������Yjjjl���f�6�l�[v�m���fn��_+C��n7�F��|�X�@��鴬���%Pe�ǂ����)S�LQRk��9"o��� ;ڸq#�!""[�l1�{LGG���L����G   iR�Dªk�W���7ܑ˲sM
2�    V��������$�I���[b��避��Vy饗L��622bY��7ҕH$�ԩS2k�,�{�����z��fo�4fnp�
��s�ݺGP���`�d)**J�A�t���������!��������mڴɴ�������:$g||\�	  �z*�i��q[,! ����;     �9MMM�����K�u�Ν���>�Cmmm�qU_�җt��q-	�O�:5�כ�fYť���,�����n8)�3Y�Pȴ�&�:;;	��p8,;v�0�����ٳG.\hJ}d�m۶I8�=  H����+�8k8���܁��]g�G�7��    d6���np9���l�f͒��*�� �$Zҧ��8�P���AWC��Rfn��}�9�L��{%�~�e��%�c��F�Zg 쬳�S���1��֭[M�:���iZmd>  �|�v���P�@���6���     ��!���F����o'��m۶�8ͻZZZ,��
�n��\��³���e������Q^^n��V�>}�e�T���p߹s������[o��{hdv����S&&&L��7�   `�G����;l#�5��    i�5k�������)m�;z���8�y����� rI ���ԩS�~-�hkp��������R<����Z�/+���x�ԙ���~���L��ѡ{h�������@@v��mj�׶m۔�L  ��z�J�p�w�7j     Vhjj��Oooo�o�}�v&�Ԝ9s�����>@����J%�n6��Y��uf����̝;Wú[GgϞUR��r)�3�XL�=��?�)6o�,�XL�Р��K"���}6n�hz�ӦM�t�   ���J��%��g`��eܑy��    HCcc�%}&p���2a�jii������r��hk���K�,�=BZ/^li���A%u�n��:�188�ҩ=@�e�v��*x�e�����qK�   ��|>%u�r����O�t"�     r�a���`z�D"1���޽{-��J�P�ʀ���<*辔���י����ؓRÐe˖Y�36���o rAgg��`�P($===��
�s�NKz�>���mb  ��z�J�Xy��jT����\��0Y���	     j֬Y)m@����M��&&&����� z]]�TTT�ɓ'M��+�D�r3���Lݖy��)�jg��|�+�Վ�b�Նz�aȚ5k���t�����)++��_ Pvl8w 3lڴI~�a����ֶm�$�X֯��S�.]jY?�ǃ3  d6�_w�2�     �����dI��lo����ے�---��+����v�xܲ^~�?����ࠉ�����u� ��[�7ސ={��%iyyy�~�zK{>|XY-�ۭ�V����@@v��%�/�=
,bu�x�����#���㱴/���۷�  (�ʵϫQ�0}�"��$��Og$��\f� ���v    fkll��O:���.K������ rA�����d�0��G���Rݣ$����Ϥ���ҞTV�ʯ��g�I@6����=,
�dǎ�������ciO����m��   }^�WI�����ӌ<�J�,��    �d�444X�+�����%����꤬���>@��r���cz�oڴi��o~S***t�rM���e��Ֆ�=p���Z�j���;��-[��y�#����zR�C�cӦM�G   
e[�]���3�r8�P��E���s�
     �͚5K


L��رci�ضm��i���pHKK��}�lge�]�M ֨���g�yFV�\i�/~�_�q���>���ʀ��Ɠ�Ŵ�2Q(b�v������w۶ml�����}�v�c   ��~��:�p��Y�a�^��}     @hjj��OoooځW+�""������w W������o�����,N�S�H�����;��{N�-[�e��Ǐ˩S���ӹ���ri�d��7�&�� C8&���o�n��  H���+��3���{^^��:@��     �	��������M�ơC�dppPJKKLte���RZZ*�������7@HN]]�|��_�����꒞����ӧO[�Lii�466ʢE����Y�M��ڼy��z�HDi�T�EH�֭[%�����toQ��씶�6m�a>]'   �Z���Su���;rw؆a$y�@"a�     ��c�444X�KE�=�HHww��^�Z�DW�p8���E~�ߘ��f�X̲^v�� =EEEr뭷ʭ��*""�hT�?.Ǐ�3g�H(�`0(�`P��LLL\�Ƭ������w��qV��ǿ3�ȒƖe˲$˖�Ex�X!�9%,i�4��6'%iB�S���$)��_I4�Ґ�$�`��;0���-k�Ͷd˒��c-#��g~�&�xь������uN�il�~�%!����|o�̘1C���$33S�^����IAA����/��Iu�=
)]/��X6����444��͛Mo1b�|\WW'ccc���5B����ՙ�  PL�k���Q%��w`z(��1�@    ����b�5kV�s,˒(YKG�]D�����;�u�-�0I3BYYYڲ�< @��x<R\\,��Ŧ��MWW���K��,��s�Nee%�5>>.��PWW'�]v��} 6��ꌞ   b#33S�:cccJ�Q��;0=�w��    ���ի��:tH���]�v���x�/\._�\�Ν+1�A|(++Sv,�c�;�D����KX�I�&Kn܁����J0�g:��5�����{�2}B   �U�8��)�
�\{@�b��	�    �XY�j�����&ekMLL�޽{��w.n��ɉx�mۦ���� �?~\�n��uM��D�Ԅm$���j�[���5�(
��� @����P�܁��w8w    @,��nY�b��,�w��;wʆ��y6�����+��<�G����n� �o�=���B!��,�ggg����
#�w�y��߿�Hv�]~����/�H��������>S(��;w�>���Ǐ��o�9a����'c�����;��  �QUpw�C�܁���5x    @$���e֬YZ�T�kkk%+]�lV�\)s�̉y�/Q���;�x���./��RL����l(�ѫ��5VT-//7����[]]��Ac�g���2�;{�lm�떖�&�ׯ7�o�s
  bO�	i�e����hQp��;"p&�    ba���Zr������_���ޮtͳq�ݲiӦ����L�15\?��СC��㏛ކ#ٶ-?�яĲ���
�dhh(&k_ȬY��M��M(���Z#�>�/!�1c��]��X���7�}62<<l$���ɍ������
�����H6  �-��#)))�^�I[�Pp�+�~kGܚ�:n�    �nժUZrTOo?EW�#Qo�#2ܝ���lCCC���Fv��ez+���s�IkkkL3���c����\.)..6�$SӘ�Ν+���F�ci�ƍJ&_Fc||\���d��eY�s�N#����	������   b+33S�:���J�QebbB�:ܑ��7*ĭD�    `����v,x��W�^-YYYZ��\�m���#V�����#�8�8l��~�<��1����yƹ�����]CC��J">�k�|\WW縉�""���Fr���e���F�c����ƍ��z   Ğ�b��0��	�iiiJ���b8Ɣ'�3�
    0E���2k�,-Y�*�������PL�~/��-�7o�y��	��������{��6���Y����ky����#��z�jc�@��BRSSc$���<���oƌ�~�zc����Ʋ�g����d'�C�֭SV>�T(�6    ��"�=p�w`z(�    ����l���=&k۶���D����MNN��΃	�@�x������ކQ�v���Sv3�B��ڴ��%�\")))��xgj*sNN����Ɏ����++Ej||\�ﭑ�,Kv��a$���%�)�&Ohhhp�DV  ��Ϗ�;�U��6��7�		L�    LͪU��䴶��eY1[���.fk���ի%++KK�)
���#��g ��������[1⭷ޒ�|�;Zo,8p���I��+�6m2�$���F6��H��,���;�L�^�:��Ζ�˗�V-55U6n�h,?�  �eff*Y�i�I)��C���HG     �s�ݲb�
-Y��������Z��)))�����)��N8�� �LNN���߯�A5'��zH~��h/�OLLȁ�f��G>�c�@�3=a;�Qz<ٰa��|������#Ǐ7��(Q�]�V�^���P($���F� ��N"
�J�QEU�=--M�:@����H��G     �(..�Y�fi�jjj���ccc��;��4��S�`���&��gllL��y���!��/��z�lݺ�����e_|�Ųn�:c�@����2����#˖-3��Һu�$##�H��Ą��Sa۶l߾�H����;�k&�444��許|  {�^�2�H,����Ex    ��^�ZKN8�������*�Y�FfΜ�%Σ� D���d۶<��#r��wK���(����Fn��6�����M�=��t����Ʀ��nϞ=�d'm�����z�����C��ٲ|�r#٪�>���X6  �C�w�=G��
�p&�    TZ�j���Ç���H�sv�����7�7nܨ%�311az8
�@|kll�[o�U�q-�biddD^�u��W�*��{�����ޒ��<xP�;f,?//O�򕯈��1� ^Y�el�vEEE\ߧ�x<F����Ʋ#�o�>0�]VVf$W�B!m�C  �9�&��A%�B��
�p�)͖�Ǹ    ���vˊ+�d555i������N-Y�0��a���9����A��o~#��/?��ttt��Ҕ����{�W���/�O~�ioo7��ӄ�ay�7��a͚5r�wȬY����G�&l����ҥK�d��v�Z���4�
�����Hv�l�6������p*//7�����I�  @=Uw��,D���T�      P���X[�HW�]������]�V�^o�O�E���lLpG0�W_}U^}�UY�`�l޼Y.��)--UvSw:lۖcǎI{{��߿_v��-�۶Mo킶n�*7�x�����êU���_��������8�;�#���2g���>��1�QD�d�����q%�����r�5�hϝ;w����j�~�JJJ�lڴ�X~uu��l  �����dE����Lp    ���ի�e577k˪����}�c1�IMM�M�6��o��,8�� ~�_������Jvv�\z�Z�(����ѣ���ʳ�>+)))�p�BY�h�,\�P�͛'s�̑9s��ܹs���*����Q9q��������Hoo�9rD�9��Fȶm���+�4��ٳg˭��*7�p����˲}�v2�'��lۖ;v��W_�=���.��{L�qv�tJJ�lܸ�X�����ڿ����ɼy�g�|��,�_|�Œ��e${rrRv��i$  蕞��d��U����dE�݁��
.���     	dժUZr��tuui�99-�ĉZ�ӗ��))�����UW]�`G�g����D��p��_�Z:::���ʊ+�ܙ�$>˲���]������n�[222dƌ��x$##�}d�^�ض}�M�`0(�e��ؘ����eY1�w����O��_nt��)������^>���I[[�477Kkk�=zTzzz818Cee���{NN�,]�4�]�VfΜi$;
I]]���h��a����믿^{vyy��򗿌�.@YY�����F~N �$233��㴇���Lw8B$w�P�    ����+Vh�ڿ���Slۖ��F����c��n�:��Ș�ē��T���������������ܦ������-+�";�pzFGG�e�"�Jdb۶���P�����y���k�1��w��n)--������|llL���exxXFFFĶm�,�q7�#���kz�SMMM200 s��՞]^^ww��ㆆ�MȜ���*#���)--�z
�t��n�_c~��X6  �+##C�:N{}:99)�eM��D��D*��!a�    Hl%%%Z&������kkk��=�lܸQ�m��DB�}�0UW����Ǐk��m�ڲ���,�?���_�^���Mo�222$##�B8�lۖ��j���k�gWTTȖ-[��ᨔ�ٴi�����*c�����*���F���|��*��Z�J����d[�%;w�4�  �KOOW������O{B��㑔���?�8W[(^.���w     �gժUڲL����]�,//ג�H(�O]��N�Yh=qℶ, QLLLhˢ��,�`P~��i}����ӹ���d�#��X�z���q(���Z#����}��|���/n�@cc#'�  �DTMpw�ih���J�a�;�W[(/�Fr�?N��    `�t�C��8p@K�{���h+�oذA��d�m��x�X��s��А�, QLNNj�J��)�޽{��3� jnn���^#�>��Hn4L�A��ƌ�O���7����#˖-3�)��-�7o6��'  ��*�;�5�����3���
�588hzZERp����    z��nm���6	�BZ��TWW�%���Ȇ�d%�x/7����x�eŒΉ́@@[�((���矗�^z��6 D ���ۍd�˄m��cSqU��ڤ���HvEE���H�X�B�̙c$۲��=!   D����QpG2���PG�5��"�P�w    �9������Ւ�k����ܹS[��#��ѬY�LoaZt�e�����eY2::�%H$:F���"��#�ȳ�>kz "PYYi$w����x�b#ّX�z�dee��B	Q>���6�/Q����ب��k  `���Rr�����AS511�d
�HF\mu����[�*~�    8����"f�ڦ�mذA���Xs��ܜ��[����a	�Z��|ff����ǏK8֒$&�C��4�-[��/�K�m�� 񠵵U����d�|>#��0Y>nhhH�/M=D���#˖-3�=Un�[��ʌ���	   2iiiJ�8qz�w`:(�;TWW��8q��6����N    p.:�---ڲΦ��NKΌ3d���Z���)������´;vLKN�O�?Eש===Zr�D���HKKӖ����rf;��    IDAT�w&�)�@�25a�����ù�n�\z���M}^Tkoo���N#�N�⢋.��s�ɶ,K�u  ����%���)Uצ(�#Qpw0�7�u��"s�     g�v��ܻ��dhhHKֹ�*����8UN(���nY�p��mL�����ٳ����̙3���:�H4�@@[��^0=����}M^x�	�B���<LMq�?�,^��H�T�\�R�̙c$;
%T���ט��0y`׮]2<<l,  ��Y��2D��wۻw��#*�.�cF\T�    gQRR��X��ܬ%�|��ݫ��ƍ��xjY��ݜ]jj����)((H��̽��Zr������%���[K�h��ƴM��?���嗿��|�_�g�}6i�� ������s��2cٍ���-Ec۶mFrsrrd�ҥF�/��r�3��  0'33S�:�>���������9�B!ٻwo\>]N~B    tMoijjҖu.�eIcc���Ō3d�ڵ�cǎ��׶����tM�>�K.�����Up���גk���ӒC��^ P6�|<�dff�]��?��dggk���w�#���Z������e�y����/�|��d����~�_>�Oh���|�e���v��������e�Bgg�>|X-Z�=���Ikk���Y�l���q�dY�����  �ddd(YgllL�:�1������Q���D2�]�Lp    ��΂�����e�O]]���h���mk)�;a��5kLoA�cǎi�),,Ԓk��܁�?~\[��B�t�(����ijǏ�_|Q����˭��*�<��������I����Hn^^�,^��H��,_�\�Νk${rrRv��i$;�LM��|�g��ݻw� �$��D�ܙ��d�w��m[����ꫯv�/��$�    {n�[[�}ddD:;;�d]H]]�ضك�Qڴi�x<	�B��eY1�cVVVL׿��3gʺu��A�Çk���ʒٳgk-��6o�<-_{�eIWWW�s�D544�-+//O:::��M����z�T�M�X�����Ny����v˂dѢERPP �-�5k��$���9r�,\�P{��瓃j�=���edd�X~�TVVʍ7ި=777W�.]�)�7o6�m�a  `ܧ�	�HFLp�G��]�v��FLEVpg�;    �t%%%��z�d577k�H>�@@��ڴd���G]��qa9///��s�W���1�U������y�B,,_�\KNGG�c��`ppP[VII��,rrr�<(wJ�}/�m[�9"~�_�y��կ~�G�UUUFr+**�䞋��2ZpO���ѣG����Hvyy���sY�l��߭-˒��#�  ��D/�OLL(Y��;��8QWWWS_"���2�7��    8�ΒlSS�����yD|�e
S�����љ��"��G�dǂm��&U�^�ZKN��n��Ң%HTG�і�x�bmY*���k͋����咕+W������w��]�����& d�������JKKe޼yF�-�����n&�p�I�&�سg��8q�X>  0'==]�:N-�3���8�孷ޒ��n�[���&ĸh�    N����~mYSQ[[�-k���QM)��nN���"���1�9��|�#���k$;V8�%���E6��A�^�lذAKVss�� Q�s���Չ���Z���>�|�ԧ>%=���u�]r���KQQ��mI����� 0��g$�lLN�nll���)�������먇�L�M=d   �S5�ݩ�(�ѣ�G,˒�^{M>lz+�E�d:�v    �{��nmw˲�����]z{{�dedd�%�\���`7��ަ�T.���:����6]�k��F�t���L��k�qu:Ś5k�e���jy�m:-Z$��r�<�����O~2�`♩�
�&_7'z����G�)Vgr����ŋ����Hv��   �/33S�:N��>11�dS'�&Qp�3�������q��+�	�:�    � %%%��z�d���;�"i}}���hn�����`'���~0�S�)==]��(�0�$mmmڲ>��O�����\��G?�%khh(aOut	��]}��ڲ�#''GV�\�-��ѣڲ"���%��r�|��ߕ+��2�~.ɠ���HnAA�#NpX�l����ɶ,K��a��*�WTTD6.FL��w�^���  ���"��{7"Lp���{
��RUU%o����B!��Q"�����    8����"���u�.��RIMM��}t�

��.Ӓ���&_��Wd�ҥZ�t;z����
�����,<�|��_V6Y�Bjjj$��0`�:::�emܸQ�����E�O��O�>��ե-+W]u�<���r�W:�`�캻��СCF�+**�侗��qcc��S�L���4�{����x�b�g*++3���'  ��S5@&*YG5
�@�(�Ǳ��6����u�V�輈    H,:�MMMڲ"�g�eI/�����_������h7�w�M7IvvvL3fϞ-����*�ׯ�i�i:���������hedd�7��Y�|�����jmY@"۷o��,��%����a:͛7O���Z��N+�{<���(_����`zLMqwB��d�����֩��OZ[[�dGsR�JEEERXXh$۲,���1�  �AU�}ttT�:���w����d ��*�sccc���o�s�='���iN�����    P��vSp���	ٽ{���Ho��,�eeeɝw�)YYY1Y��+����_JKKc����<��r�-��"���g#;�O�����w��]Y�z���'N�޽{������^k��ŋ�o��o9<55U���/);|��=�5�|���������V D����ȽЂ��'s,Y�D���d[����W�LM7]p7��g�	�� �y�N�S��jLp�G�=A���˛o�)O?���������-E�	�    �h���h��900 ���Z��QWW�-��K/�����ѡ��RTT$��w�lذA�z)))RVV&��s�|�K_�Yy�i��ݫ�����k��V��~���+1�855U|>��u�]r��Knn������,Kk&�����dddDk�?�a����;�x<Zs�'55U���QV�\�=�)��fee�7��MY�x�� �бcǌ}/)//7�k:{׮]2<<l,_7��/�mk����3�s�d���  ���v0T��j܁虿K�������Q%##C���dΜ9���-�����x">�������M�H
�Λw    0E���}��iˊFmm���a-�bg͚%�W��]�vM��GFF���_�͛���ܹs��n���y뭷d�Ν�3g����ʺu뤬�,iJ��599)���RQQ�5w��r�-���>�9����ݻwK[[�9r$�eo��+EEERRR"�\r�\|��ʎȍƶm۔���F'�F���P[֚5k��;���䡇:������_��_Mwk��<��_�BT�F����QO��m[v�ڥ���'�'RZZ*?����sss������[{�������F�|�~~�_�-[�=���B���G{��HYY��\���d���/��Ͳb�
��>�O<�=wѢEZ_w��m۲c�#�  �9T]e�;�x(�'���19t�:tH�z���2{�l��͕��|���WVz���n��A    �3�,�755iˊ����<xP�,Y�%���|�w�h-��RZZ*���r��7Koo�tvvJ__�K(˲$==]f̘!�f͒y������e�ܹ���Do������)���r����_.""�e���������ࠌ����"'�ｉ199��������iii���.��z%;;[�Ν+9992{�l���s;|���ٳG��+W���k�*_7�͙3G�̙��uuu���^��i�Nm1q�>kkk�|N�������ߥ��^^z�%ٽ{���YYY�|D���zc��޽�H�n��fm���ò,	�266&�Pȱ7��g�����nzH@�����OZ˃��`�)**�������Ų`����X�%555F�M���2Rp�����\{��׫{��@ `,  8Cff��u���w z�1e���2::*]]]�k�.�x<RRR"]t����Mk�H
�"�    '���~���Zm����2���~6����l޼9ƻ:���\���5��x��� }}}FN8SJJJR}_z�%= �UWW�g?�Y�z�ڳ].�lذA6l� �@@jkke������*G�QZxOII���ҥKeӦM�n�:�x<�֏���^y�r�W��ƻ,˒��Viii���6���cǎɉ'�> +w�}�\t�E������/---F����˵�M��w��-�����M���r�M7Ex�z���򤤤D��2yB�t^  �A��ѧ��8w z��P($---���"����~�z)((�j�H.��     p���m�`0(���Z�����Nn��-YYYY�jժ)Odu��VDƶmy�W�ӟ���$���^ٺu��m 	g||\�n�*�]w��}deeɇ>�!�Ї>$"'O����cǎI��8qBFFFdxxX,�:��IKK���,�9s�deeI^^�/����ؘ466��̙3�3����=����"�������$eqP����H����.���zJkfyy�ּ����ƲM����k}���ϧ��^PP EEE���˶mپ}��l  �.�KIq��i�N411�d
�HFܡDww����˲x�b)++���&�    "��fskk�c/��W[[��ܹs�䕗�O��~��a�9s��xWP��^�?��?���,�[IO?��LNN����^�u���k��r�(���T)((�z���m۶Mٴ�h�x���uuu��?,�v�2� TUU�g>���,X �-�Çk�+**���B-Yg�,Kjjj�d;Aee����O<�-���B[֙���+�@�X>  p�3f(y]�� N`۶�B�i#���d���~$�������F�dyJJʔ���w    ��-�755i˚�p8,����ʦ|�9KUUU�w�X��������4ZZZ���6� auvvr��F�pX^{�5�{�3g�|��6��?���կ~�r;���࠱��tNT/++Ӗu�={�ȉ'��V]]m�!���)..֖�	  ����%�8��."J�w�ݎ:�Ё�;��B��oJ]]ݔ���vG�$V8lG�5    @�p���ϡ��V[��ٳe�ʕS~�m۶�p7ΰu�V�뮻LoC�_|Q���Lo#�Y�%?��OŶ����O<!�0'��P__�@ծ��z�7��x�����o|�=�hL�c/��2mY>�O[֙����@  ��l]S���򤤤DK֙lۖ�۷�  ΢����+��	���)Y��3�n���H�������    �QRR"^�WKV8���-Y*�ڵKB����H�
�����Çc��,˒��~:!'NNN��?L!4ƞz�)9x��m 	���5�{:ض-O=���=���ȕW^i,���E~�a\b����o���P.\�ȢE�b�s6�e�Ν;�d;���
�l�U�?�w�yG���|  ��
�J։U�3f(Y��SC]�n��y�&҂�7R    ���~��a֖7]�`P�9��7����<��s1ޑ9o���;v,a/2�ڵK^z�%��HX�����Ϛ��4~�_����x��[oI[[��=�_�^fϞm$۲,����o���4�$���!ٷo��l�`���{�R>��Q��^PP EEE1�)//�yƹ�!  8%==]�:cccJ։
�@t(�#�g����s_IMM�lA��    ��tܛ���e�R[[�-+;;[�/_>�߶m�����pGf˓O>)"�}�y˖-���jz	���Sx�&�?~\~򓟘�F����_��W��a����oHWW��| TVV����y###�g�#ٱ~�!77W/^ӌs�m�  ��233����+܁�Pp������M;��1�    	��M��t�,��|aY�<��c1܍�>��S�"s(�{�G���Lo%a�����w�-###��$��//����m$˲�������k.�K֬Yc,��W^1�$��۷�eY�s-Z$.������R\\���ǲ,���1��D����.�WTT���iƹ�۷O�d  �a�{d��p6ܡ�KDV.�u�2{�w    @2+))�׫-���Y[�*�����ѡ-���\��_f��������H/��/o��ֻ�;-���'���!�뮻d``��V�^OO�|�[�J�S�x�裏R�S�W�������UTT$s��1����*�6�$�@ `�����˵/d�޽�>��;vH(Ҟ[PPӇ8!   8EFF��u�^p���P�w$
��&=�u�i��Lp   �d�sz{ ���.my*�,�ϝ;WJKK#z����g�'�����!?��O��d�����%��ַ�رc���������o��f۶<��R[[kz+	�g�q�T��.��Xvcc��l ���~#��,S>v���ٵk���X}����ҥKc���ض̓�  �4�Rpg�;
��(,��������Ȗ1sZ    �!V�^�-���I[�j�'�Gz��رc���m�1�Q������w������r����[n��6ٷo��ĝW_}U��_��阀C�B!���d�֭���lۖ'�xB�x�	�[y��ŋ�e;a�=�,���errR{nQQ�*_w���ƾY�E��,L=DQQQ�u}>��\fn��۷O�d  gRUp�J։
�@t(�C����rIAA�i�w    �T��nY�r���x.�755i-�Fs����Qy�	����]]]��o~S��w�t�9ȷ��myꩧĲ,��q������{���P(dz; �ò,y衇��?���c������{���3Ϙ��iJJJ�e:t�X6�lFFFd���F�c1a�d�xϞ=<�y۷o7��`���h�"��<!���  �������4%� �;�����999�}��t���k:     ())�׫-o���ڲT�m[�����Ȳe�"~��_~Y~�ӟ��$�}��ɝw�)���g��d��lY�<���r��Kss���8�eY��/ʭ���TL`t<���/�?��?ˮ]�b�������n���Z�[y�����a#�@����4��	�&�����Ʋ�,Jcc��l�_s�Ε��R�kN�m��.  �'==]�:�RpO��:�wh䒓7\.��������én     5V�^�-+
Ɂ��ł�Y�7�_�uy��ڶm��o+���������|�d��|����;�{���tvv�ގ#X�%o���|�K_�Gy��_� N��������<������gz;��G?���~��r��Q��y�׫�������1�$�;v9���H
�����#K�.U�^$lۖ;vɎ����˔������6Sٿ�YO@  �-33S�:N���D�d������l`:��Ė��#]]]""��x"[�~;    $�U�Vi�:p�����JbY����h���|��c�E5a���Z����[n��y����v��,---|�d������R�~�\z�r�5�ȪU�ĕdG�y��7�W^���~���?��RUU%����я~�X��I����w������222bz;甗�g,{pp�X6����Ƥ��Q6mڤ=���L�y�%kUTT{ݼg�	F��Amm��AeF����P.\(G�Q�^YY��u�����e  ����P����Lp�C�����vFF�x<	�BOpO���    ���v�e�ʕ����߯-+VFGGe����&����ʒ%K���-�����o����~P>��OJnn��F���K~��_˶m�Ķ����;V5�ٶ-۷o��۷K~~�|�����r�.�&J}}������z���4�% 
X�%���RYY)+W��+��B6m�$s��1�5�ZZZ��W_�����x 0;;�X6w����*#���
e�hO�R����Xv<8�Z���iϮ�����zj��dgg�����(r�   �EUa;Y
��,�xG�ڸ�7�].�deeɥ�(�    IDAT�ࠤ�F�e�w    HF%%%��z��555iˊ���Zmw����h�"'o|�������^>����W_-���
wxa�eICC����k���0�b�)\d>]ww�<����OJaa��Y�F.��"Y�b�̛7����f۶ttt�޽{���N����O �۷o��۷O~�aY�t�l޼Y.��)))�vZ�.�PH�y�������Z���3���̚5�X���� "SSS#�_�Kaa�tvvNk���)--U��Ȝz8��������˕������v+�Q䚚�d``�H6  p���L%�$K��	�H6ܡ�Ǔgff���p�G�1�    ��Β���I�����V>��h˫���-[�L{���Iy������_���b����eÆ�p�ܔ���&ٳg��ܹS����^+���HT�k۶���N�m�qBlgg�tvv��/�,"'�<˗/��.�H
%//O�ϟ︢���tvv��Ç���S:$---��qr6���Q}���x���&''���t��^-ˊ�����뵑^�����X���c"�m[ZZZ�}���xd���RZZ*K�.�H~~���crrRzzz������&���r��A���0���eee�v��)�l���444��͛�g���M{�{yy����gڻw�#�񤮮N���$##Ck�E�d�r�ȑi�c� ��o,  8���VN�NK��w�����p�	�    ����yy���Mo#�=zTn���ۘ���vioo�-[�����˗˲eˤ��@rss%77W�̙s�B�eY���/������'===r�����x�ek%���~�������w�,%%E�͛'���2�|�7o�̚5K�^�x�^�5kֻ�{�~lۖ'N����%����i��9rD�����Ou�������c��|�ӟ֒�}�v�����t�C��M7ݤt�Xz��G�������В�C(���finn>��gΜ)������'��ْ��%�f͒��l�9s�deeIjj�x�^IMM���t�{:�@K0���Q9~����744$ǎ���.����'S���w����J#w��7�{YY���D���Ԍ��K]]�\v�eڳ}>�<���Q�VV��X�BᎦ�  �������;��(�CW���iiiF/2    ��322"uuuRWWwڟ�\.���|� ���.�`P,˒��1	�Bq=�6�X�%===���3�����
����2>>.�e�6bb�"�����Vimm���̘1CRSO޺q�\�err�?��4�Ds�ch�7 sjkk%j��XRR",��G�F����ٲ|�rŻ��Ǒ���4Rp///�V������)Y�(  �Eհ�_Qu���;�wh�r�>y=55Uf͚�:�w     p�p8,###""r��qû�N�P贲z 0� ������n��M���$�S�+**�g����o~�������V���y�wx������IR�***���B�����}>��M'  �sq��J
�bY���w :f~SFr
�^LOII���lC�        �����>s�> �L�i�S .//W���TUUˎG�PHv��i$;گ���,Y�j���L'  ��IOO��5�u����&�TM�?u�)�,(�C�3'����D7E%�w        pv&'��� R[[k��x�b)((���fϞ-+V����.̶mce�xfꡀh�ؼy����(���455�����l  �|���J�I��;ܑl(�C��mz         ���hF�0+
Imm��첲�����6s�~߾}288h$;�544�������b),,���L�P]]m,  8_ff��u(����;�Q6y�	�        ��Tq-n6晚����"~��cS�xgY�����~�x�^Y�zu�vs~�pX�o�n$  ć��%�Ppwh�f��K�]�        �fY��쬬,c� Njhh���Q�K�,����)�}VV��Z�*�;:7۶����Hv"���4�[QQ��o޼���"MMM���o$  ć��t%��A%��w :ܡ��	�         �B������lc� N
�B���eee�mJJJwsn�����A#ى`�����Iaa����	���Ʋ @|PUp7�pk�B�����SpG����(�       ��2Yp���5���������|�)������7��,�r�C^�W֬Y�ݜ]8��۷�  �#33S�:cccJ։�p8,�^����M�Ƀ�vh�RVp�(        ��d�����X6�?jll���a�K�,��������U�Vi���ٶm���HL=DQQQ1��۴i�����x7g���,}}}F� @�P5�=*Y'���ǧ���咴�4��w�VTLW�        H8*��Ek�̙���c,�I�eɎ;�dOe�vYY�������e``�Hv"ٳg�?~\{nqq�^��8!   8]FF��u�a����k3f�P�(�Cu�        ���w�5k��p��	�S)S>��m���ۍd_�!���tY�v��ݜ.��  ���lw�E�	�H*ܡO�V�Ey        p.�@�h�ƍ��8iϞ=F�,[�L������^�W.���;�#۶�M�ODN}���K/�ǣi7�kii���>#�   �Pp�ܑL(�C���b:w        pvCCCF�7m�$s��5� "�e9r���M�$55U�n����I�d'�}���x.^�X


����  @r
+��顪���k܁�Qp�6�&���c        �������������I�ʶ>�/���5��jٶ�(222dݺu�wsR86��   �[pU�N�Qp"G���m�;         	�t�]D�뮓��"�� ��޽{�|OX�l���������e͚5��#b���Ȝ�ņ$--M�nNjmm���^#�   y�cccJ։5
�@�(�C&�       �XbY��=����׾�5���2� �ٶ-;v�0��y������1����&0������/}}}�s�,Y"���sMvס���X6  8��7����+Y'*Y'�(����}MpWV�        	ǶmG�8����[�������
��*++��m�vyy����dj�x���R]]m$��2��3d���F��9!   ������PpG2��m\�
�B�        �GGG��-��HQQ�����\w�u���jz;@R25�|ٲe��������Ȑ�k�j߇�ɲ���15��̇(6lؠlj�Z[[����H6  8����MLL(Y��;�	wh�w        {����.��+7�t����?���뿖��Rq��E�b۶�	�.��	�6l���4��1W�O���K�,9�N   �%k�=*Y'�TMp7�;`�"��+l)Y'��        ��I�S�������|�����19t�>|X%��А�8qB���ell��rB8���û�~8MUU�\{��s+**�^��c�d����J>���i�.++��{N<�lذA{�);v�0�  N�,5�<]T���p�ܙ�D��;�q)*����        աC�Lo�222d�ʕ�r�J�[�Bss����Jnn���e˖Inn�Y�n���S��l߾�Hv2���F
�>�O�{�9Y�~����k�99�����H6  ��x*���n%������fr=܁�1>ڨ��        p>���266fz �T���rIYY�lذ�X����I����d'���6���Ҟ�t�R���7zB���7�  N�m[���bz�������
�LpG2���=-����        ��mKcc��m p���J#�W\q�\u�UF�ED����e'S�k��V6n�h$;�5 �LNN��BDT܃���ut`�;�T�@�pQL      0E���_]KV[[��'ۺu����e0<<�%���7:������Jww����k�]�d�ּ�25�>YUVVʟ���kϽ�k�g����&ǎ3�  NJւ;܁�F�ڜ,��E�5�u$~�S      ���F�/k����� ����$��5�� Guu�|��7�m��������6�F{{�tvvJaa��h��v  �!�
����J�U��܁ȹMo ��VPNW�        HhCCCr��A�� � ~����J��$�ǜ  0/�]�]��`0�d(���������`�
        �������� �A8 ]]]���E8�|l��m�LoA���6���6�  �^(2����*����)YG
�@�(�C+W�R��       �����qu�@�%˄햖���3������)�6�-��%  ���{|��D��;�r��'��)�       �)�Lqp���J�[Ђ�9���   �!���`P�::LLL(Y��;�	wh�
O���rQp        S��+�0<��:::�ȑ#��S�p��A��Ł�����6  Hz�e�mO���ܣG�Ʉ�;�RQp.B       �):r�S�������b���Uz{{Mo#i=zT���Mo#��eJ=  N�j*�nܣG��$��DDjjjd``��6�СC��;*&�+�        H�>��lڴI�^�� p���*���Mo#f����������6b�  p�x-����+Y'�iiiJ��#
����	�3Nr��#Q��        �.�SO=%���gMo�tvvJGG��ފr�p��TVV�_��_�˕x��8 ]]]�� @ҳ,K,�2���dff*Y'�
�>_)))�Z�	�H&n�@rq)��>�?�       �9�����;���!u�ykk������F���鑃��FL��~�[   ���E�s����)��.��;�RQp?1�?�       ��m���Jww�� p���J�[�	��Α�QpB   Π�,m���{0T��.�>gLqG�����ӟ�>8_O^        g8q��s�=q7��z���r��!��Pnǎ����SYY)�p��6�:x�tuu��  IorrRl{��fM���P���訒ut��D��;�r����'dx,�`7         �9rD��>J� n�{kk�������O__�����ކR�  �3����3eff*Y'�>J֡��dA�Z��
���p_`��        ���{�n��;�����V TUU�P�);OUU��-(�}�v�[   ��aeEiS��ӕ�o�3��w襠����X,;q.6        �:::��;���v�[`ȱc��������c����b�
��9��C���ѣ�� @�SU�6)##C�:�ZpOKKS��tܡ��	��pX&���V�#        ��z{{��_��lٲE&''Mo��2a���UzzzLog�����f��P�  p�`0hzӦ��n�v�M���D��;�r�-����~��$Љ�        � ˲��g�������������k�$�y���gz.�K��&��E��(ے;2ǰ!$ b���_��@�|�c8F� ��N�$@��Ol��D>�l)��M��dD���r��ٝ��{O_��=�������Twu��~ ��ݮ��5���_��}�k_�4:>��sU��ML�&
w ��u�ݱ�;L�ш���]���t��kQV�}ff��u`�	�3T�(�E������fi�     {�ٳg�~��W~�W��_�z`H���&bs����z��g�.|�vgϞ��/V= �y�ۿc��3SU��v��{*��ja5�?�o�k     DD=z4�=���㓟�d���`����d�<�L|�C�z���<y2���XYY��_=�|�ɪG�ۤ���8��z�eY�c�ZY�V�U�:�$�;#��p}W8�k�n,�m��w���     q�ر8v�XLOO����Ǐ�ȏ��~���w�Q�h@ɞy������������>�l�#p_����:�� P�����G(EY�q�z����3T��#�����ª�;     0�^/>����|0��x�'��G���?��|��lyy9�;O<�Dգ�E�x�=��s����h4�e�Ν;/^�z �Ӳ,���������R�i�ۥ�3L�3�mc�����ܗ�۱�ى��<q     �u��Ÿx�b�����""��hĽ��?�p<��q�]wšC�����q����뮻|�c��g�ˀ��S�baa��1�����x����hգ��3�<S� ��c[�����n�[�:�c`�pg�jQF��;�8��{��ݯ     �y�����-��z=���b~~>fffbff&�����Ǽ���GЗ~=���cيy�ܹ�G`����o�裏V=Ǝ���U�  {Z�������4���3���ܛ�f)���pg�Jhp7WVZZ�    ��TElnn���fգ 7���_���	v�ԩ8u�T�c  c��jU=B�fggKYg��ag�U��RK���H7	ɿ~����        ��eY6Q��sss���n�KYg��jppg�pg�j%4������W6;qeY�	         �m���#����צ��{��,eu�W	�[9vq9���        `�u��Ȳ��1JWV�}kk��u�I�;쌀;CU�����hu�8����s         @Ʊ�|;�
����R�&w�w��VB�{�[7�����|�M�         P�v��-J`����l)�hp��'��P�p�t�{//������         C�R���v���>���3�Wʇr�sW�c��ʹ         `�Z�V��������v��u�I�vF����E	/��xϋG�.��\         0`Y���U{9���vKYG���B��������R���]_oǅk�>         ���f�#���l)�Z�R�&�3�Um���[�~���G���P=         ���V��������KYg\�S�~��f��+���;y���G�/���         P�<�ckk��1�bnn��u���UE�z�]��l6�V��0�6w��%4�;[ca�WV��$         L���ͪG����]�QEt����N���5��zLMM�0�6w��6��^;����p=         ���nG�eU�1��ӥ���v_�QPF�="bff��u`�	�3\)��}��;�<�]���s        �nE[[[U�14sss��3�_3w�>w������5.\ۈ�����\         Mc�Dޏ���R�ppgopg�j)E�._�w�?r�Z�:{�.         ��V�Y��rl���Y�v�}7+�|��x���(���7         FC�׋v�]�C7??_�:�p�v���#��^ ���|w��7�GD���q����f         �(�"666��sss��3Λ4���	�3t�]�S�]�="���j,���N.         ����f����������j�JY�
eܛ�f)��(pg�j����������v�&         �����^��1*��]�;섀;�Wd�:<�op����x��b��q         A�e���U�����/e�q�:
���	�3t��mkzy����v9w���         ���(b}}��1*7;;[�:����]=�=Eٕ��mĹE         �'����Jμ�#��n�[�:���]-��}@/�G�/������        0Z666"�w��� ���3�w�}�_��}h*v��~�uS�˧���Vo �        �w�Z�����n���+e��f�Y�:0����4��4��{DD��x���fv�        ПN��v��1F���l)���U�;l��;CW�EH=�T�$���d���(|         &O�׋��ͪ�9�#��n)����3|)���bp�7,���Ӌ!�     �'�z    IDAT   �v�yU�1����KYg���a���Z��>6���˭x��5!w         n+��X[[�$t��fggKY��n��N�a����n�Chp����F=�4��        0~��o����ww�w������]ۏs������C='         �(�X__��p���Ԯ�o6���1���������"���
.�\]��W�~^         FWQ���E1���*�6T]F�=��^o��T��햲��;{��;CWKy�Ǧ�.N\Z�3WV+97         �%����{"�q�w�}l�ٌ���]ϐe�X7�w:�R�)�F��;C���{�7�~a9޸�\��        �ލ��<�En��}��}{�]w�2���z)�T����w�w�����{T�����j=�T�         Tc/��#"x����}��K�aii��{�n��u�������4�s9{u=^={��2y         �,��X]]�brl�������cy�RfX^^.e���z�R�w�����.�S���6���1         ����bmm-�mF��>���}��O�2���B)�T����z�������l���z��="bi�_?v9�ݬ�Q         �N����{6��h4��莏�������Ξ=[�:U*#��l6KYF��;C�������^<w�r�n��        ��h�Z���Y�#���Ď����?�w��۝?��u�TV�}ff��u`T	�3t�	��bt�ohw�����q��zգ         P��R���E�ݮz���O|"���wt�O��O�r�^�gΜ)e�*	����3t�"��ѣ��~C�"^=�G�-EQ��         �^�e���Y����䙝����ɟ���������?��R�}�����z��U%w�w�n7�Qlp�n����/��V��Q         ءv�kkkQ�xV�*���������c����{Q��S}��JY�j�=�]=�}���_4ll���/�����G        `������h�ZU�2�:?��?}��=���7���(�/��RikUI��G���KyD����{DD^�8rn)�c!6;�[        �I��vcuu5�,�z���S?�S��SO�����������V��r����8v�X)kU��햲��;�N��JԊ>[���/�����k���յH�e�        �������^��?���8y�w����l��/�R��=�)�|_��ף����hp��p����N�q��ȋG�_��_��ֶ�        `OK)���V���hm������_��?��?��������W�W��'�,�\_��WK]�J�=SU��TOy���j��7l�{���+q���x��C�of�����H��Ջ�V/V�����E��o��v/""R���X��n�cf�[oP�L�cz�����c�w�M�s�1?��    �)����-����w�w ��n����k�Z�j����Q�ף�hT5�@u:�h�Z�J0??������~��bss3z���q���8~�x��V��햲N��,eU'T�V���>�YXnŕ�V���|<����7+��^�Z���W��qee+����wc�ՍV'�zL ؓ��807w�+�~�s�ࡹx��x�ۿ�7�H    {]Q���"��Ȳ,�<��(���(
4 �H�V�F��母F#���bjj*����^�G�V�z�m�v��j�����n�y�Y�C�šC�J_7"�K_��@֭�w�i*QK}6eOț)�5��=��w��z��wm��.�ŉ+�qfq#�_ی+�[��m '+R,ovcy����w<����x�ہ���w >�������t����    ���E�ۍ^��^/�,��!3 e)�Ȳoe�z�޻>�F�}jj*��f4�͑iO)E�Ӊv����>?�p�cl���r����y�c�J��G��J�S��R����A���V�����9��3ӣq�W��"�]ی��^�W�.Ǳ�k��Q΋; 0:�7:��щo�[~���Z|�=�ɇ���]����]    `���u���t:���4��ʲ����z=���cvv6��fLOO���Ʀ���ē������~�bjj�?����>wӍ㪬��f�Y�:0�F���T+�mp����w[������������ٸ��|�}`6��6cL��k�N/���_�o��+o�� {I^�8~y-�_^�/>�z->����>to����ݻ��   ��Ȳ,��v��m�2 �Ê��N����@�V����7���˽�sJ��;�t�]��n�����g�g���߮z�[�|�r|�+_�z��ip��p���_�=��Ĥq}����1ݨ���3�ov:��N���tL5����6ԝ��������W�kǮƫ�#+\\ oU)޸�o\^����N����?xO��S��#��z��U�7�    �^��v;������
 � ���VlmmE�V���阛�����m��SJo�SE�yEQD�e�����&������'>�8t�Pգ��g>�ko���v�)}pg�	�S�~��7��L//bqu+W���4)E�[jű��q��P; �#+[���^8w�o��ݿ?�g�x��N]\���ɹ�   `���"��7�e  ەR�n��n7VWW��hD�шz�>�e���j�����ħ?��GyW�>�l���KU�1�a{$@�D�nV����X�,g' ��-mt��7���K�������`��l�c   ��J)E�e������4155SSS��C���},~��~��Q���������z�����#�N%jE��I}G�6;y�tf9^���\{ P�"E���'�l����9�g��    `bE�^O[; 0P76�5����t�����s|�C��￿�Q"�[ל����kkkU�20�a{�U���o����x���������>/�[n ����V�?��r|��qf�U�8    0֊��N��NG� �<ϣ�nG�׋�R��L�V���k����U����g�ȑ#U�1P�=�T���lpw�2�<��O^�����♕�
�� �Ỳډ������_�K�I     {�`; 0
�,t��g�Ư��F�׫t������/~�����햲N��,eU�T�V���^����Yl��={>�Z�,wQ	 T���V��s�/�.F��@    p+)���z�� �Hɲ,:�N����ȑ#�k��k������������Vr�ak�ۥ�#�Τp���gP=yeT�����K��~�r�mU�� �튔��k�{Ϝ��WG��z    0j�<�N�Y�x =)��v���t���K/�����X[[�9SJ���[��[{��iY�333���J��J��lpOF҉+���g����Vգ  �R���_^�/����kK    ��Nk{���3�" `|EaSހ?~<��?�Gq�ر����j�o��o�g?�ف�k��Ւ/�Τp���߭bR�3���+��� ��q��f��s���r9�   �q%  �#���ի�˿���/|!�|0y�W^y%��?��}m 돲v��ϨܙtSU��T/z}'�>:�6���������_ Tm���^�?����9X�8    0tY�E���> `|�yEQD�ٌz]�oY�,����ߎ/���3?�3�#?�#��{��������x�gJYoEY�������L:w*QK}����n$��_=��\k; 0ފ����K��މ�x�jԪ	    ������ `�RJ��t��lF�Ѩz��r�����_��x��ⓟ�d�����cvvvGkE���7�+_�J<���A#����:��h4bjjʝ��X�T���"�d\��O^�ç��V `����+�^|��ioz   0�RJ��v�(�Y �������TLOOW=��9~�x?~<~�~+����/�|��x���㡇�����<���ŕ+W�رcq���x�Wbqq���GS�Ӊ}���z���w&��;���=%o�T%E�׎]�o�[�z ����։?:|)����7���Q	   ��$� L�,�"��f��Q&���V<��s��sϽ�g��ӱ���������h��N8:�N)�4�����,e-5��`o�yD?��h�D�R|����� ��[����_�+���8    ��(��t:�� ����<��n�c��^/���cqqQ�}�������)eE�T$E�����0��R�W^�G/�W=
 �P�oe�G�/�ږ�;    �A� �k��ee6�äp�2�|灡$�>tO��o,lT= �P��y|�˱�s�	   �xK)	w {R����)�b��p���$p�2�b��4
�����s+U� P��V/���+Q�T�(    з^��{\ ��eY�R+F��;ܞ�;������C��э�]�z �J]��/���   ������ �=���FQ(Vet���	�S�~��Bc(R��󣋑�  ^8�����   ��REdY�� L�^�W��&w�=w�����!%����ŵXXiW= �H(R���v5��   �q"� �6�1J���ܩL=�p�5��f'�g�/U= �H��։#ת    �%˲(� �-�,��Պ��sqw&��;��;���}����k�ͼ� �v�_�͎�Q    F[JI{; ��p�Ĩ���'�Ne꩟���� ]\ފ�W7� `$u�"�9~��1    ����  n.�sw��r���ܩL?�E�1s��?�\�  #���f\�,��    ([JI` �6l�je5�7��RցQ$�Ne�E
���V\\ުz ��V��O�   �h��z�R�z ��V�M�T����w&��;�����S��}P�?y��  �+qm]�;    ��(��� `[��S%�p{�T�^d;>&�97�7��Z9/�  �.��ç��   0Z�l矿 �U6R%�p{�T�V��2%�Ax��� �N���   �I)	h �w�"��'�Nei���V]&��p}+׵� �D��o�[�z    ��, �~�$HU���ܩL-�Y�eQ���, ���qy=6;�Q   ��` @��,�z� w�=w*S/v�"��b@��]�[�8{�U�  c�H�^X�z    �8�, ��E�\C����fܙd�T�V�����'�{��j�T�  ���k�.�    ���v ��q=Űip��p�2��V�}����͊8zi��1  ��V7�c�]S   P�<�#i� ؕ,�\S1T�p{�T�������r�����u  v�s�U�    ��eY�#  L-�SY�f�Y�:0�ܩT��n��E�͙2�vQ�( @�6�qe��7     `�����Ph Pw����r� �L2w*��woΔea�K��\  ���vq��    �c�� ��(
!w�&�����{333Q��J�F��;�ʷ�$���F{; @��X؈n�z   ��� (��+�����]�k�ZLOO�0�w*UO����2��"N\٨z ���   �a� (�k,����{ķZ�a	�S�z�����F�2h w�   `X��  �u�"��&�N�vpOy6�I���.�U= �DZXm����ߡ    ��R� �,�Qc8��r>[pgR	�S����][��ƕ�rv~ �NG/iq   `��� �(�H)U={�w�5w*���B�}��]ިz �����z��   `��� ��-�A�nM��JՋ��fC����"� 0H��<.���   �	�Q `��1�a(+��l6KYF��;�����N�ڎ���� 菻�    0(�D /�$���ip�[p�R;kpwѰ�V  �q��Fd�-    �WE�#  �	��4w�5w*��A�{�k�W�R��*� 0ݬ����U�   ����<RR�  0�à	�í	�S�Zэ��	�
��:����� ���qE�   �r��x 0T��$w�5w*U��z���c�L�{��_�� 0Lg7���m!    �H)	X ��/���^n�vܙT�T�^l�:�n�ҏ"E���A `��"��E�`    ��(�)  [��R�z&TY��f��u`��S�z��'�B��/�Z��
 0t'm2   �$�C �a�!���nM���5���S!�ޏW6� `O:{�]   (�` @5l4dP�jppgR	�S9�S�g[U� �'�E��K��    ؝<�#�T�  {�����;ܚ�;��ۻ�Fp߱�׷b�g! @UN��    �$T P���w���{��,e5�Tn�w�;w��f�#  �ig�����    ��e��I �$�� hp�[p�r�|��7nv"�o�  �N��8�   �>io ���;� ��&�N�������������  �vꪻ�    ���  �Aȝ�	�í	�S�z��'�"�x��rR�
 `$��֊�HU�   ��I)ip ��(��;ܚ�;����m=�ȵlW
M�  ���qn�U�    ���R��8 `�y�ڌR	�í	�S���{鮬�c��� 0*N\٨z    �L��� `T�|Hٺ�n)��3�ܩ\-�Q+z�`�~�	!@ 0ZN/���~    ;��> %6 R&�pk�m����6B�DD��k��G  �t�"�/�F   `{�� FOQU��ɲ����f�Y�40z�	���S�H.���Z'V[6  ���W7�   �1!< 0zRJ6"R�2Zܧ���^f���f$��[�}����v�� I��nF�R�c    0�  F�������{D���L)��(pg$ܮ���5�o�fP �Ѵ����J9oP    0�RJ�%  �$)��;ܜ�;#��ݺ�=.�c�Ջ��n�c  p�   ��d��[ ����wJ#�7'��H�m�{��};N\٨z  n���F��   �V�� �6�k���-��V��I$��H��kp�R�'5� ����,����   �ɓR��T$  �2�E�nN���0u��\��v6;y,
K ��S�6%   ����  ��(
�)E�SN�O��I$��Hh�.��+g��$;��.�  Fߩ���G    `D�y^�  l��6� �7'��H���������휺�	 `,mtb�իz    FLJI( ��p�eܛ�f)��(pgd4��7Y�r��'U7+��uM�  ����͉    ��� ��(���� �������!�vzq3
e  c��w    x;w ��eY�#0�4���	�32�z��:��� `�,������%    ߡ `����[�V�z���nN���1u��<�q��)�-	� �����   ��? Ə;�[�n9ſ�L"wF�T~��^9;�&ѹ�Vt��� ���^p   �[F�� ��������nN���ѸE�{���Sii� O�mT   ��� �Ө��uQ�q$�7�Y�����<��kpWEJq�Z��1  �C�"κ�   ���<��R�c  ЇQ٨(�>���r���f)��(��Ȩ�^��w�����.�tb�;�  ع���   ��J�'  ;�R�����x��7�Y�����=��w5�����U�  �.������7�    ���; �x˲��bjj��胀;ܜ�;#e����5�IF_J�4~ ��,Oqnɵ.   �^5
m�  ��(lXl4U�@�
�7��RցQ"��H��g�����ҎV���#  v���F�#    P�Qh� `��޸(�>�4���	�3R��+���"��{c��N,�{�=  ��̵��嚺    ��Qh� `��ܸ855UٹٝI�����	"��Hy��{���T�V�4�+���W7� �dy�sK�X   ��T��	 @y�ܸ8==]ٹٝ���f���o�v���u�U�    IDATFގF��'�zэ��f+�h4]ZiG��� `R_بz    ��ʖO  �W�F���땲���������!�N��9ooqo�ݸ�`9O�����z�#  P�3�6��k�   �K�l� �|Ul`��j��X��.e���+j�Z��:t��9�j��wF�t��zщ���.�'JJ'�nV=  %��疶�   �!��� ���bc���9)���V)�����8x�`���w�}��!"byy��u B�����In*kEs�w��T4�h�����6 �Is|a��    �*�= �aod��>��_�^�:?�p��~��|O)3,--��D�3`)�3Ӿ�]�^�}+�����K�j����� `����\s   �^PE�'  �7̍��ZM��(+���c��u\�^�G}��4�S&w��#�^�;1�]y���y+""�k_4굛�'�q�fO �I��)�-mU=    6�VO  �g�gff�:���Z����|���y�طo_)3����X��s�����Ʒܧ�x���R�W�V�b��� `R_��   `��� ��ֆ�~s�Ε��SO=��;�W���P)�o�Zq�ڵRւw�����k~�lDʣ��ʿ�b����Q�hc�ĕͪG  `��\��{�(    �a���  �064NMME����Xw-gϞ-e������k�Z���h)�?{���P*w�����L#ߊ;���Lk!"}��������lY㍕"�8uU� `�ey�3�ZU�   �� L�alh����9�'N��)�o�Ϳ���?������r��_��u�wj�����k���g����ϝ�il�_ڊ͎� L��/�W=    2�6O  �7Ȑ{�ш��龏ײ=Z:�N?~�������G>����ݿ�wK9oDī��Z�Z!�΀�nvw��;_L�s.�����襵�G  `�/mE��6�    �hm�  To�w��^���*3��?��Q��n���~���}��s�y����	�3P�����݇<4�uGU'+��b��1  �"�x�w   �I�� `�H)$H�h4��l�}�p�h:|�pik}��������-3;;�������ꫯF�%�H������@ֽ��l�}��@�E�6"/\\  �G/	�   L��  {GJi ����:�5�h:q�D,..��������c�=��W������,�|�<�Lik��T���Fg0/�O<tw�o'��p��Z�#  0DK�X\�fQ    ��(�(���1  �����f3���w����hJ)ų�>[�z����+��+��O��ϧ�����G�GK;W���������w��zw �������=J�ov�ʚp �^��   `r �=eor�m{{DD�e%L� |��_��Ri��߿?��?�������OƏ�؏ſ���:~�'��sDD<��󱺺Z�1U� L��k�x䞹����������&��W�ko ؋^�����]1ݰ/   `�	� �My�G��������JY�u��p�B9r$�z���l4�O}*>��O����}�K_���m������֞j��{�g`�W����e͝  {Q7+��卪�    `��</�� ��QFcz�ш��r
f5���?��?�z�9w�\|�߬z&��;wfq�������?�sT����f�ݦ �����n�   0  ���^��_^6��땶�;|�p?~��1����ͼ��;wram��x���b~fj��6�& ��mi��V�U�   @�����Ph ���&�>??�F��9\����}�sU��-gΜ��{��1�`��٫k��ݥ3ը��}�ި�z�����Kݪ�  �b6=   �/��  ��"��7==�������ʢ��Çǋ/�X���_�����@	�3pY^�����N�9?z����3,/�d  �䕍X��A(   ���7� ����ua�^�����:C��+u=�3���H���˿����7�Y�L8w��إ�������k�P�5H�ֻqzq��1  E�x��r�c    �C�� �!��(�bۏ߿�j�Rg��>>�����]����o��oW={��;Cq���������w�7�v�A8|z9ܼ �^����   `���� x��6r�߿?���J?���x��?��x�W��-RJ�����em��;C�깥���^����/f�C;g��6�q��F�c  0B���o�(    �#� ��Eq�����h6�/wͲlG�T�(�����ߎT����|���U��!��P,�nť����7ۜ����13=~��O]��� ��9ra-6;y�c    p)��s��  �N��933���9o��Ⱥ���r���Ocss��Q�駟����߯z���K�2�^:3ܝD�f���?���m~e�'�V�b ��ɋ�ޝ�    �O�e�4Z �.�<�&�f�����y��׹s����ף��U6��/�����;w`��'���;|bq��<0׌x�=Ѩ׆~�*R�?��v  n�����p}��1    ����-[9 �����SSS�����/��Ng`�3x/��r���Ϣ�j���?�|���/����	�34/�Z����w��7������>��ֻ�   {V���8�yaW$   ��I)�#�  o�ݛ"������=�����ꫯ�/��/ǵk׆v�/~���տ�s�pgh�"���+9��w�����ޑ��m����U� �Xi��3+U�   ���yE1��/  �O�׋z��Zm����-w���O��O�����O�<�V+~�73���/~ơ2��_��Pٹ�?�/~��c�1Z)�"��ʫW#˵p �=�O]��UM    �"��^��1  #�^o������	�j��7~�7�������?�����?�����*}m؉Ɓ�ψ��z����V|��'�S�쭘������V��hʿ~r9�-lT=  c$E���v<���h��6E���c��w0   �=(��N��1  3y�GJ)fggv�N��Vk`�S�ӧOǟ��F�׋���}13���#G����_��bss��)G_�V{e}}��W=�$��P)Ń��G��W���S����j+zy��ϸ��q�Z�F� �q������c��׿p   �^�EQ��  ��n��f3�������jd��'U�eq�ȑ��?��8w�\����=���Fc[�/..�W������?����#�]�6��G����̳"��x>>��}��0?3?����'��Z�[��n�ʕ(�x;  �9yu3^��O=tGգ    �Iy�G��U� �[^^���oۡ����ܝ���^�O?�t<���155�����p�}��q���8p�@�z�X__����8{�l=z4����nJ���;qy%N-����W:Gs������/ŅkC=wJ_~�j���� `w��ص���ٸ�@��Q    ���R�z���  `�E���q��wG�V+m�V�I�ꞓeY�������W=
�J��؛����U��z-�z�=��G����޽�H��������gf�k�ك�A!q��-YB�E�@��($(DI."�"AI�$��	H��U�$Hq�X�0�m�'����z���L�twu���1�������V�WU��I�~�K��o���������7�u⥓�] �͕e<���H2c�   NS�$
�  X��l��⚴�e��ha��6�T�_|1z����<���?)�v�?��7���Y{�� ������s��c    �i�FQh8  �������fYk2�D��Y�

ܩD���'�V���ێ�~ǃ�M��-����Ǟ��F  ,�3W��A�1    6^��e��� ����tR���n� UX~�j����������cgku���j��]�z�x<�箴#�W�^Fħ�|��\�ʲ��(�}\�}D��sY��>n��1� �|�������j�~��������fkqc���V<p�N�s~��(    �(�H���k�Fg}��o�1��q� �7?�{��_}�7<뛿ƭ��<��n��mo��5f�Y�i��T �O�;�鏓�ē���}��(����.�oً�_<���x!k~��^����B��y�_�(�"�,��(^��) `���h4n�aS�ei^�cO����UG   �H
�^�,�W��]�w�� ��6/���F�Qu̕1�Nc8ƅ��������>�T�~����w>����̹�lĻ�������/�D�����Q�\k����|Lc�e���ϊ��[1���zc��Flmm���V4��h4�l6�d��a��ID�   X�4M�l����}~�w��3? ���'�Eq���������֙lv���b{{;��oor�l63q�
ܩT��o=~�/?Tu����{��[/��3��qо����.���י�eL�4�$�$Ilj K7�5��^�z�Ѹ���l6��l���'_����^�:   �Ƙ7t:+�{m�3?���e+���t����u��o{{;���F�c�Ӊ��ﶚz��l���'=+�W���k�| �:���;n7��r_|��wųW:�Lo��ʈ��SGџl��|sk��u�6� �՗�yL&��L&�r�������mw<XeD\i���>�]�   �,ˍ�iL��k��g�S= ������8"^��jww7�͜l�eY�����{o����d��[���q����F�N�A8�Ҭ����w}�=UGyC��[���.�=vb0I"�^c�_�Ɠ/�N)���������1�N#�2] �Z��<�$��x��(�4��,7n�aY�|��h46��   8m�8�x^�?�����p8�$I"���]��3��>��b4�x<�<ϣ^�o\�{��Q��bg��K<˲�v��~nS�V{b0<Zu^ku[fs�������.�7�{��(��mw���~�Cq�5��1K�׼�Jg���v�#M���1�N#�_�� ���(�ux��z������q�ܹ�(
/�"�4��N�    ˖$��	�e��4&�I�f3�� ����<F�Q�F�h4���{{{sF�����l����M�3#˲SL�\:��ʈ�ҙ�_���צ��V����N����b�و�,�4ysk4��_8�$_�ͮ�(b<G�׋�`p��) ��ʲ,��i�F����P�e������UG   X+Y�mD�P��1����d2و�	 �fʲ���s2�DQ�l6צ&�ff�Y������/��h�7�+�&�W�wV�aw��b|��竎r[�Z����w�ߎi�ǯ}�r�GI���X��1����t:ݘ�  �c��5�͢V�E�٬:���<���o�   ���,#I���/"b:�F�׋~��� p&EI�\kn�h4ֶ�UY�1��������u:1�Rྺ�� ���O>���o�{ί_�P�q��{���_��Τ�8wd޽a2Y��  ː$I$I�~?.\�{{{kY(�$I���ev   �Ӷ���eY�d2��p��	 �ʲ��x��8�������[u�ۖ�i�z����6�c:�V�
`9̨g���i|��ź6�����?�R�1n[�$�n����Xq; �M�y�^/���E��UG�-��u   �4$I�v�˲��hGGG��v� ���uR��x���������/6����������y��UG�-W�����|zm��uo  �3EQ�h4��x���q�����Z�ZEY��M^   �Ӗe�Z56��U�F��+� �R����vc0����coo/������v��lF��wl,U��<�T�����ᷮ�(�i��O>�d�g�_(>�3�js `���L&���.\����c��4M�V�E�Ѩ:
   �J)�"�4�:�-I�4F�QL&���:
 �J�<�~��� ����+�V�e�Z-���F[�G�8sҬ����/G���f�~�+���a�1^��f���0z���v ��N��j���j�t:�:�J���'   �uʲ�$I���f�Y������q��c{<  R�e�F�8::�n�Y�ڍN��NwV����'���7���(�룟{)~恵UǸ�,�b4�� 8I�D�ݎ���k�k�Zձ^c~`����    �m6���Y�t:��p�E�  �,���1�cgg'Ο?�L�
�Yi�x��x��o��y��UG���/w����c�P�$1ע�( ��ɲ,z�^�8�|�?>����5��p�=�T�   �Z�nw%;`�e��$����w �D��,f�Y4��kͭ 8
�Yy��⑷��_�t��(��%�S�>Y�Z�to  XEQ�`0��p���q�����Z�������ގ���W   ���(F�Q�1^�(�k�V�� �I�4��n��p���Nq�$��Bn ͋x߇�4.wV�y���RtF�QD^�e�F�8<<�v��� `�̻m���Z�ۍ�lVu   �S�$It�ݪc\3�
xxx��@q; ����<z�^\�z5z�^�y^u$������0����1��ո)��'����Uǈ�,c8��ᡛ& �51�N��jE�Պ�t5��t:�%  �3%��h��Uǈ��;�v:�8::��he�Z� x�y3ң���t:�eYՑ 6�w��Ag����c�T۩�cz9>��J3E�� �����  ���$�v����1�L*ͲJ�    �a�_��!  n�|����Bw�S��Zy�J7���/�4����+Wz���\%׎x�����K �A�����+��$It:�ʮ   pZ��n�f�ʮ�$��M� �����ݫ~�`(pg�<�b;~��OE���h��p?�蓑�?�,��qtt���XB ���i���h�Z������F�\   �4T���eYt:�h�Z�$I%  X�y�{��U��&(pg-}���x�G�<�N�yQ�O��q2<�B�ya���a��}� ΀$I���$NNN"M�S�~��u�
   l�4M����u�<�N�GGG1�LN��  ���,c<��ё�/�;������W���}�K1�-�I�~��x����N�q||�& ����fq||�N�����   �F��<NNNNuRrY�1� �Q��GGG�(�&g^jǏ����/���o}�J<������ji����I���Ȳ�Ԯ �j��1��v ��y���S�   �i�t:��@�x<�����ZT ��)�"z�^�l6�:�ZP���{����~6��Z|׃�/w��>���׽��,��ﻑ �5��8�{�$I���ʵ    ����ڞJ���j����� �+��V1�`�(pg#�����_�\<�Rak���>Y���
���ZWN  ��,�Nu�k<�G   ��h4��x���e�� Z�V$I��� ����G�Q�Q VV��ŋ�������E���#�[���Z��J�"������r7����n�k4!  �%˲�L&���[[[K�V�$�l6�~   �E��f�n�O�:'''1�N�~-  6CY�1��b6����v��zCj�����Ѫs�Z�Td��eć�������LL�;�hY���cO�W��Ff�Y�d2Y�u  �Ly�G��^z7��,���D��K�   ��eY�����,�����ɉ�  �H�$q||��;��(pg#����/~�3�������W�����g���eeYF�׳� �BL&�8>>��l��kE�V��!   `-�e'''Km
��i�Z��K�  g�z2��j\�x��SuX��4�O>q%�Z#��CwE�V{ß����6�U���i���,�� ���,�k��vv��ϻ�("M�8w�\�n��   �*�N'�$Y������;  .��L&�l6ckk��8p&�j�'���U��tpg�E����G?��x�=y���t2���ͧ�XRW��d�V+�,[��  0�ڝl:��`0X��    �����5X��,���F��3� ��(�"NNN��g��	��4���(k�xǃwLz�  hIDATwE��ʎ��I��ПFg��N�~?���R� ���y��4�����h,|�$I��lF��\��    o�d2�^�����<7� �S�$I�i����+��ྺtp��ȿ����~�3�u_��O=�d\�.��CY���tb8.|m  ��,ˢ�j-��u�c�   nW����t��v�Պ4M��>  ��t:�V����� �LwΜ�$����x�p����K�g�G�-�:EQD���� ��L�����ZJ���l�Ν�z�s�   @���XZ��l6���EE  T�(��L&����\�@�յUu ���?��?�֞o�eY��� ���'
E�ϟ_������w���   @eʲ�V�y�/|��t�N'�r'�  pk�<�V���{olm)����p�-�����Dq;  +����h4Z��i�F��v�   T���D��_w6�)n `eh�
�5
�a������D �7����x<^����4�����   x#�~?&���ם�f� `�h�
�%
�aAʲ\Z�  X�^���l���åt�   ���x��`��fY�s;  ++��h��QE�Q �J�;,Ȳ��  `Qʲ�v����2�ݮ�a   �T$I�Ng���y'''��  XiY��8l<� ��(��q�1  ��'-㠶�n�   ,U�eqrr��u�{&y�/|m  X�$I���W`i�Û����  �J�e��v�nQ��   KSE����=���H�d�� ���F��L&U� X
��&�;9� ���N�K�B4�   �HeYF�ݎ4M��l6��h��u `ٺݮ)D�F�G��\�C�� �,�:  ܑ~�����l�Ng��   gW�׋�l��u˲\ʤ;  8eYF�׫:���(�P����0g�@�e1��  w�(����q�=�,|��x��$j����   Ζ�,�6Qy0�x	 �Z�N�1�Ncww��(�vj�ڠ���VDL��ȓo  l��d�ϟ���텯���g   �7+���FU�  �7�����Ύ�Sp�j�Z���X=��mK�t)# �
����  ��g8z8 ���eYL&��c��)�R����G�?��6�ê#  ���f�HӴ�    ��(���U�  ��Q�wD����G��kp�<����  6�q�   �Y2�to `�dY�٬��Vj��׫����#���N���.  6�d2q�   ��� ������)���Ug���q���Nto `�e��   p&�iy�W  n:�jj�nxpp�b�!��zY��U��uQE�iZu  X
s   g��� �TeYF�$Uǀu�TDx"dE�����p��� �&�0'   p� `��߅[�٪ps��x���.�,�:  ,��]   �,� �&s���(�߮:7W{���7�~�\��JY�1�Nc2��l6��4� ���h4bww7�����lV   `!�<��d��X�  ��l���^�;w.�u��p���w\un����>�^qX)i��x<��dEQT  N���V�����ޞ�/   `�e���Z#+  8kj�Z���Ĺs�bww7j�ZՑ`%�e�[�Wunn���s  \'˲�������m|�;w��   �Ғ$����tf  β�,c:��t:�z�~m����v�ѠR�Z�#Ug��mED�j�ϖe��U��*EY�E�ٌ�ﾻ�8  ��V�)X�E�F��    7�eY�ey�A} ����(
�9˺�U���mEDdY��F��3U��*�����٩:      p����bkk��  ��T���ە+W�U����#"�/U�          `)�<���3�Ʈ�1�Xe)           ��ѫW�>]u�ص��(�2          ��eY�X�!�5�
ܯ^���x��,           ���T�[S���""~��            6��j?^un]�U��BD�U          X��,�ʕ+�����k\��`0�]�x�[#�]�          X�O�p�!�=���EQ�/"�ӏ          �����QV���x���{����#�=�          x3��������:��5ܿ��#��4�           ,��������CpgnX྿�ߊ�v�Y           �X�V������Pu�\�f�a0<{��ŷGĻO1          ��xloo����� ܹvp�K��#��S�          p'>�����/��¬� �9�[��j��f�oF��O)          �������(n��[yӥK��Q���0"޺�<           ������*"�������}������(�J��          T/�������PܾQn����#�<�`����w-)          ��\���ɕ+W~�� ,^�v����;;;����j��\V(          �������]�|���������z�.]���Z�D���          �jW˲�7��� ,�mup��p8�������j������          ��YD��t:������W�����{�G�-���G�?���"�          ά�V��J�V{��˗_�:�g!�s=���eY������E�          l�Y�V�p�V��˗/?_uN�Bܯ������Z��eY~oDܿ��           뭌�O�e���f�#/��b��@TgY�׫_�t����k��{"�]��;          �e݈����TY��~pp����N���5~�ᷖe������,/E�#q�V�={eY���݈�          �G�x���_���Dĳ����/}�=�
�d�-i�\�    IEND�B`�PK
     �k�[�ޗԅ  �  /   images/2832311d-4ed1-4369-9d2b-9063d9d0cda0.png�PNG

   IHDR   d   4   |l��   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  IDATx��ipTU�Ow��`��Ȁ,��.�Ԡ�k�NY�E��b�˔U�X3�X3Z֔N���c��
��+*�,�P .D�%d%d뤷���}��N7��D�S���u�w߽��{ύs��g�-"�I
)**�X,��W����hoo�p8��M����Prss%�z�6�G"���!��c�1��X����ő4`�N���JII��L����f�����|
D����TTTHAA��m�Baij8,���{"�=�x�k�Œ r2u�q������&)..V�ɖ"FRZZZ��Ȑ!#p�`�lشY��2�X/�0JSs�,]4Y*J�ˣ�m��P$m��;ӡ�1|��ׇ��G��W����ꫯ���r���@)�I��aR���I^n�'�"Q�pR�\3k�89�2��L>�Y'�Nf��v֬Y
ʷ�~���M���1j�DbxWYY��9R�* ����⽍	?�}��pT~3{��/��b)^tB��̮��Je֏?���ژy���C0]^  'M���g�r�P(�S�ʔ	cdۮZ��q$�� �y��1�w@"y�!�' 8r�jD^^�tvv&Q��S�ʸq����������>Nsڴi
�<�~���t�@|�>ϖh+ߘ�?�{��˘������e���<�u���)Gjj%��1G��R))܄���a�]��y睧&�?���ٳg�̙3�>P-�� 2g���OdϞ=�wq]s�5I?FX�=�%+4������v�vs����-�{�>Gd��q�?ܩ�9��M�:[��8F�$�R����S=���=�����[o��+W�V��@$ �O���1c���<�w���r��* V��T�˚5k��㯯��1c�HWW�466��ŋܟ~�I.����~�A?MN��=t�` L{�\`ԨQ��ښ/>��s���;�t�_�ĢH��H ��TⱿ<��}�'�/���J�;v����* ���IO�3f��Ǐ��w�}W���z���ÕQ�}�M7�9� } <� �'�#� |�ݻw�3#F��\�(��YUU��4��8q��9 ̘h���?�\���_�W��N=d#+�Y�¦�h8$��z��$��G�kܔ&p37� ��0l�ƍ*�n�������{̽{�*3�j�I^�f�����b�x/L����7�Pf�<9Kuu��)�@`���/���zH�n�*k׮��{L߁�[Fo޼Y���K�ٱc��P�T� �ʋdA�d�4���Ѹ/��d���2��S5Sȟ���Ihe?�ɐ�;\p����Ȕ)ST��ϟ����G�������n�ɻ�� �	��袋�^�o�Q���ɓ'�o�o�������4�M��v�;Z�Y��Ga1n� �=ݎ��� �3/a���"5�T�m2ݔt�� #��ӷ퓳� �	�<��曪	0�����Y�j�j �����Ѫ?�P&L���sXh(A �AX�s�Nmk������4.\�PaӦM
Ș��>�H���
ٵk�2�=�8��G,�S�>5>%r�d8	fA���PO�+T�����/���;L˫��������K/�2��(��q	,�p|�����e˖%� 1+� 
P^L�N��I@0�j��4��t�6�dB6�wS�w��Xr�zK�e:O}����-S�{J	��N��^�ӵ���~�Ę��I�A�ޖF�7��ܹs3�� P&��s��0����\i��)�vV>��;7%{�#��f��8�;p�9�/���F�VHr��4�h�$ A��b}T����LW:�~Ƒ/��Νy,��-(í���SB/����}��
TИ�%��U�!������ 4XQ��"Î.G6��S��r��Th��I��2�16�Vh���淴\���j�C��+�"%vU;���;S��!�NH��v��6e�����Ѿ�S����&��ue�D�����+ 0�l����>���P(B8��4���w���x�Q�l���	@��N���a_�b+~+�G�.�+ �$fR�y��q��VC����2h`~�]��c�r��`�s�ȑߗ���gK��A�d�	d�n����A��Q�/1�����äj�#���V��8�+M0���Y�^��;YAS��?묳�x@p��e�r�
���t��/�ݸO��m����ӌ�k�@�D�W4�< lo?"nl��l���ΐj��l=%+��5b¢Ma.` 2ޖ��~(2���hH��=�Y{>��3V���F3�'̌�]��HT���ݕS��T-����z&Ҏ��w�:����%=�H����1�5>��>π��JgQ� �f�g��y�x�1��O'��oOD����%���L���|0�l�;0�� �E���\X[[{��� hGQ�#�5A�z�┌A����W+0���g���:�v ���b�/d.k���,)S��ws��[��r�ߚ����[O�;V�1�܈��.?��&͞�j����ĬAi��O��<۬�B'w�`�<\|��Z�a3�����M�!�źv|:8� �M��/t��)�P�DT���Y��)8���d�7�H�����[�����~^�6W�"���*9� ����=����Sc �O%DB��ě��E���$�A�Lv�p�]n��ߥ����RV�
��rb�tG��sL���,m����b�:�|�Z�)55��[U�s]׷ł�+�	L?�; �N�f��H�a��iQ6Z|��d���(=G�+b�JCm�l߱O��TB8��h���}�2U���g���jNR�Ot�ɐ��u˶Θ9�L�7u�@4����َ��u#̪f�C
��-��"O=����V��P;l�Xy���ppnKb�F"y�pm��])o9�p��w'ϧ�V?Y��m��
Ό>$���$��9�#�G���}��y睚`�%�0��F4�rS�!/��r�k���{Z�H��v����Zk�m�,��O?��^#�>�����MS�}��j(������7߬�t7�5�V`2mXrR̨��S�e��7o����LC+ ��o~�V��O?U��z)�fœk����}��^l81���>���Z`�X��m�M�<���R���;�h����k�0}��D�VB���vg��[P=˶Z�d���ZH&Zq�7h��5A�]v���܏?�X��r�h���{�-4���zg�q�q�Z�673�T@f_Z��O�5{M �瞓�M�	�����Xgo��QrM�m�&�6m��ݦQ��$��bu���cBtXl-` �l;f����K/�T���9[0g<Gf�*(L���H;��I�i��� 6��~���D����,��*(թ�rT{[__'y�i7\t�B��^;�|��x]���v�:�pPJ�a6���_}���I�=�����w���
��d��اm�E;�.]��o�]�%�/>m���֪x�{P
�3h�'"���+�$�N�AC��lդ͍��[#8���,��a��� ���K�=Y�K��u��{�>��[o�	c�(��"������o��� �@��v�Vpn�����R�e)��3�t˷-M2sB������a��(�~V �nfhS7
�����:|�����AlԱ3��2�$�9��܋���v��?Q���>߅%�sX����!���>	ˡ�v9����O�~� {:��2��bbY�,�9Zj[����M��`�}��t��Z������L�~��ѽ�3��C��@�',�}� _�j�<'�2���v���s��"���4�em=�Ś�l�n׶I&��l�g}J:��1���PM	��4vI���SO4�=��2��г_�%���gK�� a� �j^�	�މ�����Q	�������J���x�`�M{u�AՎ��p�y'�Ӹ?m�i�5y[�	RMWJ�n�q�[v7Ȣ�+d����f��PO�'��G�'MԳu�HA�!S7l��
Q\�kE&�,�Ѧ��{��4�#�>. �u�Y�G�}W';v0`�ݑ�1�.��q�r��Ps��j�x�4^��(�$0a�!���/#	ӓ��5�zs�=�A�3NT��ڤ����H1/Gj��P"�G��kAp������A���/t��    IEND�B`�PK
     �k�[�c��f  �f  /   images/c88b2895-5e8b-4a57-9f9a-b80dd50058b1.png�PNG

   IHDR  �  �   ��ߊ  TiCCPICC Profile  x�c``RI,(�aa``��+)
rwR���R`����b
����>@%0|����/��:%5�I�^��b��Ջ�D������d ��S��JS�l����):
Ȟb�C�@�$�XMH�3�}�VH�H�����IBOGbC�n��ₜ�J� c���Ԋ�_PY���Q���Tϼd=#CsP�CT�%���X�}�����ߍ�������k'BLÂ�A�����΂ĢD�33��10|Z����� |�'�8��,������z����j��N��������.j���p  !e�2���   	pHYs  %  %IR$�   xeXIfII*            (           J       R   i�    Z       %     %      �    o  �           a���  �zTXtRaw profile type icc  x��S[n�0��)z^�8~$R��b;^eW�J�ё"�@`H�n-|DI�D��@ȴ�v=L�"�	�s,`�ۮ��z����"H����pz����3�ͬ,9&�h'�tN9#���(���d>CQ�h�|q�k��R�R����mOi�q�6�Z�ܶ=���C�>hrK$>���U`�͚t3�s;����%�S�T�c��\���~�y§b�_"%�G"a=}J�H����|)�Ni����2��yl�c���r�E��|�7$��8��s���.PJ����
��wq�8��P'��j����[ܞ�c2����g�+��|����RM�=�c2gҥl��ϞauTh���҈�\�z���줡㜥   %tEXtdate:create 2020-01-31T21:31:09+00:00��y{   %tEXtdate:modify 2020-01-31T21:31:00+00:00	�   tEXtexif:ExifOffset 90Y�ޛ   tEXtexif:PixelXDimension 1391c�   tEXtexif:PixelYDimension 800�요   (tEXticc:copyright Copyright Apple Inc., 2017���   tEXticc:description Display P3�y��  a�IDATx���|SU���M�M��ޣ {��Dq�����~�V*�~���(���(�"{�Q6-�-�M�{�'I�M������K��{onn���cU{�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!@��-[a츱�aC�5?�q8�^ݺ"���0�
�"���l�a���>C��p���Oo��vn����"��mE�9F�1\���?ۛ�����(:���c�X���_wlP(�ʔ{���=��|+��#}�Y��mo�w��k��]�o�������?�O�0�?���'�Q���W?s��3��"Sڶo�dՊ�}�I���i�f����gf^�t8Z������^d�g`���>�n�q�0K���k|=Ϗ���5�1��}���I0�p]�y��U��'3r��~'_{���G���ߢ��h������1o��v�#�����޵{�I��z�}Պ�ged��x0'""��!;;�߁�������t8�ADDDՎ��4���N����E�l4"""��L�����QQ���ԿTP�UK���	���sn������BDDDՓ}����{�������H/�=��|!'""�c�4a��sh׮ݔ�#F���u�}�?_+.q��p8PPP��o�O���m+�p���DDDG�}ǎ툯0;+k����C���PA܉��\��+z��I#<r䑓�\y���O5�Q�?�^D��R]�]R<�5k����q֦=11Q�s�*Yǖ�Ull,���0�C�Y6'"�`V|֠g�HKKS�o����T���Ύr���������GXd$���(T�:����=3+Y*��D�~2+3K��H�h#"���sx���_����`:͈�����O��;r��"""
f����6.��p�)�ggg��oDDD�����R�7Mgx�'�����"""
n�Cii����p:M{�'��]��QP3��SSѼE�8���,�3�:gOݟ�F��:�������y�
�DDD���";+;ơzI2�kff&���(��j����H�4�L��at""�`&��:���K@/3�^�a�Љ����nC����E��J膻��0���(���*w�^���(@VV���(���*����:��D^^>���(����p�Yo`� ��;w@/;�����FDDD�Mr�0��mPP�ϵЉ����iB��'ԭiՆ.������Q�V�%""�Qt/w���^J�&�΀NDD����m6È𶁴�{+�Qp�/^�T���t""��g߾m�*���6�Q𲧤�H������]��1�'���i��*w""��g����m*`��r���/��Ä�m�����NDD���3��G@g�;Q�S%�Æ����˝��(��3�����G����ΐNDD�Lس23��i�I��S��)U�ge���'{�3{NN�
����%�;Ճ������zdDD�i��K�DDDA�T=&&Ff��Н*�;Y�NDD�L{xD�t�S�:M�~Q��l6;|T�;�&L�Љ����=L��*w�Su"""
^v�a�ax�&�܉�����0�QN	�U�DDDA�T�\J�׉e���U�DDD��.K�|tV�3�|�i�̽t�U�DDDA��%���F��8tV��rK��U�DDDǀ�����t�K���˝��(���K�z���X���(��E�{	��7���t�,��ʝ��(�ٝO	�:��:űʝ��(hI����4�r��YB'""
fv��a�iz	�n?7�)���(�ٝ�sm��NDD��r���SQ�n��^�n��GDD�쐕�L��T07Љ����)U�J8|�r�Nq�DDDA�n+/�K�g@����<����@=?""�F��0;�*��乸ҵ033ii��k�.$'�@jj*>�����9	�QQ��S�ѨQC4k��6���\���1%>�|��%rpq��+�*3��?V�Y�?���Eb��-طo/<���<W�C=��,|��\`�!6&u��C�V�ЫWO0 }��A�&�f�1�Qȑ��i[�I@���p�{�W�܌���X�z5���;�:��V�ޯJ��(��Q�w�{�>)ͧ�Ė���/s0i�$t8�#�=�\|���ܹ��v��D$<�����pU���Ʉi7`��r��s�C��\�U�^�x1�����n�n٬��E�ۆ�)����`�E���Oq��W���GR���yv"��\�g.~��w|��g���;п_?�i`7нN��¹�}�\�-[�b����Gcǎ�p�W�����=轢������i�O��P\p���������O���u����拓�'�S��o�T!����>���2>�͘����3������_��p���T�Y���tf������ذq#��nԉ�cP'��'������ix뭷�|�2]�Y�^�z���'��2���V�{!�Pz^�0���*RS�µ��Gݷg��g'a��Mw���������{���#R�۟���#G���x䑇Ѡ~}u"
Zy���7o&��f͚���8��yHo���;�1��&��ޔ�y~&M�\�f��`�
���hܸZ�h�:�E˖z8Z�*UGGG#7'�z8ۆ�n�:lݲU�TU�[�Z�QV�a����HOKǨQ#� 1�A������K�,��߁�����Qi�tn��lC�C�����g�><����!??�oF׵kԸ1����3���&M��v�ڈ�{o���b�ʕ�a�:�~�:w���Gf ?/~�$��'�@LT�:�Ca�^��,���eʐ�0���or�gf��_�G*��`���9Q'>�>n��V=��v�Z�ϖ�|/C:�5i�H?�~n��L�<S>�\��S�5��s���[h׮n��z�~Y�(�2+&K�"��n�f9U��W\�Á�U	x���s���Űa�p�9�v\-�_+Ƴ�L�׭Kg�;��|2��֮�ù�J������ѱc�ؿ?K�DD!Nt�s����!�{Μ_���~�2�M�!����#г[7�_+O���/�	u�b��aX�l)�36�6��ѥK�� "�P�c�i7���*w]-̀^�n�ꫯb�d�z��L����p�Wb���hռy�Kƞ��u�@����~�H޶�����{�	�_xK�DD!ɕ�۝�i���q����0��)���_Q����p�����FTI0/N�}�Yg�����ǟ@���(�/3p�@*�y�m�4` ��cP'"
9�����rg��#���,F�9Y�.;ѵ[�G�M�VG%p��,2����/�L񲕁?���?���%]""
I�L�곛�k�Ԛ]B����i_c�jo��L������ރ^=z�R�'�N݃~�os�o�X��3��0s�L�{�DFDT��y�"X�X���x�����X]��:Ne��.��� ״������͞�}���[8�2{�u@|�ٸ��K�ɲ'8�w�{���O��������m=�c���xbP�p�ٟrss�����f��u&"B=�ߞ��y�v����y���Cn^���OV}���a+���N�[�8r��!�1�(ǲ��V�Nq�|����EFxȹʵ)p�>[u�rm��ץ���u}]�����OC��:����9�?���"��\}��ˌ���^��Пc�{�hU��)}>޶�R�5RT�y�s�C~J�@~�V�,�[9C�����57"��_@��U�?ϙ��+V�ۭ%cͯ��zԍ�?�7�/&:�^v	�M��C�0���-lطo�-_���Y"v���X�vV�Y��6`��]f��S�P�,�B�Z�ШQ#�n��:u�q�uD�����JZF233��]ۺ		:�*�>��)�f���X�x֩��s�N�I�##"�{hѲ:v�^�{����k�}^ŏ�r�*,Z�k�5۵k���t@����36o��{�@��]о];Ԋ�����u�8��W�3K��t�	�H��r��!���Q�X������u���lչ5m��}ջW/���u�9��a��5X�p�>Ύ;�q$C�����M�4E��ѭ[7$%��k U��{2��3-=[�l�K!�9n۶�))�����C��(�OL�3A��E�ΝѦMk�V���~�:��.�����MIJ�)���+T���6mB�>y��zK�D��f͛��,�u���㐘X��ZT��gVvv���}<p����_�X�����)�T��21g�(��t���k�8t�(���S_om�&���O<�R�>}�]}�������֊����m����ޭ{w�P��螛�J|���f̘����[�nEzz�����u^��t ���x�s�98��S�P%���w���x���٧��U8r%���5l�/��2ڵiS���C�o������
+T�g��>އ�";4h����õ�^�A�����8;U��n�����/�l�2���w/�k����(u�p�)����N>�$�R�ؑ^�/���<iR��r]d��_��*Hz����ᇙ��/�x�b��>>_�͎z�����5�\�s�g[O��J��`��F�ܰdrd�$���q�#T�T�9���u�	�$xUU��\�M���5�'���X�d����Hp�uT�.�6P�]O�ё"��*�W6�{�U�~1#G�ҁ�0��j�L�#�<Rbd�<������ս>Uw�MNNF���zoR����Z�.�1�sp��#�}{���� ���'��o��H׌2*��ґ��,X6�����?��v��#����.�С�)��^��C�`�l�R������;�ޱ�A.ǭ���*�4h�=z�K1�tP���>��U�ɫ3U[����{����z�g����t��.��c�JXd:ܛo�Y�ʮ'� ��%�ϕ�X��$�9[�
y���N��r��z�8�ޭ2�|��~��^v)U�gR�ve�]�b���ٳ����:���q�*w{�6|���0�Ǚ�Zɇ�J�͎��T%���_��u���<�+�ȿ����_�sGvv�_�+�lʾ��5�����y��ǟxݺv-���I�����B��Z�'_�.w�ځi_}�9?��ŗ\��{I����'g�k�|���z9ϕ+W�i���-�����nՏg�T���p�������KGb�*����?�{���K���Uk���̾R�����'[[��>'�dIAa����G��o֙)��L��M�����Z[j�֬^�u��T&��ge�ԯ���(g�pKU0߽[� �=�%~�q�I�������5�گ�GZ����[=�m؀�^{��9N;{$�6%������/�E]�r�Z����5�m��֩��,ǘz� ^U��7����}(���\�;=���}lٲ�����]J������7'��^��=�ܯ��5sm�?5o���ά���:v���)푆V*4u��p����N����|���f�?c�u�!�_L�[�n����|��"�>� /���]ŏ��VJx�n�\��cǢo�^��r&�9�UeXe�sU�-//��<{s][ɠIFsŊ�駟�裏�_����2��-�S�-��⟩��]x��gT@��&��̊ٵ�̮Z��?���H,���>��I����6��x���r�#����D�Х�2���>���:wB��m�Ӗ���[*J>�9*Q{z���믿�^�)��2�J(2���ч�R�J�H<�!C�v'T�%���'�x����d�k����~����@?���B����3�{5j��4dee��2?E�q80��oUf-�Ox�<�$�*�9
o��ffT�|ſ���Gzo�3�up��8���J�/�_R���>������O���$}�+S%57�F���Ƕ-��f�x��r��0��iذ~=�}�\tᅺ�_�SXO���/�£�<Zl�)��m[6]��������۶n�NjA@�����:lM.��t�t�2[�зO�׉�:�\jf���C����໻����m���WJ�Y��d��bX�w��_�h!��^�����_���*ڋ�	Z�1�w����a�B^���t|߁�'U
�4q�Q��-,���1a�J�=U�9�����NJ��= �r]���1��W0��	�ζʼ�������yx�����K/�Nco��^;i(��?��@���u�ȑ#�h�#!����F����9�[f��zH��������|���ū��s��z�
���zg㪫�
�gYڌ�3K�b�c���+�������Ǚ?⥗�cܸ�������eR:����ǝ�Tk��g��Ѝ�bz͹xť��`Ϟ�^����B�.]t5o(]!OR4��Y:t6o� ��ê ^�~��8ӻw4k�u���UT�h��]z���˖��]	��=gö����Ï�k{�E��T�ק�~��%���#"Ѵi3�B]Su���7';�R��Ҕ�n���VS�JЎ||�ɧ8���|�
_/�]	hLl��h��m�"11QG����uo�;v�;�Yg|�T�H��E_�.�W����=u�4LU%9W{y���D�=M�4Vץ�>o�$��RSS�a�l޴I��[_W�2L�:_r�
��0�L0w]���u�4G����u��n2�Jz��]�V]�dx_�X����(��N8�_�������ȑ��v� ���N��B��I��K�.�3�����Qڵ7oެ۶�'|��C�.Fq6=���=�;�^�I�$��t�2L�<����\ރ|O۴i�{�K�HG�C��r�򹦧�y9w��LӁ��}s���c��A>�G���}��/��\=�7mܨ�[�d��%�ף�t�S�֭[6+��)s���2>�����ak2�H!�ک��H 5��_�|9�?5��`�Db���T%�W^y��#פtu���ԗW��M�:����k�Nx�;�oÓO<�F�h�8Ce�Ru tu�+
�R��ۯ/���J�v�ih�����̈;)q�P�9����oM�R�1�f�Ϟ{n֫���]7�
�u0��3p�:N�޽Ѥq#=��s9���6�k\�����}{���#Ìf��:��^��"�>R�s�v.
�a*A�ޣ7�P���[�j�;W���W�dΤcۤI�����e�	�34t�x̘�طgRS���v":�N9�\}�U�qӦMu	�s]dH�֭��ݷ�����W`���"C�O���}zW����3�ǘ����yp'��o�駝����,���!�1�S��߅�����Y�,2K�s�{]VN����y"����}��ΕΠի� g�u&.��b=�q�ƺ7���zA~>RTfm��%�����H�Qِ�o�}�]�pB=����m곸��{p�-7���]���;u������gj��Q#1��u?�Lɐİ��?��kf@�R�+���D6Х�P������*p_Ub'�|*~�a�q�@Ĩ���'9��x��W�������6g�l��X��mX�z%�W	�۪�Ѩa�J't�P�\��T%���;q뭷��JPQ�L�p))�҅<������>V��t�Q%�����[���x��Gq�E��P��8R"�ݳ�w�'��?��*SeyUR��N�m\�а�8T`�*�G��"�*�ȃ�Եi�Jp�+c�\��-[��u-q�
�R��
�e��B�u��l�kޢ�=4LW97�_��K�jת���ҹ���N�ñ��?��IUb���{�͚4���^֬߀ѣ�ww����'�n��s�mh�2c��:��&������Izʿ8�E/�(ٰr�r�S�O|�Mԫ�P�{]�냅�Q������O�Ї���멈s�m�y2��|�q��aʔ)5r�:�����$C�j�9��nE�Bf��Gq��Յ���2����4��>A�I	��zg�'�q��ϬH�Zž�b���u���1}��qc�}˻C<��&g<�[��c�=�i_M��8B�)�|�ɧx���T�V�6j�Q�G��7�Ꜽ���R%����믿�vxz���T��^��K�DwZ�VaoǑ`0d�`]���۱g�.��lܸIWG׫�$.֊�K|ݺ��8����I����[Ǥ$<���X�n}���H&�ƽ8�{��1ͅ-���?U�1c���nƖ�-�c`��d=#�t���a�ĉX��[�թJ��1b�H]����ɞ�V_]O�II��V�	V��3f`�*9ߦ2��Q��J��u�_��T�3�9?o��!�Ho��]Z��~oSKK��|��:��^��X锸��Zzj|j^�9bz.w��멚�)N:rI��+�['P2�HL%&�6�i�ܵ��.2K5�u7p� =L+�]�#z�����J��t5���H{�|�ǨK/��\gW{�C���]����ݯl'��I�ᤷ�*wk�.=��`^ѡ���:^t�:�D�g=6X�z�J�+��;�w�q��ů"ץW������1F�t}��H�[O<�.8�����{��N��T`�>��C�aݺu8EmW���]���-��V�e��O>����+0��g���L{����t�{�+6��hˬ��z(��g֥〥)�|��a�葅����h*�I��K/�K�,յVs�H��c��	�N���Ց]���g��m�vM_d�p/SfVWs~��ŋ�[0�j��숃���V�ǞxLw[�'�([)�l~��ttx�� u��8��tӍ�ڸ��A�L�������mE��ύ7݄s�����9IIpР���O�x���1t�=iK'��֝�RʖL�ۓ�Fj�>x���J\~�e>k,���*�O�4��C("7JG+����S�#S�Ju�Ν�U���|�M�A�n+̋�Ƌ/�Pw}a����$C}��1�����Nt�p�Zb���W^#�j�G�)S�m�U��y�f�?p $k,��Ͱ�۳�&��KG���l[�V��P�i)��~��7�Y��~i�'�T.��SN�|;�����}�}�a���k�������s7�p�n���qM=%�u�]W���:w�&M���`��G'Z�l��.��2:$�~b}��f���A]�&"#�����)�Oj�V�Z�:�y�xm�>C�u�Ǒ���w�5)P����蒤�NS�*	����2��:wŭ�ݪ�D��.���o���f��.�+K��e:��^�\���0��$��a�k׮���B�{��]��Cꚻ:�ѱbJ��M&a.GMkC�_:Qe����B�+�ۄ�y���$\q���L��OI�.��=��?�:�X�b��5hr�9�<����uĀJ�엨J;�u@_�u�SO;�U��� �p��z���L��U-��V�[a���+���ؼE/S|��s��ǣg��*�JB����m�uQ��^�s��Uj+�2�aa�ͼC��z\�ަuk�{޹z� ��ҿ�.�M���[�5h�Hw@�L�kO@�*yw��	�M�n����̬��б�>k��]/�jb�db��[J�6�`�=D���3�:�[�
h��Kz��w�y�c�UU����0�!�^}UB)=g+P"UF�a��^����r�#��.N����72C��- �>=z�@�J���u��$��ye�лO�J��/���KH��uY�C:�z��(���3o�<����^v��F���,u��x�	i�8p &�5�G��ۇ*�"�Kf�c����(�;YAN'���*s��"1tL�v���u9�����M�>f��ܵL�*�W�L�b���:2ɔ���B�F�4i}�7\�c,XY�K�}9���B:]�t��{��_�׶BSO��1 �Ԇ���qb�>/A+�g��IV�mV�5�ef�U������U+Cw2S׿V-�m��zQ_v�ك��Vx}�k�nh߾j�Hr7M<����J&ϑ9�s�n��^r�ש�������"B���VMcNgH��Ւ����yU��n��sTt�ϭ$G*������٧�`)Î��z�Y���j��ڷw���n٪�l.=����� �+KWT��{�ԓ�4k��e�����H:�1u"ݮ]�J��}]t3���A�?�l��%ǩlgTڶ�ː@���;�`0���I����K[7o�|�y�w53+���m�Fe
7O�d�$3lU�.�Ռot4�_˫r����$ш�Yb1��4W�Ȕ���ɬ�i�u}TsV��]R�����<�b�0��;v�eJ��(qq�t'�ʒ�k�')=���y?�u*�픡��&ޛD\%t9Ve�U��쨌M�7##����=\��[Uj�_��d`�e|v�ڭgᓀ~dLDFE�q��Nz%�*ڼ-��b��/�$t���g���3�I�!���*s�I[]%�Ƃ��͝��Y��4C��I�oU�	��!+�Ig$�6:�t����W+N=j��IЊ�=�Z��k\�V2TU-Zer�t��*S)&	�nݢ�}�H&j��=���_�HaS��L�*�Y��?x�S�W�8��A�@L:TD������YCg&~U���JJ2��M�����۷O�U�w��`���4�eɼ޲�CU/BӴi]��(�8��;��[��.�?G��X�(U:�N�H���Q��H�������܇�}޷G��YO�����Ǐ�믿T�o��ѽ��z�����d�1�F��(8I	�^4o�L��]KJ����MWz]=��i�suj);�7�����/�yJ�99e�2�:Oα2w�T�JG��&�;F5J�$�v42 R"=��M��R�&��x#�k2��q6e�&5��؏�d����j�k�#�\m�5�m�Q�ƈ�]���:�i{�w��`&��[�M�*>
U��1���Idsr+7,�nS�+�����]M��W���e<���X�����z�Uѩ��jH	���n����dLm�zu�o���.;�Ɂ������O���V��G��*@Ib���C���l5s��J.�J�*��<�f"W]HG���e��@u�*��d�;Y����r{��jh@o�X퓒�F�3^�kv$Y6P��7o�3e5o��u�`>?��>�P`��+\��U���Q�*��SNUC�1G9��qk%�Nӽ�0���pk���a��򎥚�gϞ�V�;���˗/׳N�`��ʒ�F^}�5|��7�бz��޽{��%�KOfo3_IU��`)�hf��0HR��g=9�!c��5>�'
��L���C�v�\�3G�f3u���@T1�Yn���5��^*�K`?�a=fu��eض-�:f��#%g�/%EO��c�6����l��ZĐ�3z��K/����)�N�p"	��(�H�`)�W5�s����OT͝Oǎs��
M�?��$&�?f��:U0��8ӟznC�u:N�n[`��(�mHNކ�9�]�]��7�B<�*=Ʒmݬ���ڷo�zi����A�p~PzȘ*�gdT}�_��Z+�و���Ы��`^+�{'O�0J�\h�8��TT�Mu�H�ʽRU}'�zY����?���_�e��]	؇���%����t򓕮�ԫ[O�Ѷ��(��Ν;u�۪v�59���v��1̍f63�٤������Y����mT�:1������]޵Ls������U���v���_�d�R8�rF[�nÌ߫�J�̭>RS�v*���� Q�������*K:ffe!.6�J����]�N�L*Svq9������m�2��Uږ����۷��~�]���R����ft���;�-^��k���Æ�;vbʔ/зO�c6C��gb����|�z���#q֠Az-i�O�^�zhּ6m�^�e�Mz�}\_s-������6��u2;�$x�����BNN�I�d�����K.�Z�%yd^�#��n�Ն^3'��%k�r�U)}���^��u��]vN9i�Q�b��yr2>��s���d6�����mZ���O�܇gq����1��_,�"��u�֣e��
[�n�ƍ��mXY�֭u��(ڨ�^�nv�*��|#d	S�z������H���.���R� 'AIa�������������t�m6\~�e��/�q�:��ٰ=y^z�%t萄���G�)�L@1y��X��?�7��s���0{;�������`�1�Х��Qe
N+LtE�i�쟱{��>���٫�^~��ߊ �y���T@�a񬁕+WaŊ�8픓z\��������s�~��*cQ6@�&MФqc�h���:�����N~3u�	[yU�5��]�}�Νqɥ�`��qz&'+�&M������ȣ�e�i�l���{((��L&�hּ��'A��9���[q۱}�f�*���]wމvm����ٻ3�NG>���ckšO�����}'R �=$�����s����>uON�2����.\�_���Ԕ�أ�d/:��]�>�p�'�se6s����巽BL��:/l�
�W]}��6�[��e����+HHH��s"�ë얔m�*�?�̳ػ�[�z"��.��{�*w�R��ۯ�;��f����0u�T64`S�����|K/���ŤI��úw>ё����3�w��S8�����^ݗ�^���k ��r�ÙY���U0���;��2�UI=�S]�h�����z�I�YN�l2����~�m�a�S��p���؟��}N_��o����W�|�^�/��,^���dNt��7�|�.e�:ݎ^��?�|UZ����&m�'N���N9�J�/9�e+V���^Cf�� ({+JO�s�=͛5�B
$��ڧo�4�GX�1�=9/�8mޜ����W|e�Q���o�nW;g�uV��i��ЭÏ4�y�d����Ə:sJ"\݀7� ��*O��+/��6]���O�^<p?ڵi��	D ����3Ĩ��x��`����E�.]�>�Yg���y�υU_��[6���c�L%rmZ�:���j߇^��*�[�V�hѪ.��|]�
���O��UW_�y��!+Ӻs܌�CR�x��'sd�Lxz��^�cǎՙ~o��N���5ADd�^��j1���<�Kܒ%�ωe@p�v�����ª���n�{�X6d��a�oa��ŸM��SZ������6�I]6mقw�yWW��L���NJ�W_}���
�۞eY
��oT���*�;�����J4�0t�0�ya:�kW�DN��c�.<��p|�ŗ��l�$,,�^{-�w��`NU��s��_���V�z~~�|��G������n|���ҫ�ɧ��?{�j�v��|��hP�~���ccbi�?��}���3rM����t�SB7ٖQ��XRU7��0l�CؽSz�Z}A}����O=���'�����y��'�u�V��c^r9��,lܸ�~����5V�Ҭ����X�W<s }����}���~��3>��S��e%��_���}��GqҀ�^�&��Zi..Z�J*���7��/�p��	'���E�������{J��}��WGw��.:s�����q�
�����"G%_��Q����g��Y::{�ٺ�����w����<k�̾t�����z�T��n_���N�e�U�Zn	ݕ蒇L6q�嗫l�	��jއ��Ds~�	���;Z�j�~���G�����84i�1��:�K)\������{�`ٲ�X�d�.�oS9��Y�|��LO��1ϣm����}݄x�Y�իWc��%�J䤏��ٳ�f�\}�5�����!)Ig ��N:mڼ	ӿ��>�[6m.�WYN�l��?��^�`NUi����{���#��]z���eMM����q���~-[�@���}f��`��ǧ�->��l\���8ѵ{<��Cz\zM����j�ɢ֭�z���];q�}`��i�ԩ���9����ߥ�q�1��+�ak�r���6`�ZD����_�uz���F`�~�+odC��v�����٧vĨĠN|��)�H@�ǲT@Vw�����}�߳|�I'�ŗơO�^���ӫWO�5��s�^��[-Į�;0�����T/5+��e<�L#����g��)Y�p!�'o��᫆����`��0���@T��b-*(�y�ر};�y�/C@��z���xRe�'O���w��4j�	ut'���=m�r����زe�*I�.��{�F���SO���WMIg�}Ʃz+U��s�^�ru2���4���as��2q�i������G��T@/�#�蚢*\����$��z��c\r�˗-��Jg�[��d!�Çӽl��J���0���{�y1�Yt��9 7�9C�F���裏b��M�ԥ��k�v��~�=�UxD�c����<��Ư��M�5�SÇ��T����hеR*0H&2?� ���C�v�m�#遽i�z���˯��uהφ������3#��y�&x��q�X���d������u2
���X|�\������{�a���HP����z�Q^���ß�Rsx��e�^�6mZc��Q�q��ɖ��\+o�:W�L�ÿ��[q��w�I�FKdH��a�����ß��E���^)z����I���ʕ[�ҵ�J܆�63���&%ntlɽ�X}wF??J��ߞ�6�I/k�Mi�W��*�+�[^F���mݦ-�����
�\�����G��X����f
�))ػo��Ŧj�
��k����={b�ĉ��������H�|=�ze��W��SO;��s7�W���$��;g�^Fv�8���-2����U�9�s��:�	���K����ݺu�Čp�3���^��:�=��Ӻ���W^����aZ� X�E�ʻ���=22��q�}�����DU�]N_�#�=���{?v�H��A����HNN>f+\)���ˣ�����?��ުґCf�[�j5������G���!O�[OO[y�5W��s��OH�۽kL��:��x������,l.�H�M���O���O9�]w�^�F&�����^!N����5Z��W�������@�S�Z4���q��^��z�Ksp�	�>����*�e���G~y]lt4n��z=c�dοV���7��~?3��C���
�Q1�ر��Tw���6jРR���Ɏ�{��^�Z���bu<��qD��Is�|��F��}\(oi���9nӦ��=Opv�A�Н�����Ti����õ�K�L���m.���lݲUw�������HH�G�vmq�	'b��A�ӻ7��M�[�*Ty_҃]ޓ�������3�`�?ر}������К�fG�
�mU�\f�2dN:i �={+}��^�[�e�v:�zᜰ��Wmʾ���t�ֽ�LWr��I�V�!5r���֭[�kWu���Ǒ��S�Jur��=�d�%�v��!`��ʔ��{�,�w9���� ̋.׿Es�믎Ӷm�A�Hy�:��2r�sz����9?��ʕ+�����ɽe\
Oa���Eb�D����w.NS%r����Vi�٣�
n9% ��e��/=���tb릮yZڡ��/Sjk���W�\i^�fK��|���i�Oزy3���c��B��Zj3dTP||�����K����]],�J���մNG�s��gC�t�8�3t�;v"y{�^&TƖ������Y���HH�ڵ�PO���5k�\y�W]�fw���[�9��&w���ur�v�Y�F�N�e��Y%#=]�Ws�$*�j��^f��ر:w�W��#d����׫�	Z2���$�뮻���V"""W��+�I���>����QQQ~�ŕ��qϊ]�#>@���S�/�r�p��}e�#������-7�d��|b��+}lԵ�N����6m�ڵk�z��}�����lnn���bս.�=˒��ڵC'��v�{�Z�Z�
��s;��S��w�-kO�\�����S�|��/-�%� _��C�:�����Sqݮ

�����~%'�:u�ѨQC4i�T��1�2�S�
Ԭr�"�W݌�*ˣg����ِ\���5���@$��A)J%J2�Qj�����_��%�o��>�]� C��2w�zߒ ��� ��Ë����}�u�Dӓp�:�ʪ���qU{�o�VD�=��������"�LU}��qq�Q��)�/�I���&=ⳳ���ס�}��$�(:yHf˰�O�H/����r�;P�7��aUu<O�Tc��Q�9��k������΀^)f�K)C�\����b?�w,��#��L�im/��;�hݥ��8��|��8ގ)�ňp�z�����<��58��0K���0�~L��6�@;�\{u�yy�PM����Ni��f7����YB'""
f�S\�[y:�Q�ѝ8�)������^����3�-ӯ6�|v�#""
b���������(�ٝN��ֈ���7=S\�[�,HN�Љ������W~	]�9:����T:v���3M�r'"":�����,�Tn�7+�O"""
�K�ݯ8-%tFt""��d��m�::QPR1����DDDAKW��UBg�8""��e��˝Et""��U�:#:QP���U��8t""�`&U�~lU�?"""
F��ΈNDD�̊��3�)݆ι܉���;��~e/w""�����,�NDD�L��YB'""
jXm�m�DDD��"���������r�z�DDD՞S�r�5""����U*�}�k�r'""
ZR���VN�f,'""
fz�5?7eX'""
V�ߋ�0�'��,�U{�˧2�5?�r�܉�����m�r'""
b��U��DDDA��Nq�����(��~W�Q�b�;Q�Ǚ∈�B g�#""
~�C�˧2�+��^��DDDA���2DDD�ʏ�\�L��NDD���ΨNDD�����*w""���*w""�`�ʝ��(p�8""����kb=S+'�܉��B ;�U\m������K�p.w""�����\�DDD���X�U�DDDA��Q��LqDDD!����,DDD�*�˝m�DDDA�ɉe�������CgX'""
R�
T�Q�͉e���B��m�&�܉������6t"""
F�U��Gk��DDD����܉����
t�#""�`���WЉ����Dh�m��(񃈈���aT$��UBw8�HKK�!�p���� �`PS
Q���c�=�l����j���둓��ז�n��0l�C��Wæ�5�������]8
�������p����*�&6���e��-�8\yS~U��^�t1����h2�g�.��6��sDDDt�I��f4��&��� ""��JJ�:�烈���+UB7��͖n:�� ""��Hfsأ��ege�U;6�-3:::�^�n��������{�g��0=""�I&������K���;w$�Өqӻ<�t^^^/�4cTD��u�ƪ�3*8���c:1ϑ��g�#|���g��OF��x���$�����jժ�y�����W�<l��k�ŧ�O����;v����LP�F��]mn�G���E��l6�&m�v��0�æ�`ap�4�����rd��ϫXf��Ta���
�+����ſ�F�_JoWl����l�	�Q�k1׉x����󇢿B�8*�g�J����b{/���}����(:f��Qxn(���.u��{�`[�~���0T�.b�ҥ�{v�
/���G���NC�&M�T�^n7TWr�֬Y����[f�������=��ILl�o�Nɟ�f��MX�<[Q��}y�~����1�\4%�Y�wϮ�����,�{������vW��3K���yxv�c?%�l�Kb�R��\��W���)|q9��,q%��[����ĮK��}���n�a���{��_�]�r)�'�z_/)���N�l�b+��(�-6-�Y�b����J�-��ڨ�9��G�}{ΧԖ����t��pJ�e���%���-:�b�G�J�JM����.rџ�ݠ��:IϹ��\�������0̘�hg|BvIIs�����Saw���ʇ���G4�΅�Ϡ ?W?j"�gY"P������Ӑ@�p��ÐB�l�S�t8W pr�����T$u:�Õ��p?����w���&���\]$�b��$�o�^ܙ���kѾ����m6�����u�]o�ٽ�ً\t�Ÿ��[Bnn�;z��͸�λt"Q���N���on���'�<�������OOL�<O�EyUw�g��&�%�f�L������õ�Y�I�?\���u����hY<u���	S�,�;u):/��s�]6
ӛb�r�����
_��G���R�����̰�^����kc��4�ͦs�6Wy��-5�0�\�����6�]^cs[�e�._�CA��o��0RB�zHٿo��>�S?�� O�l٪UH��7�

���Vtx�is8t��4��J4�m�j��m�w��/�(5�_�O!_ega2�J%J��#��X�]<�g�إ{�i�'6�^�٧�Lexb�Y��Z�;�'���|��������Jl��2y�.�-�܌Ȉ��Zu#WD ��x���\���j�ژ��~̯s~Y߿}���E���[_a��p�2�mW|�ҥ�R��(�P�F�s+��(��/��(]�*��2�M��x�k�9��?ós�t�<�t�B�{��#�?=�Og^�{Tx6�k��F��'�����ܙ��r����w��=��M\�C���x�y0e[��|�}������vU��2��pU"R��Ɂ�
��c8�Զ��r���گ�S������r�Jt�ܹ�ug����e�,���o��� ����W;����"�#

�eF���e���سgZ6o�/S�T婌���o�c��-]:�mҬ�ks�u���'`��u���+AD,Щ���T<�$$$����J��ʬWr[�l���kt@�`.�;���*CS���f�^��?�>��t��6��{�Q0a@�2ڷh�ǞxR�����v��V&����a�?�`��A�>������_<��sػG��R���Jn߱ø���vh�] "
F�d�q�&�ݧw�_|�^�ڵ����������:��m;����x�駱j�
������f͚���/s�~y��6�w�� "
6�d)-��p|n���V���]*�J[�j5�nۊݺ�:ҝ���1f��y�l�i80ԫW��O>��/��Lꐄ�cǂ�(1���N�#:&f�
�y*�G��¦;�-Y��������λ����(�	N����h׾ݘO?�$%'�0���:Y�6�6m�ʔ���#���5*�M^n6����\s"��Q����{���K���@��0�=�Q��o��}�'�?�fM��;�"�`ŀN�.��b\{��6�#""|Wf��Ȫ/���K����^�jӎ.�bي�1b$��މ��\�����g��w�;��>�Y'>�G<"�`ƀN^����۴9�����U��Uv[�n����t@�$������ѣ�d�b�	�JtTTr��-�L�655/;DD�:y����`r�ڴi�Ff�*;ͫ��b�e8���Q���㭉1��o`5���W��k�.���� �n��O?"�`ǀN^}�~.����j���s�yyQ��q8�p�"���"*22��g��oLx��ٰ*�׊��ѭG��Np�����޻o���:`@'��M�ݺ�@TT�&e~^nS�v�U+Wb_J
Z4k�`�i75r����`��y���ϛ�����C��޻Љ��`@'��z�\vŕ��Ď�QQ۳27-���m۶bÆ�A�u��~w��b�vs�ݞݰA��+W,[8��G�Գ;n��jU��S߾}p�ק�<{�Z〭�%�:tK�.����`$����˒�����|�)�ߓ���mxi� "�N�ɧ����
���e�Ͷ��뻗�t`ѢE��ɑ�AՎ.'+��'�h7���]ٮ}����-c��� "���ɧ_�͚�D�:�W���g��^�j;iG߻oZ�h�`�״����p���n7���hܴ�����)_}��K�aԨ "�n�ɧ��.B�=l˚ի����Xt��۱~���	��SRS1z��^Ǜ6�,����\�պ�k0�|���K "��Щ\	uиq�ݪ�%=-�M�-����y��y�5�fϓv�I����v��:uz��/�ʱ���)�����b@�ru��I��9�U�a�Q�c�t`������Flt�1oG�v�7&L���[��#���7o�r�/?��y���ؽsN?�tUW�T.w�8�{�^�򚣠� �j�U+Wa�޽hӪ��x�#Gc��vsy6���s�͜�����O��3O���:c@�r͚5]��@|B����������e���ؾ�֭?f��<�`�E���_{�����/���w'OQuǀN�:��q�7�t:��/]�+++�n٭����v��:��(���y�EtL̎�mڌ�����0 ��Qv;"����_�z����/��?x�`�mLӡ�S���BlL�QoG�����7����`n���7i������3#����`ND!���Ҹi�rӍ��:���l��]y�e���ػwڴnu��MB�Ju\�j߻w,�����P��'�<��AC�1۶m��oL Q�`@'�<��Ø��iG_�J�9y+�Ihݹs'�o�p��������`���n��]�v�g�������q��_3�QHa@'�HǸ�I���Y����J,�v�e˖��AgU�9I0�/(��＋iS�I�?����#�7i����[2���ѳ[Q#��ÀN~��q=��t"۵�߅�2�3,�V3��ѳ��sƣ�4�g���k��΄U����s/�`J��]�v�Z<x߽ "
5���m����n94��S��`5��X�z��KA�U3�g��u6�y�w��˪vUX��]��Ν;��釙Y���� "
E����Cҹ�ٳW��av�� ?�2��x�M7VY@��JO�ر�������n�ڢeˑsf��)�a��_����Q(b@'�=8t(>��+ԩS{UDDxFA~^�	f��Ұt�2�y��*9��~�?|���0M'���e6���Mz��W�r�x���0⹧AD���o���Z�i���M��ѻ�23�Xm�׽*�G����ܹxy����̀uU���s���Mxz�3�5�[��ND!���ֿ�?^Ƥ����/������m�5�Wc_J
Z6o��K0߲u+F��m[7���m�ڷ����{�r���_���?Q(c@�
9����1))�s�n+m6���Hޖ�M�6,�K0����K/��彩�-�����4m�t��?��9���дi\q� "
u�T!��ɨ];			K#""rsrr"�n�jG_�l�vj@��0M|��g���>���U��a��~�ĩ���K/3���1�Y��Q���N2��3q�"22r}dT�����&V������%K�������J������k>^�"2��[���ۻ��*�<��?�����n4$kBGMk׭�bv�r�s'k7��f�v�Y�j^Rlk�Uh3#l[��dE!0�&"��*'8��e7��s�[�<|?3g8����w��9���L����ܶ�3� ���~�>*J���k������%��8m�F�Y�Dz򃴘מ���5k��\���G�|}[Ǎ�� ���T�|~�3y��' ���~�6�f��ҥm�3�t��_`�Kjj���ٳ
����Z:;e}F��������zWxDĎ�~����
� ?_�n� �pB��oK�zJ[`ƞp�m%��e����A�%-�-RRR"���;�jQ��y_v��]v�����	:���cGW@@���1��v:��Ç%.>ABCCK||}�m6k�����V)*:!]6�x�}:��W���Xa��MY+��f�����	�����Z�N��M*{��:�m������gŠ7T;v��J{{���_�|%M�&�w����74HRR��*+�^Q���ᆌ=|��W^����አc@�B�d��Sr?ʭ���0�Ӹ��*����	z_h1���ƍ�$���<��
�?w�?����/�k� W29�$��ϲ.%��*�~���p3J�su^ZZ*�Ϝ��s�ݷW�l�"6�U<͛�Un���o�ަ��RXX(��� �pE�1 ?��DG��M�'����X-���q6[�?^$֧�b4��禥�Dq�$'�H���t�����=>�Ճ���; �.\���x�ጠc@���f�~��������k�X:�=]Mk����-�q];��,)�k�d�	����N'QQQ{�WO�?c��v����+ �;��������L1u�
�k/{�$?w��������&[�n�?�#�}��Z!�!E3�e���hjn�m��  A� ����c�>bޙ�uZ���{ڨ���(��e2c�t���ҝ��'37HW�7ڢ�r�K�Z~:yrʮ���t�3R[^..  A� DDE�,0��_�Sl��~�����(/���EEb�Q����{W���%yM����Iϭv7��Fo׍��;�צ~x�;��Ȋ�� �_6w�,���Hxxx�ȑ#-�W�~�o�����XZ��亠����F6��Jj�:���/�Ӽ���ZdT�;�ߙ�>����%9�� �w:L�"uz\����-��dn�����R[S��o����)ٻ����i��%A����3��^{�g5���*� �C�1`�G����>Ѿ^��Ω����t��_� {��S�Iz}O���]��.�X����s����s�bc7�d��ߕ�P�1���y� ��:eF|��
h	)3��6���8m]��۷K��Y2g�,�8wN��$u_�WK/��i���_�Т7W�|�.�,~H  �"���ks��y��t����ߔNj��%=-]���$c}�=rD<=��]�GFF��=gv�ƍ�N����
 �cP^߲E��#gΜ)�;엺�����򤪲J*����Ԗ�u?o8j��֙�fnX���g�!�>yR  �t��%�n�Nʻ�|\z��t~�)�'��MR�e���i�L�]���훶lq���ɯ�<)  �:�d2ɒ����������ں��tz�~���w'L�X}Ͻ��ݺu���ݻD�d;A��tZ��J�:m��/>q����ā��%�GZܽ s�����j��u�̝@t�'��˧G���;�x�iʦ���X�V����`0J\|\ުU�v,8䊈���� �aC��?��{\Ǝ���?���b}�.�K��`4��W�Ǜ��j����pF�1$��^��:f츎�G������q���>��K:�n[xT��i�ؤ���[� �Cf�Ν��ޮm�r�������T����C�i�+��<�����-�  ����2˖,��/���s�J�ط���w���-���*<!!��]wߕ|������� }G�1���ِ������l�X��m�I=��������3>m�^9��ŕ���*/���  ���cH͙3Gv��-oeeɁ��"_�$�ݑ�]�Qn���z�;f�y��g�9��ӈ9 Aǐ[�x��d2���D����t:&8�UN���|�����`4�1��Eǋ���ʤ��V  C��8UZ*:�QBCB�'LL375�X::��lA:�����'wtp��u��wZ,�z�j1M�$ ��!���86ih��^��������dn�:V: `�:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
�O��Ր���    IEND�B`�PK
     �k�[��EM  M  /   images/d3694a2e-5bba-40c3-8069-8db85c4c9209.png�PNG

   IHDR   d   d   p�T  TiCCPICC Profile  x�c``RI,(�aa``��+)
rwR���R`����b
����>@%0|����/��:%5�I�^��b��Ջ�D������d ��S��JS�l����):
Ȟb�C�@�$�XMH�3�}�VH�H�����IBOGbC�n��ₜ�J� c���Ԋ�_PY���Q���Tϼd=#CsP�CT�%���X�}�����ߍ�������k'BLÂ�A�����΂ĢD�33��10|Z����� |�'�8��,������z����j��N��������.j���p  !e�2���   	pHYs  %  %IR$�   xeXIfII*            (           J       R   i�    Z       %     %      �    o  �           a���  �zTXtRaw profile type icc  x��S[n�0��)z^�8~$R��b;^eW�J�ё"�@`H�n-|DI�D��@ȴ�v=L�"�	�s,`�ۮ��z����"H����pz����3�ͬ,9&�h'�tN9#���(���d>CQ�h�|q�k��R�R����mOi�q�6�Z�ܶ=���C�>hrK$>���U`�͚t3�s;����%�S�T�c��\���~�y§b�_"%�G"a=}J�H����|)�Ni����2��yl�c���r�E��|�7$��8��s���.PJ����
��wq�8��P'��j����[ܞ�c2����g�+��|����RM�=�c2gҥl��ϞauTh���҈�\�z���줡㜥   %tEXtdate:create 2020-01-31T21:31:09+00:00��y{   %tEXtdate:modify 2020-01-31T21:31:00+00:00	�   tEXtexif:ExifOffset 90Y�ޛ   tEXtexif:PixelXDimension 1391c�   tEXtexif:PixelYDimension 800�요   (tEXticc:copyright Copyright Apple Inc., 2017���   tEXticc:description Display P3�y��  cIDATx��]	xLW~��d�(%�J"��}�%(�Z���B��_[y~R�R[u�E[[����J����ҿZ��j��B)��'s��;��Ĉ����>���=��s�s��-�37:�PTB��A%DaP	QTB��A%DaP	QTB��A%DaP	QTB��A%DaP	QTB��AW÷&��z\I���7�)I*�Ev�Z�:d;iJ�3mtRɲ�������V�$IY6��"a[�d��$}/����~�l���99��t.��$u0Z��d�M��(��5D��a�}0�*�
��?���h��dY~�`ȫq+��L��yY���@���[���������ƍ����0��`�Aк�C��"�|<B&�������r����t�PQ:�;w'N�{˧����a)y���3�t>���ʂ
E@fB\yyP� �f�3b�1�(p�3!�<ÃY=��䫄(�d���?0��&1A3vH�JIi�	�YCd��c,�p?��0���g�Ж���lqtws���%b�G��ɒ�2d'jaxR�v�Zl߈s��S�����_C���2Js;�i���8�f�ɒM>�Q.]�����С�x�g/�5J<����зO̚=�g����f6.:6lX�t]������B��5�D��;ѽ[7���s�p�0g�,�n�=_x��(���E��~/���u{���F�m�6�2�h��!����v����;����dX�i5�7�}�����ٿ�2~޳?��#n������1p�@xV�$��u˖�Ѳe��H�zi��|��u��,�Ν'�����ԩ3�/�5PP��7o���,�_���C�޽ѵK���ǚ5k�t�:>�,^|q 4�XȺ����7!&&�+{�_�~��d��ǎ	SԥkW�o؀������A��n��B�p2�7n����Na��>$3��ARLN�G��&����~�� �����QQ��wq�������Тe+xU�ºu_ lQ������͐�լ�K�.����ԙK�.��9����(�QN4|���X�p&M|�����5�OLLDu��x�"�.Y�9o��&�l7ww7�b�rD�c�)��?��޽E��jO����[���a�0�?B��ۿr6n����o�Y�}��E�E�:uh@lAZZ*�i`5]�ر�u�9Ǻ��<s�4�V���ի۽��1�Q�n�:AƢ����D�?O�F�g:b����a� i4puuÑ�#������W��u� ̜�iL8^<H�Ȏ��ʕ+Bui������®�v�u�zS����u>l�ФΝ�P�U�@.��+��������^M�5c�L�L��S��nW",�Y��e��'""#�|���'B�B�FMТœ8���	�R��ӓC��w��t�b�_G�R׿ƛG߭~=L�6U��?���קў��ݻ[��Z���\�rLd0�q�	��o@Ey.D<kI��
2^U��~�zB�!C^65V�E�6m�W���$!-^�j� ��溃��������͂�٤������m׮j׮����{��l"��e����G�fg�AQ�%{ΫbM�6��F�흚6m"�.\@�ƍD���]P��	��g�ΕG���e?h�V��\��ӊ�����ٳq"m���`1i.�[8c:fd��Y����<P��6���׻�2�sq�{dDG2kd'j	h�͛��)2;U�jW��%�=z|j���)�b~b����!JcӁ�L��+$3�i��ߪ[�Fc�8����2�F����~~���dG��?��%\�9���ɡ���3lw[wGDD���Ç�6�V�Z8AQ?��6U_"���YԢq�0��$��_M�i������W[P��@�nns+�F*Z��@'����!����ǤI��`�<a�CI�>��p������<*T�[�Cɩ�1K�,>�>}�/�h�M�vhD�*��89�-�aq�֭�M0m�t�jQt������5k?C��M�ۻ�Mk5���Z�e����ZSVY'�����L���������'����F����g(4�Ŷ��P�^G�>|<(��p������_�R�VUDK</`9rr��WhI�6��E^��9��~��΁�ʧ(��K�c��K�^���}Ѭis<���b�s���J�efp �e
���,���5��<�5o۶oD��h���%.�sab��F��%a�ȑ4I܍��u�Ȗ-�!00�==̤?�9@���������A��"���K�T����J��2
�������r�̋h���C�Шn+���\�t	�i~`�'t�dA�����Ӄ|�'���GEDCQ��z�5{zP�gA`�@��?�h����\�h*��5���]�r^^^pbb(��1��[ޒbo�ػ^8�s4�叽|�4�@����4}�#0(h�my
?A�#����Mg�<��7��?�il���_ �2Eto�����"����j�37-N^��4g��)�8����&��'�*JBCLQ�JH�C���=d��,���}X5D�2`�����0��g窆(&Q#,���!�.o���e�TF��[���9ʲIQ�[�<l�M�V��|/="D�xOR���vG�_G�3˚��7��aj�gE��s�6��ˋk�Q'I����܊�GBEiB���j���QCG�h4Z�D�$ݢY�-R��By%�V+i�T���I|3����4����ĉؙ}���2r����)���Om�fk\]�zH�|�R�iO�l�Mۗ�I6_dْϜf4G��Fk-匷�ݥe�k�\𛍶���V���_�3���X:�-�b(ڴ#ݾ���KĤ����h$�v!VI~}��+s�^����xg��p�h4"�E@�Ӈ$^N������1���	�����ǁ=j��������o��qbZW�?��i�1��wI�t�G��v��e��^3�x޹���k+�t�w��`-;q<3��rJ�r�##���Κr$55G��޶;�a�±c_�ٿΜ�V�{J9�Ԕd��=�(B���}�\�.1�7����׭w�^v�.\�[��"{x<����̣������{�"o���]�|ҵ�"#��[v��n�ٻoޚ>�Mۢ�̛;[�A���(Ks�#�����@�V�s��I������׸��������gn�fV��8\��@�*e	%F��#�n�����8v� �2�Ǎƙ3�2+yV{<6���ܜ����#d9�¡��ȏ ""�z�ז-_�M���^nzjJ�QNk��i�܇��#��~_�Z(_��?���&��2�G9��ɡ�=�gge|�yx�fY$�Q�/R~�'������ll���<����� ~�N�z�����t
s�PVQ��<^�q�s��mOrrJ@�=�t-���K		粲24x6�;�;�%JHJJ
*�|D��-KKMN!p5�olI�x��ݺ�Ge�F��kǏ�H�"A�ռ!i\�xzz�/_�<�R�u�7�u�����U�F��K0��N�rx����̬L�(B���^b���x:y9��}���E������k��%u����QTB��A%DaP	QTB��A%DaP	QTB��A%DaP	QTB��A%DaP	QTB����Blg���    IEND�B`�PK 
     �k�[�O�k�  k�                   cirkitFile.jsonPK 
     �k�[                        ��  jsons/PK 
     �k�[ċ�C+  +               ��  jsons/user_defined.jsonPK 
     �k�[                        �  images/PK 
     �k�[����^� ^� /             '�  images/67df6019-bb76-4308-bacd-6454b246d44a.pngPK 
     �k�[����  �  /             ҟ images/7de8bea6-aec6-4ad5-83ac-8e47725efc1f.pngPK 
     �k�[�I��t� t� /             � images/89718c7b-e32a-4492-aa2b-d7960b76d502.pngPK 
     �k�[�+�sz;  z;  /             �� images/8883793e-4c9f-4ae6-b420-3a6e91b2597d.pngPK 
     �k�[t���?  �?  /             w� images/e2e2c934-b375-45fc-834c-534243cbf361.pngPK 
     �k�[e���  �  /             G" images/6c1978d3-8c4d-4ea9-a1ba-37ab4b096c5d.pngPK 
     �k�[�{�, �, /             c) images/f87b1235-301d-4eff-8a86-0c2fbb955692.pngPK 
     �k�[�ޗԅ  �  /             gV images/2832311d-4ed1-4369-9d2b-9063d9d0cda0.pngPK 
     �k�[�c��f  �f  /             9g images/c88b2895-5e8b-4a57-9f9a-b80dd50058b1.pngPK 
     �k�[��EM  M  /             g� images/d3694a2e-5bba-40c3-8069-8db85c4c9209.pngPK      �  �   