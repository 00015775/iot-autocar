PK
     )u�[�G79�  9�     cirkitFile.json{"raven_core_version":15,"hardware_version":0,"pin_to_graph":{"pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_0_0":[],"pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_1_0":["pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_18"],"pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_0_1":[],"pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_1_1":[],"pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_0_2":[],"pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_1_2":[],"pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_0_3":[],"pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_1_3":[],"pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_0_4":[],"pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_1_4":[],"pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_0_5":[],"pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_1_5":["pin-type-component_b75c9246-bd39-4180-925a-8f93a01a1635_2"],"pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_0_6":[],"pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_1_6":[],"pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_0_7":[],"pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_1_7":[],"pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_0_8":[],"pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_1_8":[],"pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_0_9":[],"pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_1_9":[],"pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_0_10":[],"pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_1_10":["pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_1_16"],"pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_0_11":[],"pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_1_11":[],"pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_0_12":[],"pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_1_12":["pin-type-component_b75c9246-bd39-4180-925a-8f93a01a1635_1","pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_22"],"pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_0_13":[],"pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_1_13":[],"pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_0_14":[],"pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_1_14":["pin-type-component_7ccd86c6-4309-4eb1-9259-cfbd7ebab56f_2","pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_17"],"pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_0_15":[],"pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_1_15":["pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_39","pin-type-component_7ccd86c6-4309-4eb1-9259-cfbd7ebab56f_0","pin-type-component_b75c9246-bd39-4180-925a-8f93a01a1635_0"],"pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_0_16":[],"pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_1_16":["pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_4","pin-type-component_7ccd86c6-4309-4eb1-9259-cfbd7ebab56f_1","pin-type-component_b75c9246-bd39-4180-925a-8f93a01a1635_3","pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_1_10"],"pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_0":[],"pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_1":[],"pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_2":[],"pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_3":[],"pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_4":["pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_1_16"],"pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_5":[],"pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_6":[],"pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_7":[],"pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_8":[],"pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_10":[],"pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_11":[],"pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_12":[],"pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_13":[],"pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_14":[],"pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_16":[],"pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_18":["pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_1_0"],"pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_19":[],"pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_20":[],"pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_21":[],"pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_22":["pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_1_12"],"pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_23":[],"pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_24":[],"pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_25":[],"pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_27":[],"pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_28":[],"pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_29":[],"pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_30":[],"pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_31":[],"pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_32":[],"pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_33":[],"pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_34":[],"pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_35":[],"pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_36":[],"pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_37":[],"pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_38":[],"pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_39":["pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_1_15"],"pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_40":[],"pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_41":[],"pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_15":[],"pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_17":["pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_1_14"],"pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_9":[],"pin-type-component_7ccd86c6-4309-4eb1-9259-cfbd7ebab56f_0":["pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_1_15"],"pin-type-component_7ccd86c6-4309-4eb1-9259-cfbd7ebab56f_1":["pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_1_16"],"pin-type-component_7ccd86c6-4309-4eb1-9259-cfbd7ebab56f_2":["pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_1_14"],"pin-type-component_b75c9246-bd39-4180-925a-8f93a01a1635_0":["pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_1_15"],"pin-type-component_b75c9246-bd39-4180-925a-8f93a01a1635_1":["pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_1_12"],"pin-type-component_b75c9246-bd39-4180-925a-8f93a01a1635_2":["pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_1_5"],"pin-type-component_b75c9246-bd39-4180-925a-8f93a01a1635_3":["pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_1_16"],"pin-type-component_edfd1f52-be35-43c8-85fc-6e1e03d0b2cb_0":[],"pin-type-component_edfd1f52-be35-43c8-85fc-6e1e03d0b2cb_1":[],"pin-type-component_5b6c3c0b-79c1-4551-982f-7c6e68ecec3e_0":[],"pin-type-component_5b6c3c0b-79c1-4551-982f-7c6e68ecec3e_1":[]},"pin_to_color":{"pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_0_0":"#000000","pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_1_0":"#00f900","pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_0_1":"#000000","pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_1_1":"#000000","pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_0_2":"#000000","pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_1_2":"#000000","pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_0_3":"#000000","pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_1_3":"#000000","pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_0_4":"#000000","pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_1_4":"#000000","pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_0_5":"#000000","pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_1_5":"#0056d6","pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_0_6":"#000000","pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_1_6":"#000000","pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_0_7":"#000000","pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_1_7":"#000000","pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_0_8":"#000000","pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_1_8":"#000000","pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_0_9":"#000000","pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_1_9":"#000000","pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_0_10":"#000000","pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_1_10":"#000000","pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_0_11":"#000000","pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_1_11":"#000000","pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_0_12":"#000000","pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_1_12":"#be38f3","pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_0_13":"#000000","pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_1_13":"#000000","pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_0_14":"#000000","pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_1_14":"#ff9300","pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_0_15":"#000000","pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_1_15":"#ff2600","pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_0_16":"#000000","pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_1_16":"#000000","pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_0":"#000000","pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_1":"#000000","pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_2":"#000000","pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_3":"#000000","pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_4":"#000000","pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_5":"#000000","pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_6":"#000000","pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_7":"#000000","pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_8":"#000000","pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_10":"#000000","pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_11":"#000000","pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_12":"#000000","pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_13":"#000000","pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_14":"#000000","pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_16":"#000000","pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_18":"#00f900","pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_19":"#000000","pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_20":"#000000","pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_21":"#000000","pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_22":"#be38f3","pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_23":"#000000","pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_24":"#000000","pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_25":"#000000","pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_27":"#000000","pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_28":"#000000","pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_29":"#000000","pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_30":"#000000","pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_31":"#000000","pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_32":"#000000","pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_33":"#000000","pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_34":"#000000","pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_35":"#000000","pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_36":"#000000","pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_37":"#000000","pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_38":"#000000","pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_39":"#ff2600","pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_40":"#000000","pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_41":"#000000","pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_15":"#000000","pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_17":"#ff9300","pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_9":"#000000","pin-type-component_7ccd86c6-4309-4eb1-9259-cfbd7ebab56f_0":"#ff2600","pin-type-component_7ccd86c6-4309-4eb1-9259-cfbd7ebab56f_1":"#000000","pin-type-component_7ccd86c6-4309-4eb1-9259-cfbd7ebab56f_2":"#ff9300","pin-type-component_b75c9246-bd39-4180-925a-8f93a01a1635_0":"#ff2600","pin-type-component_b75c9246-bd39-4180-925a-8f93a01a1635_1":"#be38f3","pin-type-component_b75c9246-bd39-4180-925a-8f93a01a1635_2":"#0056d6","pin-type-component_b75c9246-bd39-4180-925a-8f93a01a1635_3":"#000000","pin-type-component_edfd1f52-be35-43c8-85fc-6e1e03d0b2cb_0":"#000000","pin-type-component_edfd1f52-be35-43c8-85fc-6e1e03d0b2cb_1":"#000000","pin-type-component_5b6c3c0b-79c1-4551-982f-7c6e68ecec3e_0":"#000000","pin-type-component_5b6c3c0b-79c1-4551-982f-7c6e68ecec3e_1":"#000000"},"pin_to_state":{"pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_0_0":"neutral","pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_1_0":"neutral","pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_0_1":"neutral","pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_1_1":"neutral","pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_0_2":"neutral","pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_1_2":"neutral","pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_0_3":"neutral","pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_1_3":"neutral","pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_0_4":"neutral","pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_1_4":"neutral","pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_0_5":"neutral","pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_1_5":"neutral","pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_0_6":"neutral","pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_1_6":"neutral","pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_0_7":"neutral","pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_1_7":"neutral","pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_0_8":"neutral","pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_1_8":"neutral","pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_0_9":"neutral","pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_1_9":"neutral","pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_0_10":"neutral","pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_1_10":"neutral","pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_0_11":"neutral","pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_1_11":"neutral","pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_0_12":"neutral","pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_1_12":"neutral","pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_0_13":"neutral","pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_1_13":"neutral","pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_0_14":"neutral","pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_1_14":"neutral","pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_0_15":"neutral","pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_1_15":"neutral","pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_0_16":"neutral","pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_1_16":"neutral","pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_0":"neutral","pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_1":"neutral","pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_2":"neutral","pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_3":"neutral","pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_4":"neutral","pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_5":"neutral","pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_6":"neutral","pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_7":"neutral","pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_8":"neutral","pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_10":"neutral","pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_11":"neutral","pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_12":"neutral","pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_13":"neutral","pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_14":"neutral","pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_16":"neutral","pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_18":"neutral","pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_19":"neutral","pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_20":"neutral","pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_21":"neutral","pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_22":"neutral","pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_23":"neutral","pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_24":"neutral","pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_25":"neutral","pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_27":"neutral","pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_28":"neutral","pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_29":"neutral","pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_30":"neutral","pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_31":"neutral","pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_32":"neutral","pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_33":"neutral","pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_34":"neutral","pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_35":"neutral","pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_36":"neutral","pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_37":"neutral","pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_38":"neutral","pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_39":"neutral","pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_40":"neutral","pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_41":"neutral","pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_15":"neutral","pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_17":"neutral","pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_9":"neutral","pin-type-component_7ccd86c6-4309-4eb1-9259-cfbd7ebab56f_0":"neutral","pin-type-component_7ccd86c6-4309-4eb1-9259-cfbd7ebab56f_1":"neutral","pin-type-component_7ccd86c6-4309-4eb1-9259-cfbd7ebab56f_2":"neutral","pin-type-component_b75c9246-bd39-4180-925a-8f93a01a1635_0":"neutral","pin-type-component_b75c9246-bd39-4180-925a-8f93a01a1635_1":"neutral","pin-type-component_b75c9246-bd39-4180-925a-8f93a01a1635_2":"neutral","pin-type-component_b75c9246-bd39-4180-925a-8f93a01a1635_3":"neutral","pin-type-component_edfd1f52-be35-43c8-85fc-6e1e03d0b2cb_0":"neutral","pin-type-component_edfd1f52-be35-43c8-85fc-6e1e03d0b2cb_1":"neutral","pin-type-component_5b6c3c0b-79c1-4551-982f-7c6e68ecec3e_0":"neutral","pin-type-component_5b6c3c0b-79c1-4551-982f-7c6e68ecec3e_1":"neutral"},"next_color_idx":11,"wires_placed_in_order":[["pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_39","pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_1_16"],["pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_4","pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_1_15"],["pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_1_16","pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_1_14"],["pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_1_11","pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_39"],["pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_1_16","pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_4"],["pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_1_15","pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_39"],["pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_1_16","pin-type-component_7ccd86c6-4309-4eb1-9259-cfbd7ebab56f_1"],["pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_1_15","pin-type-component_7ccd86c6-4309-4eb1-9259-cfbd7ebab56f_0"],["pin-type-component_7ccd86c6-4309-4eb1-9259-cfbd7ebab56f_2","pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_1_14"],["pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_1_14","pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_17"],["pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_1_15","pin-type-component_b75c9246-bd39-4180-925a-8f93a01a1635_0"],["pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_1_16","pin-type-component_b75c9246-bd39-4180-925a-8f93a01a1635_3"],["pin-type-component_b75c9246-bd39-4180-925a-8f93a01a1635_1","pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_1_12"],["pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_1_12","pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_22"],["pin-type-component_b75c9246-bd39-4180-925a-8f93a01a1635_2","pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_1_7"],["pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_1_4","pin-type-component_b75c9246-bd39-4180-925a-8f93a01a1635_2"],["pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_1_5","pin-type-component_b75c9246-bd39-4180-925a-8f93a01a1635_2"],["pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_1_0","pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_18"],["pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_1_16","pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_1_10"]],"wires_removed_and_placed_in_order":[[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[["pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_39","pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_1_16"]]],[[],[["pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_4","pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_1_15"]]],[[],[["pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_1_16","pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_1_14"]]],[[["pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_1_14","pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_1_16"]],[]],[[["pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_1_16","pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_39"]],[]],[[],[["pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_1_11","pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_39"]]],[[["pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_1_15","pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_4"]],[]],[[],[["pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_1_16","pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_4"]]],[[["pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_1_11","pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_39"]],[]],[[],[["pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_1_15","pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_39"]]],[[],[["pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_1_16","pin-type-component_7ccd86c6-4309-4eb1-9259-cfbd7ebab56f_1"]]],[[],[["pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_1_15","pin-type-component_7ccd86c6-4309-4eb1-9259-cfbd7ebab56f_0"]]],[[],[["pin-type-component_7ccd86c6-4309-4eb1-9259-cfbd7ebab56f_2","pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_1_14"]]],[[],[["pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_1_14","pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_17"]]],[[],[["pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_1_15","pin-type-component_b75c9246-bd39-4180-925a-8f93a01a1635_0"]]],[[],[["pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_1_16","pin-type-component_b75c9246-bd39-4180-925a-8f93a01a1635_3"]]],[[],[["pin-type-component_b75c9246-bd39-4180-925a-8f93a01a1635_1","pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_1_12"]]],[[],[["pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_1_12","pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_22"]]],[[],[["pin-type-component_b75c9246-bd39-4180-925a-8f93a01a1635_2","pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_1_7"]]],[[],[]],[[],[]],[[],[]],[[],[]],[[["pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_1_7","pin-type-component_b75c9246-bd39-4180-925a-8f93a01a1635_2"]],[]],[[],[["pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_1_4","pin-type-component_b75c9246-bd39-4180-925a-8f93a01a1635_2"]]],[[["pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_1_4","pin-type-component_b75c9246-bd39-4180-925a-8f93a01a1635_2"]],[]],[[],[["pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_1_5","pin-type-component_b75c9246-bd39-4180-925a-8f93a01a1635_2"]]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[["pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_1_0","pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_18"]]],[[],[["pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_1_16","pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_1_10"]]]],"arduino_state":"arduino_off","pin_to_uid":{"pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_0_0":"_","pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_1_0":"0000000000000005","pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_0_1":"_","pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_1_1":"_","pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_0_2":"_","pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_1_2":"_","pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_0_3":"_","pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_1_3":"_","pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_0_4":"_","pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_1_4":"_","pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_0_5":"_","pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_1_5":"0000000000000004","pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_0_6":"_","pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_1_6":"_","pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_0_7":"_","pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_1_7":"_","pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_0_8":"_","pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_1_8":"_","pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_0_9":"_","pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_1_9":"_","pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_0_10":"_","pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_1_10":"0000000000000001","pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_0_11":"_","pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_1_11":"_","pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_0_12":"_","pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_1_12":"0000000000000003","pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_0_13":"_","pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_1_13":"_","pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_0_14":"_","pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_1_14":"0000000000000002","pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_0_15":"_","pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_1_15":"0000000000000000","pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_0_16":"_","pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_1_16":"0000000000000001","pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_0":"_","pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_1":"_","pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_2":"_","pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_3":"_","pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_4":"0000000000000001","pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_5":"_","pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_6":"_","pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_7":"_","pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_8":"_","pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_10":"_","pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_11":"_","pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_12":"_","pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_13":"_","pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_14":"_","pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_16":"_","pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_18":"0000000000000005","pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_19":"_","pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_20":"_","pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_21":"_","pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_22":"0000000000000003","pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_23":"_","pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_24":"_","pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_25":"_","pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_27":"_","pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_28":"_","pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_29":"_","pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_30":"_","pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_31":"_","pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_32":"_","pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_33":"_","pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_34":"_","pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_35":"_","pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_36":"_","pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_37":"_","pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_38":"_","pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_39":"0000000000000000","pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_40":"_","pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_41":"_","pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_15":"_","pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_17":"0000000000000002","pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_9":"_","pin-type-component_7ccd86c6-4309-4eb1-9259-cfbd7ebab56f_0":"0000000000000000","pin-type-component_7ccd86c6-4309-4eb1-9259-cfbd7ebab56f_1":"0000000000000001","pin-type-component_7ccd86c6-4309-4eb1-9259-cfbd7ebab56f_2":"0000000000000002","pin-type-component_b75c9246-bd39-4180-925a-8f93a01a1635_0":"0000000000000000","pin-type-component_b75c9246-bd39-4180-925a-8f93a01a1635_1":"0000000000000003","pin-type-component_b75c9246-bd39-4180-925a-8f93a01a1635_2":"0000000000000004","pin-type-component_b75c9246-bd39-4180-925a-8f93a01a1635_3":"0000000000000001","pin-type-component_edfd1f52-be35-43c8-85fc-6e1e03d0b2cb_0":"_","pin-type-component_edfd1f52-be35-43c8-85fc-6e1e03d0b2cb_1":"_","pin-type-component_5b6c3c0b-79c1-4551-982f-7c6e68ecec3e_0":"_","pin-type-component_5b6c3c0b-79c1-4551-982f-7c6e68ecec3e_1":"_"},"component_id_to_pins":{"2a286633-8d58-4d0e-a66b-e5c265b1c5ff":["0","1","2","3","4","5","6","7","8","10","11","12","13","14","16","18","19","20","21","22","23","24","25","27","28","29","30","31","32","33","34","35","36","37","38","39","40","41","15","17","9"],"7ccd86c6-4309-4eb1-9259-cfbd7ebab56f":["0","1","2"],"b75c9246-bd39-4180-925a-8f93a01a1635":["0","1","2","3"],"edfd1f52-be35-43c8-85fc-6e1e03d0b2cb":["0","1"],"5b6c3c0b-79c1-4551-982f-7c6e68ecec3e":["0","1"],"5b7dade3-fdd8-4f95-986c-ffa4274ae6f5":[]},"uid_to_net":{"_":[],"0000000000000001":["pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_1_16","pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_4","pin-type-component_7ccd86c6-4309-4eb1-9259-cfbd7ebab56f_1","pin-type-component_b75c9246-bd39-4180-925a-8f93a01a1635_3","pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_1_10"],"0000000000000000":["pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_1_15","pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_39","pin-type-component_7ccd86c6-4309-4eb1-9259-cfbd7ebab56f_0","pin-type-component_b75c9246-bd39-4180-925a-8f93a01a1635_0"],"0000000000000002":["pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_1_14","pin-type-component_7ccd86c6-4309-4eb1-9259-cfbd7ebab56f_2","pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_17"],"0000000000000003":["pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_1_12","pin-type-component_b75c9246-bd39-4180-925a-8f93a01a1635_1","pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_22"],"0000000000000004":["pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_1_5","pin-type-component_b75c9246-bd39-4180-925a-8f93a01a1635_2"],"0000000000000005":["pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_1_0","pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_18"]},"uid_to_text_label":{"0000000000000001":"Net 1","0000000000000000":"Net 0","0000000000000002":"Net 2","0000000000000003":"Net 3","0000000000000004":"Net 4","0000000000000005":"Net 5"},"all_breadboard_info_list":["d4a0d558-beb3-4ff5-847e-afd45f379ae0_17_2_False_722_243_left"],"breadboard_info_list":["d4a0d558-beb3-4ff5-847e-afd45f379ae0_17_2_False_722_243_left"],"componentsData":[{"compProperties":{"mpn":{"version":2,"id":"mpn","label":"mpn","description":"","units":"","type":"string","value":"RPI3-MODB-16GB-NOOBS","displayFormat":"input","showOnComp":false,"isVisibleToUser":false},"manufacturer":{"version":2,"id":"manufacturer","label":"manufacturer","description":"","units":"","type":"string","value":"Raspberry Pi","displayFormat":"input","showOnComp":false,"isVisibleToUser":false}},"position":[1229.31025,375.44717],"typeId":"9d987227-334c-49a7-9e0b-80422ab638f6","componentVersion":2,"instanceId":"2a286633-8d58-4d0e-a66b-e5c265b1c5ff","orientation":"up","circleData":[[1022.5,230],[1037.5,230],[1052.5,230],[1067.5,230],[1082.5,230],[1097.5,230],[1112.5,230],[1127.5,230],[1142.5,230],[1172.5,230],[1187.5,230],[1202.5,230],[1217.5,230],[1232.5,230],[1262.5,230],[1292.5,230],[1307.5,230],[1307.5,215],[1292.5,215],[1277.5,215],[1262.5,215],[1247.5,215],[1232.5,215],[1202.5,215],[1187.5,215],[1172.5,215],[1157.5,215],[1142.5,215],[1127.5,215],[1112.5,215],[1097.5,215],[1082.5,215],[1067.5,215],[1052.5,215],[1037.5,215],[1022.5,215],[1157.5,230],[1217.5,215],[1247.5,230],[1277.5,230],[1036.6615,531.6770000000005]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[618.1357344999999,634.0469494999999],"typeId":"d41d5606-8708-4dc6-b0f7-7b5da01a1617","componentVersion":1,"instanceId":"7ccd86c6-4309-4eb1-9259-cfbd7ebab56f","orientation":"left","circleData":[[752.5,635],[752.4991315,619.753367],[752.5,652.1525]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"mpn":{"version":2,"id":"mpn","label":"mpn","description":"","units":"","type":"string","value":"SEN-15569","displayFormat":"input","showOnComp":false,"isVisibleToUser":false},"manufacturer":{"version":2,"id":"manufacturer","label":"manufacturer","description":"","units":"","type":"string","value":"SparkFun","displayFormat":"input","showOnComp":false,"isVisibleToUser":false}},"position":[537.0136134999999,-16.50356499999998],"typeId":"f7a95729-a811-496b-83f5-7789de376adf","componentVersion":2,"instanceId":"b75c9246-bd39-4180-925a-8f93a01a1635","orientation":"up","circleData":[[512.5,49.99999999999999],[527.4992245,49.99999999999999],[542.4999985,49.99530950000001],[557.4984445,49.9937495]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"Resistance":{"version":2,"id":"Resistance","label":"Resistance","description":"","units":"Ω","type":"decimal","value":"1000","displayFormat":"input","showOnComp":true,"isVisibleToUser":true},"Tolerance":{"version":2,"id":"Tolerance","label":"Tolerance","description":"","units":"","type":"string","value":"5%","displayFormat":"dropdown","options":[{"label":"0.25%","value":"0.25%"},{"label":"0.1%","value":"0.1%"},{"label":"0.5%","value":"0.5%"},{"label":"1%","value":"1%"},{"label":"2%","value":"2%"},{"label":"5%","value":"5%"},{"label":"10%","value":"10%"}],"showOnComp":false,"isVisibleToUser":true},"Number Of Bands":{"version":2,"id":"Number Of Bands","label":"Number Of Bands","description":"","units":"","type":"string","value":"5","displayFormat":"dropdown","options":[{"label":"4","value":"4"},{"label":"5","value":"5"},{"label":"6","value":"6"}],"showOnComp":false,"isVisibleToUser":true}},"position":[684.1735537190082,335],"typeId":"72c75556-baa3-04e7-55a5-e13f447c8c5a","componentVersion":1,"instanceId":"edfd1f52-be35-43c8-85fc-6e1e03d0b2cb","orientation":"up","circleData":[[647.5,335],[722.5,335]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"Resistance":{"version":2,"id":"Resistance","label":"Resistance","description":"","units":"Ω","type":"decimal","value":"1000","displayFormat":"input","showOnComp":true,"isVisibleToUser":true,"name":"Resistance","unit":"Ω","required":true,"validRange":[0,70000]},"Tolerance":{"version":2,"id":"Tolerance","label":"Tolerance","description":"","units":"","type":"string","value":"5%","displayFormat":"dropdown","options":[{"label":"0.25%","value":"0.25%"},{"label":"0.1%","value":"0.1%"},{"label":"0.5%","value":"0.5%"},{"label":"1%","value":"1%"},{"label":"2%","value":"2%"},{"label":"5%","value":"5%"},{"label":"10%","value":"10%"}],"showOnComp":false,"isVisibleToUser":true,"name":"Tolerance","required":true},"Number Of Bands":{"version":2,"id":"Number Of Bands","label":"Number Of Bands","description":"","units":"","type":"string","value":"5","displayFormat":"dropdown","options":[{"label":"4","value":"4"},{"label":"5","value":"5"},{"label":"6","value":"6"}],"showOnComp":false,"isVisibleToUser":true,"name":"Number Of Bands","required":true}},"position":[760,305],"typeId":"72c75556-baa3-04e7-55a5-e13f447c8c5a","componentVersion":1,"instanceId":"5b6c3c0b-79c1-4551-982f-7c6e68ecec3e","orientation":"up","circleData":[[722.5,305],[797.5,305]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"Comment":{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"Servo SG09 motor:\n  RED - VCC, 5V\n  YELLOW - GPIO19; \n   PWN enabled pins (BCM: GPIO12, GPIO13, GPIO18, GPIO19) if available.\n  BROWN - GND\n\nHC-SR04 Ultrasonic sensor pins:\n  VCC - 5V\n  GND - GND\n  TRIG - GPIO16\n  ECHO - GPIO26\n  \n Make sure to use voltage divider with two resistors \n for pin connected to Echo. Otherwise the program \n will not work and Pi can be damaged!\n\n Instead of connecting GND and VCC individually to ultrasonic\n and servo, a single GND/VCC is connected to breadboard\n and from there distributed to ultrasonic and servo motor. ","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"backgroundColor":{"version":2,"id":"backgroundColor","label":"Background Color","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"backgroundOpacity":{"version":2,"id":"backgroundOpacity","label":"Background Opacity","description":"","units":"","type":"decimal","value":"1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"textColor":{"version":2,"id":"textColor","label":"Text Color","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"fontSize":{"version":2,"id":"fontSize","label":"Font Size","description":"","units":"","type":"integer","value":"12","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"font":{"version":2,"id":"font","label":"Font","description":"","units":"","type":"string","value":"Arial","displayFormat":"input","showOnComp":false,"isVisibleToUser":true}},"position":[1193.7483777763432,-66.77272727272734],"typeId":"9a5a4baa-44d4-4aa0-8d82-488487322b20","componentVersion":1,"instanceId":"5b7dade3-fdd8-4f95-986c-ffa4274ae6f5","orientation":"up","circleData":[],"cirkitStudioVersion":"1.3.3"}],"bounds":{"top":"-213.57273","left":"393.85321","width":"1101.67354","height":"904.84073","x":"393.85321","y":"-213.57273"},"cachedBreadboardPrettyViewWires":["{\"color\":\"#000000\",\"startPinId\":\"pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_1_16\",\"endPinId\":\"pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_4\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_d4a0d558-beb3-4ff5-847e-afd45f379ae0_1_16_4\",\"rawEndPinId\":\"pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_4\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"887.5000000000_290.0000000000\\\",\\\"887.5000000000_140.0000000000\\\",\\\"1082.5000000000_140.0000000000\\\",\\\"1082.5000000000_230.0000000000\\\"]}\"}","{\"color\":\"#000000\",\"startPinId\":\"pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_1_16\",\"endPinId\":\"pin-type-component_7ccd86c6-4309-4eb1-9259-cfbd7ebab56f_1\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_d4a0d558-beb3-4ff5-847e-afd45f379ae0_1_16_3\",\"rawEndPinId\":\"pin-type-component_7ccd86c6-4309-4eb1-9259-cfbd7ebab56f_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"887.5000000000_305.0000000000\\\",\\\"925.0000000000_305.0000000000\\\",\\\"925.0000000000_620.0000000000\\\",\\\"752.4991315000_620.0000000000\\\",\\\"752.4991315000_619.7533670000\\\"]}\"}","{\"color\":\"#000000\",\"startPinId\":\"pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_1_16\",\"endPinId\":\"pin-type-component_b75c9246-bd39-4180-925a-8f93a01a1635_3\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_d4a0d558-beb3-4ff5-847e-afd45f379ae0_1_16_1\",\"rawEndPinId\":\"pin-type-component_b75c9246-bd39-4180-925a-8f93a01a1635_3\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"887.5000000000_335.0000000000\\\",\\\"962.5000000000_335.0000000000\\\",\\\"962.5000000000_65.0000000000\\\",\\\"557.4984445000_65.0000000000\\\",\\\"557.4984445000_49.9937495000\\\"]}\"}","{\"color\":\"#000000\",\"startPinId\":\"pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_1_10\",\"endPinId\":\"pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_1_16\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_d4a0d558-beb3-4ff5-847e-afd45f379ae0_1_10_4\",\"rawEndPinId\":\"pin-type-breadboard-sub-pin_d4a0d558-beb3-4ff5-847e-afd45f379ae0_1_16_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"797.5000000000_290.0000000000\\\",\\\"797.5000000000_275.0000000000\\\",\\\"812.5000000000_275.0000000000\\\",\\\"812.5000000000_387.5000000000\\\",\\\"887.5000000000_387.5000000000\\\",\\\"887.5000000000_350.0000000000\\\"]}\"}","{\"color\":\"#ff2600\",\"startPinId\":\"pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_1_15\",\"endPinId\":\"pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_39\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_d4a0d558-beb3-4ff5-847e-afd45f379ae0_1_15_4\",\"rawEndPinId\":\"pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_39\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"872.5000000000_290.0000000000\\\",\\\"872.5000000000_125.0000000000\\\",\\\"1022.5000000000_125.0000000000\\\",\\\"1022.5000000000_215.0000000000\\\"]}\"}","{\"color\":\"#ff2600\",\"startPinId\":\"pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_1_15\",\"endPinId\":\"pin-type-component_7ccd86c6-4309-4eb1-9259-cfbd7ebab56f_0\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_d4a0d558-beb3-4ff5-847e-afd45f379ae0_1_15_0\",\"rawEndPinId\":\"pin-type-component_7ccd86c6-4309-4eb1-9259-cfbd7ebab56f_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"872.5000000000_350.0000000000\\\",\\\"872.5000000000_635.0000000000\\\",\\\"752.5000000000_635.0000000000\\\"]}\"}","{\"color\":\"#ff2600\",\"startPinId\":\"pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_1_15\",\"endPinId\":\"pin-type-component_b75c9246-bd39-4180-925a-8f93a01a1635_0\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_d4a0d558-beb3-4ff5-847e-afd45f379ae0_1_15_2\",\"rawEndPinId\":\"pin-type-component_b75c9246-bd39-4180-925a-8f93a01a1635_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"872.5000000000_320.0000000000\\\",\\\"872.5000000000_305.0000000000\\\",\\\"842.5000000000_305.0000000000\\\",\\\"842.5000000000_110.0000000000\\\",\\\"512.5000000000_110.0000000000\\\",\\\"512.5000000000_50.0000000000\\\"]}\"}","{\"color\":\"#ff9300\",\"startPinId\":\"pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_1_14\",\"endPinId\":\"pin-type-component_7ccd86c6-4309-4eb1-9259-cfbd7ebab56f_2\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_d4a0d558-beb3-4ff5-847e-afd45f379ae0_1_14_0\",\"rawEndPinId\":\"pin-type-component_7ccd86c6-4309-4eb1-9259-cfbd7ebab56f_2\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"857.5000000000_350.0000000000\\\",\\\"857.5000000000_652.1525000000\\\",\\\"752.5000000000_652.1525000000\\\"]}\"}","{\"color\":\"#ff9300\",\"startPinId\":\"pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_1_14\",\"endPinId\":\"pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_17\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_d4a0d558-beb3-4ff5-847e-afd45f379ae0_1_14_1\",\"rawEndPinId\":\"pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_17\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"857.5000000000_335.0000000000\\\",\\\"857.5000000000_110.0000000000\\\",\\\"1337.5000000000_110.0000000000\\\",\\\"1337.5000000000_252.5000000000\\\",\\\"1277.5000000000_252.5000000000\\\",\\\"1277.5000000000_230.0000000000\\\"]}\"}","{\"color\":\"#be38f3\",\"startPinId\":\"pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_1_12\",\"endPinId\":\"pin-type-component_b75c9246-bd39-4180-925a-8f93a01a1635_1\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_d4a0d558-beb3-4ff5-847e-afd45f379ae0_1_12_1\",\"rawEndPinId\":\"pin-type-component_b75c9246-bd39-4180-925a-8f93a01a1635_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"827.5000000000_335.0000000000\\\",\\\"827.5000000000_95.0000000000\\\",\\\"527.4992245000_95.0000000000\\\",\\\"527.4992245000_50.0000000000\\\"]}\"}","{\"color\":\"#be38f3\",\"startPinId\":\"pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_1_12\",\"endPinId\":\"pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_22\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_d4a0d558-beb3-4ff5-847e-afd45f379ae0_1_12_0\",\"rawEndPinId\":\"pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_22\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"827.5000000000_350.0000000000\\\",\\\"827.5000000000_372.5000000000\\\",\\\"1375.0000000000_372.5000000000\\\",\\\"1375.0000000000_177.5000000000\\\",\\\"1277.5000000000_177.5000000000\\\",\\\"1277.5000000000_215.0000000000\\\"]}\"}","{\"color\":\"#0056d6\",\"startPinId\":\"pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_1_5\",\"endPinId\":\"pin-type-component_b75c9246-bd39-4180-925a-8f93a01a1635_2\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_d4a0d558-beb3-4ff5-847e-afd45f379ae0_1_5_0\",\"rawEndPinId\":\"pin-type-component_b75c9246-bd39-4180-925a-8f93a01a1635_2\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"722.5000000000_350.0000000000\\\",\\\"722.5000000000_365.0000000000\\\",\\\"542.4999985000_365.0000000000\\\",\\\"542.4999985000_49.9953095000\\\"]}\"}","{\"color\":\"#00f900\",\"startPinId\":\"pin-type-breadboard_d4a0d558-beb3-4ff5-847e-afd45f379ae0_1_0\",\"endPinId\":\"pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_18\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_d4a0d558-beb3-4ff5-847e-afd45f379ae0_1_0_2\",\"rawEndPinId\":\"pin-type-component_2a286633-8d58-4d0e-a66b-e5c265b1c5ff_18\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"647.5000000000_320.0000000000\\\",\\\"602.5000000000_320.0000000000\\\",\\\"602.5000000000_402.5000000000\\\",\\\"1292.5000000000_402.5000000000\\\",\\\"1292.5000000000_230.0000000000\\\"]}\"}"],"projectDescription":""}PK
     )u�[               jsons/PK
     )u�[�fy�(  �(     jsons/user_defined.json{"type":"user_defined","version":"0.0.1","subtypes":[{"subtypeName":"Raspberry Pi 3B","category":["User Defined"],"userDefined":true,"id":"9d987227-334c-49a7-9e0b-80422ab638f6","subtypeDescription":"","subtypePic":"67df6019-bb76-4308-bacd-6454b246d44a.png","pinInfo":{"numDisplayCols":"34.16220","numDisplayRows":"22.82490","pins":[{"uniquePinIdString":"0","positionMil":"329.37500,2110.89280","isAnchorPin":true,"label":"1"},{"uniquePinIdString":"1","positionMil":"429.37500,2110.89280","isAnchorPin":false,"label":"3"},{"uniquePinIdString":"2","positionMil":"529.37500,2110.89280","isAnchorPin":false,"label":"5"},{"uniquePinIdString":"3","positionMil":"629.37500,2110.89280","isAnchorPin":false,"label":"7"},{"uniquePinIdString":"4","positionMil":"729.37500,2110.89280","isAnchorPin":false,"label":"9"},{"uniquePinIdString":"5","positionMil":"829.37500,2110.89280","isAnchorPin":false,"label":"11"},{"uniquePinIdString":"6","positionMil":"929.37500,2110.89280","isAnchorPin":false,"label":"13"},{"uniquePinIdString":"7","positionMil":"1029.37500,2110.89280","isAnchorPin":false,"label":"15"},{"uniquePinIdString":"8","positionMil":"1129.37500,2110.89280","isAnchorPin":false,"label":"17"},{"uniquePinIdString":"10","positionMil":"1329.37500,2110.89280","isAnchorPin":false,"label":"21"},{"uniquePinIdString":"11","positionMil":"1429.37500,2110.89280","isAnchorPin":false,"label":"23"},{"uniquePinIdString":"12","positionMil":"1529.37500,2110.89280","isAnchorPin":false,"label":"25"},{"uniquePinIdString":"13","positionMil":"1629.37500,2110.89280","isAnchorPin":false,"label":"27"},{"uniquePinIdString":"14","positionMil":"1729.37500,2110.89280","isAnchorPin":false,"label":"29"},{"uniquePinIdString":"16","positionMil":"1929.37500,2110.89280","isAnchorPin":false,"label":"33"},{"uniquePinIdString":"18","positionMil":"2129.37500,2110.89280","isAnchorPin":false,"label":"37"},{"uniquePinIdString":"19","positionMil":"2229.37500,2110.89280","isAnchorPin":false,"label":"39"},{"uniquePinIdString":"20","positionMil":"2229.37500,2210.89280","isAnchorPin":false,"label":"40"},{"uniquePinIdString":"21","positionMil":"2129.37500,2210.89280","isAnchorPin":false,"label":"38"},{"uniquePinIdString":"22","positionMil":"2029.37500,2210.89280","isAnchorPin":false,"label":"36"},{"uniquePinIdString":"23","positionMil":"1929.37500,2210.89280","isAnchorPin":false,"label":"34"},{"uniquePinIdString":"24","positionMil":"1829.37500,2210.89280","isAnchorPin":false,"label":"32"},{"uniquePinIdString":"25","positionMil":"1729.37500,2210.89280","isAnchorPin":false,"label":"30"},{"uniquePinIdString":"27","positionMil":"1529.37500,2210.89280","isAnchorPin":false,"label":"26"},{"uniquePinIdString":"28","positionMil":"1429.37500,2210.89280","isAnchorPin":false,"label":"24"},{"uniquePinIdString":"29","positionMil":"1329.37500,2210.89280","isAnchorPin":false,"label":"22"},{"uniquePinIdString":"30","positionMil":"1229.37500,2210.89280","isAnchorPin":false,"label":"20"},{"uniquePinIdString":"31","positionMil":"1129.37500,2210.89280","isAnchorPin":false,"label":"18"},{"uniquePinIdString":"32","positionMil":"1029.37500,2210.89280","isAnchorPin":false,"label":"16"},{"uniquePinIdString":"33","positionMil":"929.37500,2210.89280","isAnchorPin":false,"label":"14"},{"uniquePinIdString":"34","positionMil":"829.37500,2210.89280","isAnchorPin":false,"label":"12"},{"uniquePinIdString":"35","positionMil":"729.37500,2210.89280","isAnchorPin":false,"label":"10"},{"uniquePinIdString":"36","positionMil":"629.37500,2210.89280","isAnchorPin":false,"label":"8"},{"uniquePinIdString":"37","positionMil":"529.37500,2210.89280","isAnchorPin":false,"label":"6"},{"uniquePinIdString":"38","positionMil":"429.37500,2210.89280","isAnchorPin":false,"label":"4"},{"uniquePinIdString":"39","positionMil":"329.37500,2210.89280","isAnchorPin":false,"label":"2(5V)"},{"uniquePinIdString":"40","positionMil":"1229.37500,2110.89280","isAnchorPin":false,"label":"19"},{"uniquePinIdString":"41","positionMil":"1629.37500,2210.89280","isAnchorPin":false,"label":"28"},{"uniquePinIdString":"15","positionMil":"1829.37500,2110.89280","isAnchorPin":false,"label":"31"},{"uniquePinIdString":"17","positionMil":"2029.37500,2110.89280","isAnchorPin":false,"label":"35"},{"uniquePinIdString":"9","positionMil":"423.78500,99.71280","isAnchorPin":false,"label":"Power"}],"pinType":"wired"},"properties":[{"type":"string","name":"mpn","value":"RPI3-MODB-16GB-NOOBS","unit":"","showOnComp":false,"userVisible":false,"required":true},{"type":"string","name":"manufacturer","value":"Raspberry Pi","unit":"","showOnComp":false,"userVisible":false,"required":true}],"iconPic":"7de8bea6-aec6-4ad5-83ac-8e47725efc1f.png","componentVersion":2,"imageLocation":"local_cache","hasComponentImageSvg":false,"componentImageSvgUrl":""},{"subtypeName":"servo motor ","category":["User Defined"],"id":"d41d5606-8708-4dc6-b0f7-7b5da01a1617","componentVersion":1,"userDefined":true,"subtypeDescription":"","subtypePic":"b3e67e62-159a-497d-aba3-70fd70f56319.png","iconPic":"ab942d8a-eab6-45a7-8f5a-30ef729b6f10.png","hasComponentImageSvg":false,"componentImageSvgUrl":"","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"6.29614","numDisplayRows":"19.69562","pins":[{"uniquePinIdString":"0","positionMil":"308.45333,89.01923","isAnchorPin":true,"label":"VCC"},{"uniquePinIdString":"1","positionMil":"410.09755,89.02502","isAnchorPin":false,"label":"GND"},{"uniquePinIdString":"2","positionMil":"194.10333,89.01923","isAnchorPin":false,"label":"SIGNAL"}],"pinType":"wired"},"properties":[],"propertiesV2":[]},{"subtypeName":"HC-SR04 Ultrasonic Sensor","category":["User Defined"],"userDefined":true,"id":"f7a95729-a811-496b-83f5-7789de376adf","subtypeDescription":"","subtypePic":"5a738b76-89aa-4728-b8e5-f09c859dbb14.png","pinInfo":{"numDisplayCols":"17.75472","numDisplayRows":"9.29339","pins":[{"uniquePinIdString":"0","positionMil":"724.31191,21.31240","isAnchorPin":true,"label":"VCC"},{"uniquePinIdString":"1","positionMil":"824.30674,21.31240","isAnchorPin":false,"label":"TRIG"},{"uniquePinIdString":"2","positionMil":"924.31190,21.34367","isAnchorPin":false,"label":"ECHO"},{"uniquePinIdString":"3","positionMil":"1024.30154,21.35407","isAnchorPin":false,"label":"GND"}],"pinType":"wired"},"properties":[{"type":"string","name":"mpn","value":"SEN-15569","unit":"","showOnComp":false,"userVisible":false,"required":true},{"type":"string","name":"manufacturer","value":"SparkFun","unit":"","showOnComp":false,"userVisible":false,"required":true}],"iconPic":"ba153158-cccd-4fb1-9320-38bebad1b7f9.png","componentVersion":2,"imageLocation":"local_cache","propertiesV2":[],"hasComponentImageSvg":false,"componentImageSvgUrl":""},{"subtypeName":"Resistor","category":["Basic"],"id":"72c75556-baa3-04e7-55a5-e13f447c8c5a","subtypeDescription":"","subtypePic":"bbfae99c-8036-4c5e-89fd-a87441410720.png","userDefined":false,"pinInfo":{"pins":[{"uniquePinIdString":"0","startPositionMil":"-120.00000,50.00000","endPositionMil":"-250.00000,50.00000","isAnchorPin":true,"label":"pin1"},{"uniquePinIdString":"1","startPositionMil":"120.00000,50.00000","endPositionMil":"250.00000,50.00000","isAnchorPin":false,"label":"pin2"}],"numDisplayCols":"0","numDisplayRows":"1","pinType":"movable"},"properties":[{"type":"double","name":"Resistance","value":200,"unit":"Ω","showOnComp":true,"required":true,"validRange":[0,70000]},{"type":"dropdown","name":"Tolerance","value":"5%","options":["0.25%","0.1%","0.5%","1%","2%","5%","10%"],"showOnComp":false,"required":true},{"type":"dropdown","name":"Number Of Bands","value":5,"options":[4,5,6],"showOnComp":false,"required":true}],"iconPic":"a262aa33-74c4-460b-b0ad-c746896f6744.png","componentVersion":1,"imageLocation":"local_cache","hasComponentImageSvg":false,"componentImageSvgUrl":""},{"subtypeName":"Resistor","category":["Basic"],"id":"72c75556-baa3-04e7-55a5-e13f447c8c5a","subtypeDescription":"","subtypePic":"bbfae99c-8036-4c5e-89fd-a87441410720.png","userDefined":false,"pinInfo":{"pins":[{"uniquePinIdString":"0","startPositionMil":"-120.00000,50.00000","endPositionMil":"-250.00000,50.00000","isAnchorPin":true,"label":"pin1"},{"uniquePinIdString":"1","startPositionMil":"120.00000,50.00000","endPositionMil":"250.00000,50.00000","isAnchorPin":false,"label":"pin2"}],"numDisplayCols":"0","numDisplayRows":"1","pinType":"movable"},"properties":[{"type":"double","name":"Resistance","value":200,"unit":"Ω","showOnComp":true,"required":true,"validRange":[0,70000]},{"type":"dropdown","name":"Tolerance","value":"5%","options":["0.25%","0.1%","0.5%","1%","2%","5%","10%"],"showOnComp":false,"required":true},{"type":"dropdown","name":"Number Of Bands","value":5,"options":[4,5,6],"showOnComp":false,"required":true}],"iconPic":"a262aa33-74c4-460b-b0ad-c746896f6744.png","componentVersion":1,"imageLocation":"local_cache","hasComponentImageSvg":false,"componentImageSvgUrl":""},{"subtypeName":"Comment V2","category":["User Defined"],"componentClass":"textbox","userDefined":true,"id":"9a5a4baa-44d4-4aa0-8d82-488487322b20","subtypeDescription":"","subtypePic":"c88b2895-5e8b-4a57-9f9a-b80dd50058b1.png","pinInfo":{"numPins":"0","polarity":[],"pinType":"movable"},"properties":[{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"text box (click to edit)","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"backgroundColor","label":"Background Color","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"backgroundOpacity","label":"Background Opacity","description":"","units":"","type":"decimal","value":"1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"textColor","label":"Text Color","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"fontSize","label":"Font Size","description":"","units":"","type":"integer","value":"10","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"font","label":"Font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true}],"iconPic":"d3694a2e-5bba-40c3-8069-8db85c4c9209.png","componentVersion":1,"imageLocation":"local_cache","propertiesV2":[],"hasComponentImageSvg":false,"componentImageSvgUrl":""}]}PK
     )u�[               images/PK
     )u�[����^� ^� /   images/67df6019-bb76-4308-bacd-6454b246d44a.png�PNG

   IHDR  �  �   vEj�   	pHYs  �  ���R/   �eXIfII*            (           V       ^   1 
   f   i�    p       �     �     ezgif.com  �       �    �  �    �      �w��  �iTXtXML:com.adobe.xmp     <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="XMP Core 6.0.0">
   <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#">
      <rdf:Description rdf:about=""
            xmlns:tiff="http://ns.adobe.com/tiff/1.0/"
            xmlns:xmp="http://ns.adobe.com/xap/1.0/">
         <tiff:Orientation>1</tiff:Orientation>
         <xmp:CreatorTool>ezgif.com</xmp:CreatorTool>
      </rdf:Description>
   </rdf:RDF>
</x:xmpmeta>
�[n  ��IDATx���	|]gy�����w�ڭ}�-/��@B��B�Z��RJJ��a銁N�$$��t���@[�a�RJ
ek�eŉ�Œ-/�"˖Y�,k�s�׉IKbk��9�����J�%ٺ����<�'Q�z�T����g(K!�ُ���l	έ���                      ��	hI˺��{WԜ�Ҵ�'��mJ�:���gp=�b��L �E�(A��{5�V���˜'�|�v�s��ޞQ��d`��o�                       ���O�?+�m��v���lS7ކt�y{���#Z�Qe�$�2@l�êtv�έM�.����_��Q�ݩ?W�n                       ��fk��g3���=�y�иs�����񧝷���l�Դ DA1�d����Q������p7)�����ʻ�9��                       ���l�v�7�	�m��8��;�>���9�[�� �A1~���T�6;;�;;��5�lR�s�z LH                        �U��v�� ��p^�;�_!�@Yڭ���5#(�OL0L��ԲM�2�0Ζ@                        ��Rg�K!g3f��������?(K�کeX1�b��A�*�W8���l�tv�)7ҵ                        �!K&!�l��5�)=�o+�ojI_ӧ5! 7EP��<�$g��
g��Fgg��#U                       ���V��[��?��9����}UOhP ~A1^�SA��Ev�O;)rn                       �A���*`��k����_VH_�c:  A1n��p���|��ى                       �]�B�����7Bc�=���A1n�*Ի4��wޫ                        ı�1f{H�S@�ղ��'tU@�!(�v*��z�s�g��&g��                       �\�ἾCA}F;�E���Q=% NHK;T��ޭ��yo�                        p+9�����m�~����2�E�Ԭ #(&�g'�s�g�w                        �F�
9ی��C��J�'��N	�!BJ�'��u��sy�s�.                        \r����_�}�y������A1��S�����C��,                        DJ����l�j��NA}J��{|���Hy@I��;5��v�+                        �%�lwk����ۿ���mFPL��tv��S
�:��	                        �Ћ����}S��=��<���py6 fF���                         7y���fc���Փ<���pxX�׌>���                        7{��է����}ZGx A1���c
�.                       �+���6%�MzH�D��ь #(f->�\������^�i	)�IJw�e'�)˹���no'���1R�IJ^�;�;�-jqyɾyiN�PHˡe�.]�3o��hzqV3�Wu�y{i����В                 x��`��q75�ٶ�ݹ���)	I
8/���s�	JM��n����P@���`߿�4�n���U�vnyA�LM����g�׸/��W5��       DT�z�����ǔ�?�N-p!�bVc���������{E%U�����<��>��9��:ϵ'�	1��f�����]�����漽v��m�^ԅ��                �G0TAr֍�v��G�s� T3�4��uq�Θ��g��O_���W/����g�`U      ��Fg�]ֻ��ޯ��o\����ڡm�џ*�������BUg��n%�L+TAr����(=1�ni���&����s::{FG��v�I��Թk�                p���1u�j3K�׹���يRsb6��VR�Ub��<)���|1�dc�\�����gj�Ok����      �RH]
��ڡ�jI֧uQ�Ks+*M	�7�_wދM��G$�Ԙ�Q-���(��0�i��=Y�V��i�}fS���8{����I�|J��㚘;/                @�A;�5�Ru�<�DU�EJ	��5��엥���v�����Ҽ�͞���I�]��Хq;0u9�,      �R��P����W��+\�������в>����������2�fW�-�J���߻Tvb�:sk����5z��/�����I͇                ���d�f���Ը?�e&�)^�:�MY�vS���]]������>f�c����U     ��8ۗ�C����	1��7�a�hAײ~�y/(X����:u�5�#�J����3a:�74�͘_^���I�>�=����S
9/                ��1�N;r�m�{gN��Ӌ�p3&L�-��n�rhYG�L���#�s��_:��e��     <����;�CU�>��Z��g;�j-��P����"m�kҖ�Zu�T+1� �]r0��?���/ץ�Y{B}��1�������                ��JS�%��n]y�JKH����e����e/��Q/�k�������=+      ܐ�l�֌^����N	�2�b��^�(Isn}���6B�$�wmhЋ6�h[^��3���NJ�mv{�B�9���G��s��P               ��K{N�n/hUW^��R��1�Q�����W���)�]8��Oi�ҸB�      �J-iP��)}A@c|@-J�_:�6+%�-�Nw���JO$Q=����r��_�r�ݩ}��~�:%                �UE���SwmV~r��iv{���t��%}����{vPC3�
��     q-W!��v�u��_�검(������{���{¹��8ՒU����e���W�|O�L/�}�/�۳�1�>�O'��mGڔ>˾��hը�3��W�7��D�pk�2/i�jD~t^:F;���,�\(�@݀�R��W�g�Uz�T��sy�tx�a�U�R�:v(�nn)aI���i1qQ~U{�V���'�Nh�pB~�>����mb�ح�'��麧���o5iV�,E�+q���.�\�_���~�^���i�5\;,?�4�I)���R@�ҕ�+��bUNV
�v>�����W�ˉ�tp���[.k�~�'�˯�OW��\�pkE:QxB~�:���C�
���-$.h_�>���cMʾ�-�ڑ�G4���59Wr�x��sO+`�CuC�3�<�v-M��@ ���aͤ�ȯ��;��	֗+1�=�ъQ�Up9��C�J\��r�[����K�omC��
��+n�t�i/9. L8��m���S��w�O��K{�v�ڴ���0�1      ��J��zX��S�w�W�~M�Z��QH�SՐ������[�*g�M��ṡ1/��7N�ѷ���ܒ~�.�G6+�r��2��k_�>_6�L�}��"�ʘ�P�T=����Ƅ�t��V�<E�+�3ԣ=-{4�:+�)�,W�	|W*c"CII��J^LV�@�����������ݾl�3��&D
+�4ޤĥD_[�c�m��l!6n��mܮ��>_6�m:�ɆObe���`�/��6\�`����w%̾!�@��l~R~c֗]]J�F@�Jmڦ�M{5��f���e�8�}���sO���ߘ�s�)e� ���>�C��i.��|u��Tq�BX�5��~*6�ۻ����L��J�6p�v���b�A��:�?M@�J�i���&��T�s9G�#�vm�[{v}���/?��R�l��2[l��b��W�`BbL`5�˕1����d;��o��r����U��VK�/kLi��jae�P3(f�̿A�p���L�DA�^[����
Srn�Ƙa��8�����..�7�     �&jҿ�!���c��A1�f��2�8�LT�&���K�sj�DxWC�F5�߭wռJ�9;������e�s�=�t)�
�T�a�X�f��AM������B*�N�L�-��S3�Tkc�㻆���e�f����G!�ڔ�-����/�4gۨ�D��j�`?6�c��sŢ�zu�N����Ѳ���m;�M��:�a��zzl����b!]=���v�M�h�`R~q#���}%�o����/!]�ud��5�ӅL�4�An��)<_��P�j���g�̱P�b|^�\+��0����~ͦ����ҵ��������g���mUB�sO�a�{�;�˶�ZL�OX!�k���6�cɓ'����M֕�����>�)_���2�24k5lm��M�����F5�7�oX������� S�`֗&H+g������i�����ɿ�T�*'*��3�ъ����h娀H0��͹������f%X�{�h��կ�;�^�����3O�熵��5o     �HV@�j�^�DݯOjZ@�_��C�OK�������EzmI��,�Tf"��~���j/��md愾1ٯ�ݯ�K�B����|cm�֙�3�:�9��i�3�~��G!����-�[|3��Ę���	o,9WbS~h�c����h�k��l����Z���!1kUu��>_.�����+96�4`�RR�;Ыݭ�h�#�t��:��X�Ԙ(�~X�	!m9�"��9Oc&���x�������|#�����`�{�D�jN�E�D\�O3_�b�z	�Y+�.7A�{Z��b�{��fO��\�5�c�mÄ���ٷ��e�n�'z�Z2!���p���Ƌ��u����ٷ��hw�nϯ/m��VN��6j-n©�T���B�>~�C�����eo�^ͤ{����x���B�V&��<_�T����,��x�^S�Mũ�����l��d��s�O������S      V�Z�n=�7�	
���
����^��(���ڲ�tO����k��𿦬r�=P���ٽ�ʉ��5ưvR��)�n=ܪ��M�{���B��0��z�zl��WQH7&�7x���B���C3Ӝ��6�z���L�Ϳ�/��9�������^n�˙��惄Ĭ�	��>�]��vy:,�L͘%�t���5�f��'�U�ѻ�X��>���w�W��vk9��	�����9n�4�I�u����n3_��jUOT��f���T{^���	.mX�ޖ��I�n�	�+:Wĵ�u�C3!�ᑸ������ާ��9yն�mʺ�%�O͉��:VrL^Eix�ϥ{~}ij����c�����H���/©:U��	BH����:�/[���4Ay&��a�lmÁ�׃�3�[�@ix�N��ǔ	֣6�Dw���ś�`?JR���Uw��ʗ���ЗO|_��O
      N4*�j�ީ��agX?���q<�&�2��/-��[�nWuz���S���^������X3
�¯�h�-�8Y��#Ӝ�+�j����f�M棐*�Lv��N�h*�{�|R�������^��τ)���������6���f���q��6`���Ի�z��|��&�B~u'���x�qy��3�x�Q��3���f>BH��<߶��i�vؓ�|'T6Y&��������m��Ya��:}���mګ��/o����/7�B^&x�{����5�콠bBz��p0ǐ�'��}�p�ay!��e֗��oW_G���
*6!���e�B�!]�S�����1�����Bxd�f{v!��e��7�l���A8���W�B����Z`��
��pGA��g�����Ӯ�
�B     �Lg���g���)o]��k���AuiI_sn�ȇL0ȫ���-�/VAr� ���X+
�"��X���AO5�I�f�3�˄��6t�v���L3�-���#�i��P�mИ��NX�T�a��<�4��,<�̷et�m�Bx�f>�}��;�|E��z�U/s?0E�{��xf�;!��a���N�)i9I�7z���|�\�'��2k����e�.�4�Bf��z��6@M�{��τG�)��i���Ҟ�=򊌹gBH	�	+;�}d��5x������b3!��a���D�ͦz#,Ƭ/���~-]�ت<]i���+!������F������m��mv�Wӱ&{]�D�	y�9�d�?!��8ǜ���a}f�a��&�j*�;���FF��u�v��Ƨ�
CP�Bڲ*��z��^���N��7'��|�k     �52��ߧ5�Cz��w��Z���~P�QP_rne�g��m8�ݥە��,��<{2�Е	}�ط�����#:(��</5�1�9�R��ئ�����n
�lHӶ"¬�ڏ�kxiX��r;Ә�?M!U����4��\�Q�H'�:�f���.e�f
�Qx�P���h�+>_��#Ls��`'���k6���|��F^�D��f�2�7�BYII�>�݆������IMG���ɂ�r;,W8U��2B2�2�����>�7�e]ɲ�BH#���v�뉩�7�@��˹Bd�f��7멆��v�6��a����mh�L���LH�Y�ͧ	�Q1Ya�9�T������2�������|��,y)�^kM\�w�[,՝��ǒ^��8ި�g	!��}p����\_�@id���mcm�֙�3r;BH#+o&�s�p]I�D��x��V��'���aT�Q���߭�W�T_8�]���~-��     �c�Ւ~��.}R����W�w����g�ƴ����G��ߡ�D&2c��3J���{u`愾p�;�!�1xS��3H!U4�f>-K����4��H]HU��^WO棐*JBR˱��7Q���﶐j�B�H�B3�)�3����,S����&�ۧ9��1��W3����d>S��0���!����!wO~'�4:�c��t�4Z5*��;^��3Bd���7�B=�l�x�{��i�ax6D�9���f��+96���9��Cm��T�{�b!���K��o�#�4:�mޢ�M{5��ΰBH��t����ʭ!��l�|�;ח�6D�9��A8-G[T4U��2�L`���d�fhہm��;"��Z���s|��m �4:� ��o���@�^Zԡ{+^���<+U���_����G���|RK!ww      �A�����ޠG��"������>����HjB��.ݮ{�oWf"Ӳ�v�Y���z��.����KO]toA��Ls����<S4Q9Yi��G+���g����SH%���4��js��w��oCb(�����&%��4^�f>
�����|Ls�.sh��5��f>;�y�[i�X�F��'�-W�8Ӝ�ń������{5��f>�9G�Ʃ�v�|��ܦ�x��ϔ��l3__{����&��v��V%�����5�X�X�1�!����f���|�l'$&J�y��#�^�d��܆��rs3_��2B��0����lվ�}��鮠bs�<�%/$�a���C����B]&x�\��o��l����Mm�	�'�4z� s�>V6&�!�4�� T��A8��FYHj:�d�%O���B]YW�욾�ٽ�p��������W�,5_�Z���}�w�m�/�O|��     �g����a��>��Xum�T�f���=�`�޸q��)�C�I�¥5�R���s�{qL~������<
�bg�ٍ�He�jDn�r�E������$�����ݮ��G!U���Qh9��%��]��y�B�h��|�=v���f>3͹�H�]���m�Mõ�:�wFn`B*z�z�z-U�.�̷ux��lqOXLթ*�L��e��l�SOi:kZn�4��)�*Qp1���!�E��fO���6��׽�[����MqG3!��a�!�OV+a1A���NHLl���������*�($�k�!s��nCH��6Gi������ذA�#���~�.�#,���)�P���N=���������e�̰�=-{4���e�\�m�7�=昽�t�]_�V�g���0nn��3����m���c�|�x�{�B����@�v7�a1�'��6����*O+.ũ�60�'7ަύKߛ     �e*����O����*k>�]��Ћ���􋵯Ui*�9[r봹�V�?7������3D���m�F�X*�*��kc�B��2�1{�z��uO�'�QH[�ز�d����t�,��|���ʘ��*VL��[��L�w�f!6̾��p��4��f>;�y�G��Ls����l�c��V}�Z��Bl��ͣ��O~ϊm3!��Wt�H	c	�_�?�?��+:Wd��}��o��|��Ɩ9������o���o��2�E9�s��pS3_��"�ib��X����4^�f>c� !���7�/[b��W5Q��S��Ɗ9n0׉�5�;ӟń�vt��g����<N�ds샊��4��!��bY�u"s_�I����bkL)!11�q�A8ձ�c�5�^�b�M�pL�KǡBHc��D��7+9ӟÆ�:ǐi�!�����m�6�j��A8����R���ujϮ)��������	���o8o�3|      LL��!U�q}D�*����#�ӂ������I�j^����`S��Գ�Q_>�}}���4r��D���|��7(�P���v���g $��KAmܦ����5�QH�f2��=������3��=l3��v[P�f��g6��x�{MG�����'b���4����6�
�e�-mXL'�՟�W�$Ӝc�6�n�`���rb��g{Ms)�:��1߆=��T�~��ȟΧ�/����G�{l<�L3_U��LxQ��L!�l3�3a��j�+>_l�{5�kZ�xIl+L��i�KYHb+}.]���}c��gHM)bˬ/���4\;�3ygb�3B��W��ux��l�]X!��Xh���mګ��ج/��di��V֗.Pz�T	K	����`�!e]�b��ў�=�K����`CH�Bk���d��7�j!��r-�FP1a1��!9K�U�L�)ު`�냈��r=���֙}��#���     �+}X;�׏9o��~P��U���sk�<.+1M�U�Lo(���9b"%�t�N�6��c�Կ�yZ�PH��9�O��u�v��Ƨ������.�N~�o�ו�+Q��R��)�2a1fj�Het��(�r���g���wk>1��|&A�=����E����i΄ĸ�	�1Ŗ}m}Q/�4�Q&D
�`���i�nXgr����4g�ɝɍ��wBH�%��|���O�T�m����7vQL��	!�;��&����/��|&��a��}�K��C��:�Ƌv3���߭�EBb�sl���:���nPqÉ�M�	�`��GZ�����~oBH�'{6[]�]�Ӷ'�߻�`��/B�f��	j�׸O2/D�{S��>E�<�@}��B�.f}i���[�5��A8����9��<]i��c���cC�{�<�,�C�|�z�_#�� DNb Aw����/Wz"�u}�9�΢N�8�E_9���     ?��v([Y���ܸ%o�<�
�M疧�ۛPs�˕�HC.b� 9[7�Y�*ڢ�>�w�=+��	��߅�f���G!�;�b�m�io�^ͤG���B*�*=[j�T���c��{�f���6�1�ٽl3�r�o�N3�i3M!fwI�O��^&H*Za1&X�p��F���|�[�P����i�˘Ͱǭ���b&�wu���/j��4m�^���F3_�>]ȊN3_�t�����)<_���v�E��τ��}Qڵ4�]̔�h7�B�^&��K��E��/y)ٮaY_��	�����f���z��%$�uBR��&{,y��dT�%!��9���!g�м��E�!�D�ۘkU�F6i_���̉��2&_��	�q!���|p��jx**�Ϭ/���~�R�yvΞ�=�M����?��H�ܧb�A8U���l�vw1�3�bW�.�b|d��&���u*M�k�	�v(��;�G����     �#�ь��S?�l�d�My�
��~&$�NV�^�4�Q�Y�fSN��p�/�'�M����yN�2SP�4gw3�|�Ѳ��?���4�d\���6���d>
�ܯd��T�F���i���f���u�8���*&��ϲt�<�a1f��9n0žp�ԅԨM�k;�f��9lp)��w�IZ�&
#�4g�3���n���E����@�2�B�V����&�|3!��Wp�@���z���~��t�Af�0�)��|U��T3Q#��9'h�bl3_ed��L����NH�{��Q�@�#�O����2���Y_�Xñ{>r�x<�߇R�K��n}���"T�et�rfrw2�&�g�nPS�S�^�7��P;�/],�RnT�����64�d����ro�^ͤEvN��r[� �*�*��k#�}X_�_�bҍ��ɑ]_"�r�2����΢Nn�1m�>�v��75h��N/\     �Oܫ%�ݧ��/��WJT����s˳#�	zsًt�˔�����W�)�C/.h���[�>"x�)�"$���dEt2�-�`��ܘ�����RyG��u�uh���|}�9{G4���~���n渮r��[�V�F�{�i�[��*!DH��Ec2���<�4g/hoRR(I�E�i�c��w��x���B�H5�uw��N��]_�f��AM�E��τ�6�7�7��f>s|j֗�Lsv�h4�U��V��j��Jϖ��U"��S�Sm�!��gB��8���]k�k9ܢ��E
XS�]͉�o8Vr,"_�R�0��IEj}�5ܥ�YBH�Μ�nk�p��䝉��0��G[��� B:Э�BH���ު���t�tD�G�D�jNB�f�@{�=b�p���k���#�n�w�;ԫ=�{4�٠bD�mzo����.���}uKn�����7&�
�     ��(K�ک�9[d'
ó�w��C*ג�)�ĴfW��oTez� �(K��'�ΞD�ӣ����k�7�B�#Ry����s �a1���43��;�d���L棐�{�/�G���i[�c��)������|�Y�SLs���g7�f����N~ϸ�4g���d>Bb���x���o�c�����ys��B:ح�9BH��<nۏ�k�y	w3!��c��Lד-a^_.%�I�IKI�7���-�[��i�f2»��?^��3��zI�T�		w3_�|�%2�3�	K	�ZB[؛�:v(�R>�<�C�Я��.?֯�3���	��ԅT��jw��wu����oh=ܪ��M�O��k�/V�f�;� ��k�km!��c���s����©>U��j�;� ���N=��tX�.!��\
j��6���Gl¯85W﫿[�r9���LL��ۗvء�'��	     �ެ��s���:[d���Ӽ�������?9�<�՜���wU�J�/��d&����K�y�o��V}
�F!�w���ۆn�S;���G!�wݘ�W7�3��i�3ET��
�c���C!�w���p7�iQ�9�9{Q�T�m����c��w�c���iߣ�Ĺ�|�m�۔5�%xˍf��.O3Ӝ����6�/�wi1��f>c֗��R�	)��|��zW�l�=n0���`BHͤwBb��N~��f���Fj	�1�|c�_�?,_/c.î)��s��k�K{Z����φ�^"��k���r�Ҟs���4!��:��� s��I�j���B�C�]#�ԋ��6�cɓ'�����c�x�2AO�C��ݾ[�a�O5!���C.��\W�<ة��M�gNÉ�Mzv�`\˛�km�]_1���r�K�����~Ep/s�����ʗ+5�CxӦ����_��:�/��S?T�\     ��ӌ�[����+�P�s���V�<�1�Lnz����x]aJ�>�v���������4��i���g6��x��])�Rl�-�ZGXӜ���d���7�QH�}&,�6i��Y��1��=�=4�xX8�����}�
�>�n�o�#�r�:G:)��0d���[�5���f>S��y5S�&��w��珕���kB�}II�>�݆�����4��&�����L3_�b�N�X��!���LP��i޽���6�t���������r�EESE�/=,�b~X����d����z�9o�=�m�3i�*�2�E939�w� �x�Y��!������;�k��^'`�1�X�Rok8֠�bP�K���딟-W�x��]���~g}ٶ�چgBH�ynxTHj;�f�L�o}ij�L����v֗-�[_�@�m��2�3�ý�{5��A8���L�h|���x�	:zO�k՛ߤGG��s�.	     ��ީ�4���~�፫��U��Oέ-�Ӕ�ƍ����W)1@�4��΢N5dn�'G�����B��(�,W�	
�� u!U��{mA�Z�����#��O棐�?2�2�=ح���55�1��?LsƦ����n�.�-,�i��Qp�@���z���5�}s?0�A��x߳���:��Ls��R��t��*&+lc�Z�����&,�6���|���lH��n�,�u'���Z��!��}p�������g�mH�2�?</�|�:�?M��f�u���\���̈́��@`9�-�[��i�f2����5ܥ�YBH��t�Ԯk���	!�s�����iߣ�Ĺ��}�~�3أ��d���N�)i9I�7^�߯:U�����L��m�iW�.-W_�@��s��G�5�4�ɂ�5}s�P|����dϮo�K���pl�SOi:kZp����w+;�k���9���-������3�_      ����C��>*���yPi
��έnyLQJ�>��S�ȩ�W���������_���B��1U}�Z�'��0a/�agW��&�SH�Of2��������QH�?&�e-�|�L��shӚ��LQ]��\�?�f����W0]���v�?L�	�Y�d>c� ����(9[b�/TX��c����f���1d{ߪ������3У�E��N�ʘ���6��B�YBb��<�Ǹ	�Z���Y�nڪ���b=�|6�t�R?1a1��r_kߪ�^�L������#��od��5�Ӆ����P���?
��}�]u��{���GB�f}i�!���k6e�A�f}i�\,2��O*&*�s�X�ت�^��jUOT�a��{���z!�>�Z���k�>�r�E��m��ɹ��ΑN�!}�/l�|}}���A8��`��U�J���W�_e&��ךߪ�3���c_�ե��      p���C����� �?(&����y{�<掂6���ne&�X�K$�ʗ�=�J����]�$�F�ZUNT
�c�%{��ڂ���[_�����jN���c%�V��R��m��^l��f>�m��)�k;ܦUV���u�K�W���G���B�7�����4�#-���v2���luRR	*9Wb��+k�c������4��Rs�IH�?����R�J]HU�@�v�����4�o&�ԗ���G����j��LXP��v��|��lҾ�}��s�f>B�/Ӯq�܏
.�s�SO7>���'�Կ�uHT��e�fSW���!1K����y�8]a�9�V����ԟ�W�d��?�nח�5�x��BH���X�*/Z� BH�k��p6\ڠ�C�/}��N7�n�`���rV7�ӘY�7�Ee�����E�jˮ�#��WC�V7�     �UzD��煸����z�y�3��@�~��.��x��x�9�V����_G���W7)
�W�^�g(��3���;ԫ=�{4���ŖR��)��>Y���.���w
��/u~e�|Ls�?�oXi3Ӝ�/�J�����7o�+�*V�f���d��������̱f�@����*���f>�9��J��̱�i'�ԿV��G���� Ӱ��m�Mח�����g�'�O���!�?s��w���A�E��z�U�/��wh��5����|�ܔY_�@{�W�L��}��ɛ~^�D�jNB�g��]_�m٫����<������_�nT`9��ꑛ~^�x��\�W�R��lW_{���^��!�5�kZ�x��~��g�8k$u����l�d�l�OvΡ6��L�!��\�"���UJ����R���G:ީ?=�O��S�.      �2�X�L�׷����
���n��CR����l~���j@��NJ�i�_y�;���u�\����ͶɗF�.�mp�N~��*~�#���J[P�B�|R���7�]�Z����i���f�|v��`�����qAρ�n���a1Ls�����`���w2_�R�-�M\t�i"�ϭ��N4�l�L�?���=�m���̗>�n������l3��|1R���|;��ɢ� i1I���B�'������BGHL|�;Qg�/��g�G2f	!����g���b����!���6�i�vXg�~��φ�:���yBH�A��lmv֗-Ͽ�$�4~����T�S�Κ��?7�Q&Ԛ��Pz��>�>`�©Bj‹Vս�[�m��;���a�!�N�)i)I�˞Ζ�-ʹ�#�_�����eˑ��̾��p��4�aB����d}��'����Ub A�}���������y     xP���>���q˝@;�Z���M95���{��DA,u_��T��Q�����8'D��8^t�H� �3��N~�Rs���_��q
���5�m�b��?��nT=���i���������ү�붡�l��s���NW��$Ӝ�JHv2�iИ��QXL�b����Wďj�k<ި�g��O̔�-�[��i�f2~�1�L)!1q�t��>��f>Bz��xb���z��}���nBH;uBG^�����d�b칧��Z���Ϝ�lo`�G�C3_������i7�Lď��l{�`�K?!��ǜ�6�����Bօ���!�\ě��jk�����v�M��	��'��6�i٣����B�*NW�cɱ������.e�f
���ܮ]m�q!�q($5i����B�b"ic��v�Ϩ:�X ��t�.�T��+�Ϟ     ��kI��u�>�3B\r_��U���$Ot(�`�7����5�VB���z74��7��>1�W::��L$ܘ�L�L�1Ŕ�l��潚I���*��f>3���z3�T��4unڮ��>��G!U���̷���_o��V�B�R���(�4a1f�����c��G�5�4�ɂI��i�9/1�9�f>ۤѶǾ�4��e'��l��̗u%˾��2>��f>BH�Y_�����M�%�4�=�����f����0R��W~�\���B|j:�d�%O���0=�=J\��%~��	*�a1ͻM�!�q̬#;v���TΔ2�f�뙄�ħ�����SO��m�4!���ww���'5�6Ci3�s��4�F*��1�(���O���c��q$�S�x��BI/¯'�Qjz�29�<WEZ�>��}��W�o�     �A�
��S/u�Y!R�*Ѳ����Dgszb�nx�^��" ϯ,5_Ot�[��k}ojPST�{)W�_����V�m�a R�73}�m�M��(��4��f��q��!�UNT*�T�b%-$	�+e>�[��=���Ls�k!�e�E�K��:Ue���2�2m!���*�. $&��f�M7]__��#$&Ιf>���<��̫�8U���߇�t���jN����f>s�(�P`�B������^;�b�B�o��}�|��6�"~��&�|&s��x����h�QU��f}�L=����x2�2!��,�Ж�-:Vv��%Tz��ֻ�pbBH�۳�pN����j��(����Bx�c�wT�\?]�;��3� ����������}�Y҆     �1ݺ��:o��{��P���E�'FK�'g����.�T n.-!E��t��"�_���o�AHS\Y}� \W8](�0�[����`��)U���f��)ְ�m�1����0�Z	�aח�4��:���Y�x��4�K\g���H\LT�$!����t���Sv��I��f��i@��;U���	�a=������(:_����Sv���
\?�<SAPL�$�������v�9����⥪I/�'G��k�     �ޮ�էO��B\qO�V�s^�DP�QlCb
S�v��)���e*N����[-��               `����Ѷ��-�R V�E�-�d�;���ԅ��     �Ճګ'�!n�#(�a�ݹ�W�-�^���6�'��꽲x�Y��_���9               X��i��U��/ �לU�'6�[�=�y�Ϟ     ��$*�/�C��#:!ą��<�MZ�g�뽶x�~��J`�6��걎_�o}^g�]               ��k˪�G[߮�tX���<=�����/h��     xH���e�W/�gtM���|DyZ�W���J��w׼Zo.{� �GUF�>��n}t�/t��)               X�;�:�`�O*1�  뗙����v��8�����}     �^%�q���۠�y�����A{���E� �6$g�ю��ǆ�J{/�	               ���Uڣ_�}��� �OR0Ql�)�&g�'�M      ��zH������k��١��o���d��4�U��
@d�&$����w|I�~��                ��{����W�R "�0=P��&e��g     xF@����1��b��ן�����h�G���Y����6}r�+��Ԡ                ���*_f7 �gB��b     ���*���z���%�������3��s+K.�����-o���Z���@�~�����ϓ{               �@ �j^�7m�M �ǄŤ'��ƾ���     �zݡJ}ع���/E?(fF�p^o�Ke&��m��%�B �+���Tz0E3�C               ���ؾ��n��x� D�]�=6,汃�OK�e     x�������EӾE7(惺C��k�2!1���N�g�
@l�i�}�M[�ۉ]               �U�y���&�Y�) ���g���~�ֺ     �\���>�-zD3��D/(�C�Ғ>��J������^Bb 0a1�T�:-,/���               ⍩��պ��\�,���ġ�V(DX     p�:-���/	����E����%�����Ԟ���K���{�ߠ����׳�               ēwU�R�/� �xU�]]��?�{     x�/�a}Y�ҷ߈NP��ڮ�;S�	�͖��3�F �%���7kni^?<?"                �l՝zK���>o,����9}��U     ��
鏴S��6'�B�bv*Y3�3�V�\ƄP|��ԓ�( �t=������T߅��w%%%(3=:�d�0���W����JVB0 ��8}�9�E$��$*=�u��?�ڵ%��-
�����v��ny9��y!��R����}��좮-,	���ٻ��������Y4�mɖ,۲%y���ر�A�
Jp����H�r�5���+p�
d����@[�VRL�=�eK^d���K�e�w�Q&�JB4�<#�z͜$h�F����|���S~n���7�9��1�ɖ���P�_�u��sv�gS]0���)b1��?��D5:��2�r���e�����HDQ�߲)/
(+��kO�Ȭ3��2��r������3��!g߀�
��1f*�/g��eTH���t�.�0q�)�Re|96>��Y��g��|V��)|�)fg���8��d��
)-h���1�'f`&U��m�����$�_&[^n�l��`Ɨã��5$U��/'����4מ���p˟�8S�c�`�w�<O�s3�A��     �\���)g�)aQH��ڣ�+�y�,�s�n��3��d� ���b�j�;�W���#�-BjZ�$[�R��I�c�jn�ؤ�dg���వ�͒���^��I�̟I��U�*�KS�⹖�Ój���̤;��5�v�o4�ɦ>�����I�u�
��2��<Nݽ�j�V��S�E�L��{�j����o銝���Zz5<&$���kr|B᰽�s�0�p�d��ڶq�fg�e�A���VS۠F'�$�{F�����e��}CCK��&��$�(���di��~{C�#Sja|����Q_��҂v�̐����9��$�XU�#�
[|���Sg'�K7���"~��o�J߹����44*$���+559��Ǘ�]#��6�!����u�ie�LMă�6���U�3���]k���������MLJ���N��e9Z�2W���F�"jn�8s���=k��?h���\ih�u�>�|�f2UU,QV��9N��^0�'��9�?Iv�Yk��7h�M�f��e�3�f|��.[�K��D ����hbnZ?�|R      V��ݤ�z^Hy�]��q�w�o��>��B�n�6H�@H�6�[7�K��}Bjڽ�BO<�`��(�����w{Y,
��li���h�nBU<��'��މ��Og��#��+�f�ߟ����XU�D��4uv�*�l��B$&�w��bb~�{wU��ǎ)la,��o�9w`e�[6o\�õ�233USk��~��a�Qz(����g땑n߂���!�=1��ې�H��O[�'�mTlξ�S��w8g��ܐ�VYi���6[�1:�#���=g�գO�+-h�ߟ����c�;���+;+]�-=
�:���Ęq/�K7��>���Z�y��3���`��kllL1�!]Q]Y���>��Y���/�s��n�ڳ�R�=y��XLG��"�ξAp�i�����+c1&���'?�W���5�kt����XLSۀb1���,V{w�ӣO�[�1����Aq��eKrT�����+�6�H����p��1��ǜ�eȾ������X�fi<��3`],&U�&�/S���j]E$H)׬�Tӣz��V      ʧ��
���ćL).����Ƿ�G�,sq���l� ���`��zӕ���]�RS<��I)f�-'&g��=��}���⥹2���׷Y3�*�i�%�2�߯��\�G?�P��14<��As�a�E��ķ6�b��)s�-"1�2v��c_,�DbF���o��fb15�Q���[���܉���W�`Ls�:�&+3�3v��.c��9==);W��a_,f22������r֞a�WT��MW�pm�U��ZM�7����r��u��bFF#�5Q{ޞ���e��M��<��p�&��o8wo�u��ށq����SHw�X�Q�q`��XL�N�-��˨=��E/==��<���7�s����TdBp�|,�Y�){��SSsj�싏/�\�vM^^��o�/��6���q���b��M��H�Kw-/ɋom���#1�Db�_��C�w�v�3&342�����X�9g��7hM,Ɯ7�l�V0S��eʪ�)�_T_!��?j ����[�/�-5��m     ��N�*]�l�,���bnҕ���΂J]��M��J���w듇����R�����'����[&���O$�#��r��2kb1�-}���H��XL�5���b"�Gl���/��q�����m���q���̖�e��m�"�ĘǜCz"�y��z+��#1Db<2�iPln���HL�K��X�捫���4��H�7l�ŘHLO���bS,&���Db��z�,�;kO�~��2Bޏ/M$fd�H�W�W���q;b1�����">���b�<�ʚX���LN���i�VY�1����^�=y��b�lZ��#�V�/���xj~|yB>''�%�b1�HL�����9�b�Ɨި^W����GbZz`|���cÁ� ���?M���n�p��     ��b��>���U������F���oe�ՙ�t��+���4sǄ[��Ч뾯h���8���ٵ��X��Č:���x͖XL��İ��S�X�Ï�P������I���X<����ϳX��>U��">��X�Y�_X�����?F$�6�b^��;琞2���-�Ŵu)2=I$�c�vTx�!c[b1&���S�-�����z�Y��5��9��s7e�b1&s����ǂ΁��3���c�=���N�������i�\����^_���K&���J=��	�=����=�����X̳�5�n�?5=���>�=y�� ˊXLs� ���]�/�+���=61���A�=y��b�9\cs����fLA$��X�o����X���$���1���fs��=���@X�6�[�lH]�i����?�M����      ,����9۫����PL�nu�W�"E����+����]�����tW�/���e,&��!c��XL���hW(��	U&Ý���O�}��c��}+��'c���K�[/b1�HLS��,L��y�1���1"1���b��il��X�܋��� �9m��~�'����a"1���4*6���)���H�=�c1�:\���b��V"1��:���2��DyiA|�E,&�����E|�0����x�����(�Kl�Z����$c�/�c|i��p�v��],��H�Uvl�.1���~"1��:��6��hD�����9��
z0��Db:{��
�+��[/b1f|�����&s������KKx�17�;��痩.��mxg��� R�ʌ%�?ߥ[[3Q�     K��!}\w�zVHI��E������@(�Y��' ���{�95��v>%��x,����[�?19�&RY�xYn|�v,���_Db�b&^�����X��Ȕ����ƋX̋�?��x������l��~,�H�����=�Ŵu�H����ڱFO>۠؜{��im'c����x,�H]���˦��bDbl�R,�Ғ����F�#�/
,�b,���9�s��">;�X��{���cǔ�b,�pB�Db�����܋Ř;��$c�b1�=#�$c�c1�S�M}���Us<þ�&/�bL�Խ�xs�����p��;k�����Ϗ���ɋXL||��+�K���y��H����Db��c�"^�b⑘&�琩��ʷh{~� ,�sW��uo���H      ��+��s�gk~9R��O����S�,a��Y%��\]q��'zT3�$��=�+]��LEf��5�">K��i�GbX�g��b1G]�x;2Qo������f,f>�K$�Rn�bz�ǉ�X��XL<����\�������^�g6(��ݝ;�G4==I$�R�vT�����Sk'�[�X̦+]�ŘHL�E|V���T��1���^"1���b�1���$=cF���H����9{���c�v!3�!c����b�#1�,�T<s�:=�L�2\��v��jbr�kO�r3�Ĵ�)�b�/�|,f�j����Us����_�ʌ/qƗA>G���Qg7sleb1�XLM-]��b[��sƗ6��b�V�7f|��q�H���g���?��X�U64��(�ې��Z�G�/�& ��뜿���N�s�c     ��O{�q]�/�B�Y�i&�p�Q�U�|�^��d� ,N�_Y�v]w�N�GF��eb1�>Y��N�7�e22���~&RY��b����Ov(-��I4�}��`�x,fO�~��q�Cɛ@c"1=}�Db,gb1f�eW<�����K�&Y���b��]�7�H�b�ށq����P�r&s�H�Ɠ��5���^��X-''����ك�I�Ř;�Oq�w�X��4H���bL$����7pi5�b1�Db����<�x��^H�1}t,��>"1�+_Y�&3��4����Ŝ�B,�Db�F�����b�E522��XL<��C$�r!�ޙ�X�|$f�kO�s#c"1Mm�Db,WX��J,��cXss�ng�Ǘǝ�D��&����ە��#ٱ��an��ⱘ�܆��b�Ĥ�����Z�����8����H�"�1�\�_}� ,^X}�N�upCT     `�/j�~�<X(�bv�IT_�d��P����}�_/ �[A([�Z�}�з4c�}*ۻk]�b1����*��ŷɊ�4��HLj��PU��;��$�bF�"��'�*֮Y�&#c&R�$�2�BA缡2i����q���I[7�&-c"1�&�"������B,�))�;L$f�k��b��
=�L�bI��D"DbR���l\�R�G��i"�2L,�3�%-36Qw� מR�����ͩ���ǗfyNc3��T��X�Y�g"1�/S���:\מ�X����7�@��RA"��3�ξa���}cDbR�|,�I�ӑ�33���p�)%$;��9���)!5�1s��WZ�DbR�K����HM$���!�I�܆��)"1)��b�)9������Y
���}��,qC��ܩ�in�
     ��R#�J&���p���t��K�X����f.�X�6�ԇ�\�;~.�6s���'Z���u�0�*ŘXL��؂�+�)��_,��1���ێ����-���9ŘX�Y��Г���'YėbL,f�����nx����XǾ!��X��#-
�vR���/wzO-&�bE��#�����S��];+t��y��oGO����([EK�KB�enn��)��b�o]������&D�4��Y�T��S��baǗ�3�~��e*1����R.���o�e|�bL,���vu��I1&���X�c��O0�L9;��VMm�s�_�}������bb1˖�k.	�˩�)�)Č/w�f��:�{�t�^H1&38<�'vn�ܜ9$�J�܆�ե��X��}���HL�1��������?0����e�3q�Omx�
C9���o�������D9�     ��V}Rw�sR�B�b|�קe�40^Y�K��SǛW�V�x��~^               �M���D�rW	��c}�J}d����ɟ
     �BK�u��o���0����6�y�,quť��)�S�ukߨ��5�w               ��닷����S��ۯmՃ=     `��>��Н������C1W( ���{�6�Ғ�pjJ������wj::#               �K�Å���p�~�tt�M��     �L�f�1g�OH	�>S�w9�e���\}��28��g.Շ�\��N�L               �W>�n�~�2�p�
B���+t���4�     �Ub����m��z뽺P�
8��[�9_��|�r���7���g����1               ^����j}N� �2{��]~�����      ,���nr��
�{u���z��Nx[�^mϯ >�O7V�EW=w�g�               �iS�*���l@�;W���:8�(      �\�[�}VÂ�^](Ƨe������U� ~[^Z�n�z�>U�]�b1               n�
��ɪ���� 	>��ξ���n���      ,��Y}��~A�ڟ��Q�:ϻ䱐/�H� �kG�:]�|�~��                7\��*� ~גP�>��2���     �27h���<�k���>.�o�Z��L ��|`�zz�:&               $��K6�K�
 ���0����     �"e�۝�����B1�T���y�*�To^�K ��	��t㺷蓇�Q,               �Y���Zs� ���f���P��f'     `�>�<�y�0�RZ(fVw~�~y(���c�.���� El�[���F��~N               @2|��b��
 ����l}h�E�҉     �E��f����W��^y(�z-�OW�co/;[k�� ^.���3C�ꏌ               XH[���ol /��g����C'     `��;B1�z塘4��y�C�E���
 ^��@XW��Ds�               Jȟ�ֽY>�O �r�}���]����MSs�     �BL�Z��+�z�����R=�s�n�|�B�W����K6iO�=�_'               `!\Y�Z��( �R%��{�y���~     X§���l��`�WV[�Y�)���%�wjs�*���ڊ7���M�E               �k�J���=�?�ه��=���]     ���a�?��f���PLT�O��f��� ^���\�s�9���               ��U�*�� �Tfrͺ7��Cw+�	     �˕�K��	Vy���[U�i�U���󔛖) x�./ݣ���S�T�               �?��K6iK�j���)�\gm��}G     `�>$B1�y���]�<�呕K���g B����\����G               �T��W_$ X(^s��8�HtF      �D��\�U�`������Ї+.�� `��-ڨ���깡�               ^�����8�/ X(K�����=�~�o     `��f�g�ׂ5^^(�fmUL����tzA� `�}d�%���횋E               ��l]Qz� `��s�9�U��F�     �9��%B1Vyy����!�|~}pՅ�dX��L����;����?�����y������RC,��䴢��ߘBi!M�L�c`h")��¼l
�cffN��Yg�����/�@ �����!yF���o��������:��#���1��}3�a����L)�cMO/��!;+C�SB��O�q"?7[ݑ	gl!�3����8�z�?�����ch(Iמ�s��N��:fg�455������
�4;7#����7��1�?�LLN;��3�iaǗ��i����e��e*�t�I_fgjrr\HC�S����������1I0S�9V�sɅ���tdJH���I�ې��~��dn.��g�נR,SZ0M3��/S���d�ƗY�ؕ�e*�L�*b�=-��5ם���3�dn�->��Be� -ݟ�����ϟ�g     X`�n�V}^�+��P�t�<ri��� $��,�~�sP�sD#���?�ёq-_��������;�Ť 3����v/�J��/��С#M�fBUJhm�?6��}�������c1_*0����:T�,9����t�kQtnV�߉�=��('k��%K�u�h��GG��HLsK���$���d�t����|)�p]����D̅����(Sj[59I,&��k�$i�ˌp��Z;�!J�m~|��N�¼��5kf��J���k��]�$m|y�ɯΞ^�~ѹ�j�v����!��7�8��9Ɨ)���O!���%g|Yw¯�!Bũ`*2����X���eXG�[_���c]��	ɗZ��]�4Kk�4>>&�oxxB]]�Z^������[:D,&5�i���|�%�:Xע��I�~]�#�D��6�L���-��\{:��K�&��S~�3��m&�"�Z�
Ē�o�_����`?sC��':U�,9琹�!9�B,�k�Jt~�6@���l����q��     ��bz��L(�<s�v:ϕ�@��;V�- H���,]�|�~�����Q8��6�^���|RK��������� /���0��V���E3�,�Yk��f"�
�I{���e�����Y"�����0�d�kce��7k�	UV3��P0������ח��Q��\"�������
3U��:N,�z&�����D �����:X۪	��n��"1��@�^��$W1竹��X���B��#���2y�fQ�vg|y��E���`/���PZZ�ƗkW/�-b1V3���um�O��2;3�-��Us��X��L$Ƨ9���_n�,Q퉨����L$���[�9�_����u��S�s&ɵ'��HLfدd}��w��e�bR���tv*3#-i�aƗ���L,�v���e~�f��mC�iRd���L$flt\�P�=U�*t�1�w���'wnCf8M[̵��&��2�������f$s|�\u'D,�r&s�DG�F5ɒ��ƪr���ܕ�ΗO�C�<fnԕ�Ӿ��	     ��t����W���~Uo\q���r �vE���Y�������?��HLª����Zkg�X�g���&��̤�-��������������6z��XivvNuGە�¾�,�P��X�Œ�IH�bj�I##�bl�F$&aI���J?٪h�X���Mn$&�L�޶q�ԶhrrB���Ф����N�"��������������d� L,f��U:X۬ib1V��N~$&��b朝BOo�`7"1	�Y��X��c-,�TCs��I��$������;���0��l�F$&!��,��m�b,��HLB"s�H��&���ȍHL���gdM�H�5�I�{!��dƗ-�D��`����Gb֔ŷ�b��F$&���nXM,�bɎ�$��qƗC��}�p��I�!Sw�_z�*�T�
� ɶ��Z�s�tt�M      ���u���g���4>��6y �ҳ n�����������L$�`ؕHLByY�b>���X�M�'R%�N���XL�۴u��I�Z��9����@�����ֹ�I0̈́�#�}�:��Db��l�.U�Qid�X�M&&���ܣ�l��L,f.Z��ƶ�y�q�ΝHL���}���s�&�&{O��gЕHLB��<g�Us[�k�'�qnFb���F,�J&3>6�PZ��%T�Yjވ��#Fj���ms�ړ��l�Z�/�Y�g�x$&��HLB|1_�r՞0a;b16�GbN��I(*�T��2�'c��㝮DbL,f�ƕ:Xצ��1��#��EbJK��[b1�1A����!��e��rb1r3�`b1ј���I|nÑvW"1	��W�o�3;����Gbf�3�a>S��'b�g|i�9zܝHL��Ŭ_�RG�[��x�=���! ����u��#�     ���<�X�_Es�v9ϫ�7/ߥ�P� �-o-ۣ�|R��,�s����U��HL{'�x�I����m����=���L)to�eB����>�o�X����$�p��Zb1�0���@���V�X�zb161����nW#1	�K�䋕�DSv,�v$&��b�m*ס�V�=9!x�Db��ݍ�$�;�Ks�hn�`B��#1�FbL,f�Fg�Pע�ib16�"�PU�,>���'c/"1	9١����E��ؠ��O>g���?��XY��Gc��b$&۽HL����X�U⑘t����&X�mC�s٦1b1V0����ee�?�4�����/��d�#1	�X̆r�kU$�����Gb<_�]U��[Gw��#1\{��4��rgL��[��I0���+���OC������$�ehC%sܶ)�\;��	 ܲ�`���V�p�      <�v�q��`b�����4>�I�������ى������\djrnz"���b�O�f���~�?�y�gu��遴��@zFV0������/"���a]^�W�6�JH>/#1	��
�F���ݷ��e$&a>�J�ꚸ���^��ܟd��~]���4����x�,�=��I$&!�X�5���$���idtT������eKMԶ�X���&�����~�U�S�b�d"1].���w��ȗ��ss{'���q�w��αu�ty�I�^�,~.��G,�K�Q!����S�s��i=��H���D ���ҧ��W��!FꥩȬ�뻔��ݾ��b|&�Ъh4*x���.O"1	&c�=�uƗ�H=�e$&aEIn|&U���n�$B�
�u}��5kfzZ�Noߨ�UzȻk���ķ�b��e$&��b6U�T�_�1��RKۀ3���V�s꺡�Du'D,�c^Fb�܆��V�h}�K��g�����h$6<3931;��NOL�͌�Ţ��ٹ�I_@�����>(H����23��������?��{]Y�Z}��     xl�n�V}QO��O�/��l���f
����:'&��G�Gf�k�g�L�f�O�<�����{5���_�`{8<=ݟ��y��(HϮ(N�/*
�R�9Žy�n�K�������HL�"�b>utw�!�`�nݰ�X���:�<��$T�-����o�X�L$�p������f�%�/�7�*�y��޼���R�m��ww����{<��$�XL�W��Fb1^1���L��f��M�b�44<�y$&��� �%�x$�_�[0�|1s�I����&3�q$&��bY||��O,��HLm��K�ټ�\5�Z�q/מ�����i$&!>�\_��GE,�#��s����4�PT��j�$�!��H�y~pƗ�7��`m�&&����cS���/��ZiIn|K,�;&��a�4!�_n߰�X��z��448�]x��bb򩳛�x��HLBvV��8��������hm��̴g���D,��DT�CÂ�l��$�gh��r�ou��mH��yښ�F8�E�s����tod�{02~lln���\�@dr��o�?N���}�W/\�!ߙ���ف�k
ҳ�������>o�=����}Ё�     x�o������-w���e�����L��3<3m����yzxv���YS?��}����Z����gs�w��{?������,
�_���aUVqN��꧔�>hř���WBr�#1�vDb*V�狩��	Un�_��aE$&�,.ݲ~u��[��L�t�|$fҊHL���Dc�� �7��Ix��[��b\6����l�sl�XF,�&��ح�l�g$/ɖ/V��Mmο�`�M�G;��a�x"�ٸR��h�9��{�#1�VDbL,&�3w���cS$&!�ٸ�9o �6�"1	�k�ŷ�b�eS$&�D�T��Y�G,�U&��z�IH�bj�I##�b�d"1�OtX�I0��*��q��#㦣'����$�}�_�q��Ĵ��[�I0�������!���a��=�!��C�-��D��#1��������UE�B�:{z���I0��MU�t�x3���H�L$�`Ў9��Tvc�
՞����I��b*˜�N��$zW��©'27�����������O�L��7ox0)w'����7:������W�qᲜhڕy��K���m]�Y�$�g�w�}ЁB1     �s&��SxU�_��|\vQ�e3������y�g�y������w��M}o����~r}���u6���|�u��|Y+�(|ce���L;>�ER�a���A�C��#��l��$�)/�!����~��D*��%�I���[&#���m탚�O��g����ֺb՝�jl|PH��٨jN�� 7,��ehCe��~0�&T���HLB"SSצ�a���HL²�ي�LG�}�q�x��2��ٵk�O�f��^g�,�s�|$f��HLª����剦.�5G:���$��Amް�9o`|�x$ft\��]�K��b��q�OH���>R�a�"��YoƗǛ���M-vEb�9��R���GY���HL��,�7,)�t��C����ĄdM$&!�9P�C*v��XĺHLBYI^||y��]p�m����x�t�֚sHƗn�������s֮^ߞl�F8n0�K�"1	�s��U�:���'7��h&2mM$&!��;���s�`"1�'����$d�z]���d|���+�5o�pj�͜����xd�{o�?����ݫ�7'�_x�w������%iyo��.�Rηo`�g�AU9�:>ʵ     �3u���Y1��C��l_��㪀ϯ���-,n&�8����ɑ���c�?&��}��Y67��{�9/�5������[�WV�Ȱk� LN0C��w<!,�����M��]�%~[Z0��4'���`M�rsB����rs���/&$��ЄN6�*��������|f�������g�8�{�a�,�L���a�ͤ5{w�q"G�N3!���������
��58l���p���霰SBCs���œ����媵üW�x�L�ȬԴ8�K�>�B!�fag���͇ FF�=N��嫥ݜ�F����X}�,���p8]��Y<b��u�x깦x\��kO����Y;���oD�4�94[+7;K~�����2�}Ҍ/}�xߐ���<��3�ZچT�4��KO�9�3�l7�W1�L��9=�7����o�^8=�y���X�
��V�/���%�_&��Ĵ׵[�miii�mp�3����f��27O�`|�l�jl��&�-+;��.y����/�G����a>���{�ŭozd��X����_���������>�sw�Ͼ�Ї�zѻJ��W��\ʵ�x����=����     �4�����G�g~�E�+dn��z��%U.�ɹH��H�Ѷ��O����t����O���M��(ܷ6{�{�rJm��^���أ�v>��x��Є�x�IJ�w��[���3 Ƴ�:M���0;;����.H�w�d�����϶	0�e�u�����|M� ��}$� ������������.���^P{�W�108�Ǚۀ<�%�h��? ��/OMKB��y�X|���N�v���vgo�/��w_J��q�/�����y��V/��pYF�u��Vo�ӄ�圢M�v�W�bn     �O�P��~(�\g:υr�	3`q���n��eb������Es{�*�7����KW�|~[ޚ!?�Ţ8��=E�p�              �����=
���1:3=8��h���5w���Z$���?�_���������7.�(�}{~�ٹ�L��(�}~]�b����     x��\�<���>���_���U��)�Ɖ����/��}�\p�"�͏=�sg�ss1}E�;v�=;3�	)��ҽ�b               NQY��..�!,��#�����eb��t��瞏>X�lλ��gf~�5k�X�宨���ŧ�{-����      <R��k���Z���B_Lg��s�m�{���>�7up����7u��Q�B^��~����e�ܻ�ȯ��`Lj[�S�Xi               N-���Tf0]Hm�3��GN��k��]�޸H���8���7}0ky�K��}���<�1),#��KKN�?�=,      ��d!�b<�_/��s�ۨ�p�X.Ю�j!u�O��>=x����n�ʾ�D���T���e�������p}E���_������-+�$              p�1�/[��z,���t��ct����T���o��Ʉ���{�t�-˳��㮢���tn���.[�K?lT��)uo_     `�X<s������V�9�����k��(27�'��G�������{��G�ͦ�v�۶��FUvi��rvU� ����1              �԰#�����'������Ǉ;����/z!�s�{�t��ʼ�tZ~E���Z�T�$���*���1     x�,�3�5��n� �_�FH=�c���|��>������k������Go{��^��c9i~!e}�~�v����               pj��d��zz"C3O���ۯ���?腀N�շ_z��U_^�^�.���Kv�     ^Z��\_V�����og���*�VQ(GH�sS�G�j��׵����wgTxY�r�On���77���ּ5+��a.�������               ���e��*!uDcQ=6p�ѮK�q����q������?�e���̢�{̍���(�����     �'��<�Pp����u���x��:ǻF�8�>��o�^�{>�`��)��mo���6ߐ��	�+iK�jn               ��OS�RC����#�u7�q�Ͼ*�b/�u�^u�%�?3Ý���4�z&�sA�k�	     �#{D(��9�q�r���z��y�Q�N��\,������Co�o��«�kr���"��3�O�d��ֻ�d�              �E�����ӄ���PCS�T�Y߹�?څW�Ϋ�;"��.�5���]T�C?h}X1�     �{O��P�O��y}���������LF�_s��W��s������gzYg����,ٸ[���%�s2C���              ��-o�����o�:p����}�
�;Wǃ;kn���}���[�<��Z.ж�5:0�       l�>�Ǭ����i�[/�s�.,��n�����'�����k|ZXp��o���9󆯿���-����?M�S���mӏ;�               ���wv������5w^��I����˕c�E9w���B���b��      �֐*�m�����i�b���r-K��U3���\�a�����'$՗?�㫦�~�­w凲��n�s�l&              �H��Ӵ��Z�W�d���CG^��kŤ�$3!��;��ڕ����̥���,\�p ���i     �ί�"����i�[/|��͂��8v�׭�;���?+��Ϋ񭙯�՟U���႐`�9+�,=_=�!              `q�]T.�N�F��5m���_�
����_=��rl�x�����K���Uz��      \������^
�ܬ,�T�Ƌ����E��b1��?���~����}��MU��TZ�U�-X�����%����G              ���%��V��[���߳��	�U߼���+�]Q6����5���9�+s��̈́b     �7b�*��PLT[�ߍݚ�ZE��.&�`ϡ��U?�\��w���1x�6F;�6�$W��9�b               ��@H�T
�y~��阚6ܻo�������7�}Wl���fG��*�*�V)3���و      \F(�/�b�ڢ�;/zv�&�.&��|�y��{���u�U�b���W�	֨�.UI�@]S�              �Ⱛ�Z!�`�g����e��}�gO�X̦}�6<;^���j�`��/�]��u�!     ��\7(__֐���B1Qm�/�/���u�B1�y���?���w���g���?�k�W�V��|:g�f�S��              ��p��-�]�l$c�}��E���+�j��ѝ���k��d3�     �����l\��^��n�[���,�����g?|��u����C���&�4t�,sIX��9K	�               ,��t�(�ya�������Db�s���˺�-��i'��^!X��òa��M	     �U1U�P��^
���	��)� ����}����Q�ַ?�'}_
�y���O�r����e-ײ�<�D�              �Զ3�R!�tmqr�s��`��{o�O��R��o����:�Tf�(<��jg�:����      \�j�U�}5{�/h.����-ݵ�3g
ֻ�����%%;�%+�	�ۑ�N��~V               Hm�0��=�����N����C���v�X�ߥ��	f.	�ϙ�:�b     �����ܨB�97�/V.Ҋ�B�{��=OO�o�o��i!%|�_�8����Pr���}~�[�V�              Hq>�O;
�	������?rѽ7�TH	�~�����K�w>������YXߧ�b1     ��G(�m��;��wRZ��������K���>!��v�����od�{��-
�zM~����fcs              @j��*Qa(G�V����{��|��_�ZH)w_�����C������pCTo�e��i'�:     �"B1.��u'SH(�k����j�����������.9jjޚ��L�LF ]rW�f�I               HM�s3T+<�w���]���R�m���y�Ⱥ蜥�_+xjg~%�     ඕڧ��\1��i�|�}��?M��V�z���on���������}�m�Y�Qذ$�<c>$              ��v����Ѷ���MJ�	�뱎���ۺ�s�
Ϝ^X��q_a     ઠ�T�l�W$"��~��y��x�y�g��}�R!��s����ۃ׿��;�>����ේ               ROf0]�s���LFk�.�{�7�BJۿo���;��_�Y�lN03ɷ2��!g���a��N	     �5i�fI����P�OE�~���LE#�g����}L�����΢o�����g	�X�Y��P���G              ��򚼵
��w�?�������¢`~��wf|�ŧ�"x"��k{~��     �k��,�K�/l�$������H_�������@�-K�3�f���|ڔ�J�               R���Ղw�l���?�UXT�z�O�����wlϯX-xbs�*B1     �mIo��%��b�Vg�h�}�s�Jaѹ�}��B__]�Qt���ܷ)��P              @
ڐ�R����D��H��E�v����쒺�`&��=�1�\      ���qS"S��Y�]� O�Dg�l��w�߷VX��qݿ{�7o�]�~��:.�              ��t�*�Ko<�[{�=}�VX��s݃ǋ���͋���a�uk���o�<57-      �	���ٻ8��:���S����s�ؓ�a$��we�^W���껫��k���꾬CXT\��ADǰ
�����9����sj�0��z����OS�a�j��~�<O=�wfC1�*��0!�B����_�w��	J����%��3=��J�L[j�
�Ob,�              �5��1���L��v������{݊��}`yh^��Q���WW-��&�     �!�xd�x��*�O���PL!L$#����傒��u?�o�;�����Wub}��8q\               P�U�ǽL�k�D�Mw���
J����/���!��Y��[	�      �R/p�G��?�U7{AoM�B��?���^��^AYx~`��5U×/6VuJ�bB1               Ed]�PL!<?q���7=�5AY���ǿ���[��,_.pԺ�E  ��ʷJj<5bx�>��HjDF
 ��4㱾C*�`i�YB��Y�����A��Ӷ'����?,6�?G��^,�-               (��P�r1Tǥ�i9�BPV�c��1��k��#pκ���2\�5�  ��㱎��W�>Yg�#kHee�TUUI1x~�yB1 P����>�dů�	ְ�^/L��������?z뺇Z?�,�8����4               z[l�JO��Y�O{遛v?-(+�����߼ok����=��X�   ��U�U�����1D8� �Cm���#.��@��P��Y=ё��S���}���.�|^���; M�j�O               ��4�"pV"��c�W�RWr�������\�s�Yc�  �Ҳ5�U.�\,�  �b�q�G�����N�7�y���=iAY�u�_�����.�T
�4�L(              �,��b�N{i��ޯ~�ɗe����B�[�Y�j��1K�?   J�ߚ�S  ��y�����0�5�"��ƒәh������]l�E����yj�               @oK���L�3:���2����+wb��4��<   �"`����� ����1�X���ٚ��R�	���T�c��=�������O����
��(              @QXʾOG�����'����n��Ě��n����:  ��qA�� @[�����
������d6%}�ɛe�ᶇ���|wScͥGP[              П}!�_X��㑁�%��xl��խ�$pD��Z�<2��	   ��z�z @s�b��x�T��KC����o����>��] KWb���l�R��J�Tԋ��H�L               �d�q7C����d�i���D`��⟇���
�$�,{';   ��g��Ϲ�  ���o{�UQ�����ݪ|I�Y�����?�[���WN{pY��%ʹ�,
5ʱ�~              ������Qf�~��mg�<�gV��?kj��@���B1   ��c}B� �=C�r߄b�Q���F�3��{n|t� ���oC���
�ZA(              @g���������*���Ϙb^�����     �ң4��8�h��i�@r���Ls�o+���;�9P+               ��=�s,20��-O�(��<x�Ϝ�Ъ��y�����     Pj��b�ޠT��gD'n����H����#[jV�(���               Z#��������	����C�.(G     ��(�Lp�`b"y��������׶�ȭ�|p              �+�0�����KN�� �`l������Z�1��L�      �e�J��9>=�O��0����$o�}����               tU�	������y�cO�O��ǟ|�܇�F[CMA�R>k̳Ǿ�Ԍ      �4(Ŵ&8e$5�-^��?�éӿ�`xmxq�@�&���d̬               @/��qwLOl�Y^Gw|���Pӹ�챏P     @�P�i���KdRID��u�����/�\���i��e0>!               �{ܝ3���� �c49��uC(�-�ye�[      Pԅb��;�#28��-{�R�u��f�n��q@���P              ��Z���x6i���ud��_M4�����      J��PL��Z��prr� o`�g�D�"f�<�@�FX               ��y:�+2<��U{���{��n������jJq~     @iQ���ꍧ"��~���9�];�6��Q�T�7$               ��<�1��+�ILL�_Y��\�Ra��     ()JB1�aH��B��i��F�M��0��ڻV�<�R,�              ���w'L$�?�$L&�OZ7�bc�;     @iQ�	���1��FS���o�I� 'a:���Q.��               Z����%\��pf��Ǭ��(U�%     `�ַ���Y(v�\�K.�d*��$SEm����NR,��m�����|�              ��0���Q����� 'ၛv?}ٷO7C�!P��     ����W�t��=�����x %���1���$-9��y	3�򳈮P�[!               �O�<��OL0���y�e8�     ��l62���������h:v@����֖����/6�	�BaoH               ��
�O|����x��Td@�9�^3����<����$     ���Q��i�z�b�	�8"�I�`�R�q�P�Ba�               ��b�Έ�����L:�cݬ(e��C(     �;�4C�a���ń\�z�L�Y�`*�n�����              �M��=�N�e���h*��9O�c      ��a�|z�C1^���ū��W8�� sM';��-e��� 욘               @^�W�^�L�`���'P��f     0��� �C1n�Z3�x����������(eGb�⒴d               z`��3R��1� �J�����      ��B=�a��bX@Rn&O0Gi3K(�����               ]����h�� s�N�f�      ��f��Q����)	�x��+����Q*��(�5<��               @"	�eͬtF��WƜDf���b�!;A�,x9�     @ØW���f�v�$�u)yX�J2��B�9��@9bY               za�z�l��Ӷ'-�<��p�C�^-�O�c      (w�����LӬ,��\.�C1�֕�f�,�c�2����              ����PUKg�� oBZ2�k�(�     �]6�]n�[�r�\�z,%+=B1�e�$�9˘��r��               z��ߩZ��������	Ũ��b�      ��ܑ;v�����)�43̑�4#�.j�               :q�K�VV��b�d�Lֺ�T!��    �rgƊ>}G>L�JOVX�UΠ���s�@���               �=�`�;���v�d�V1  �`^�<�w뽂�c�f�\:�R�l�e (Iy� �;�cǎ�I�w��p:��`JB1)3-P�-�1w�[B�RY�@               ���$(�7��)��kG��� @9�z��o��-   �����iI$o%�v����|0%��4Hʹ\�b0w.�T
�K�A"              �V�㮞��"��7��kG9bY  �'��#�P�@  (	>�O����b���\|���=ǺY+��f��M{>SIl$�M��n� s�1�j�r|�              �����sy�}�M�<�vc�;  ����JUU�   �����\ozz�����|�;�n�l}��z�z1M���3����}�;�N�nS�T��)�PH�U�|̑+�Y,P�1              @/)"	�y]��]ۛ�v��!N�w���c��st0Ĳ  (/.�K*++  �T�Q�`0(�h�O��=����x<�J$����4�і�2zQ�:6�^y�?�ꪫ���JB13+P+��{�#�˽H���               zI�q�')+�B18i��{�@9.�
 @y�O�6C   JY �x<.v���^i��H$.�d2[��%�h�%��|�ֱY^K4JB1Dԫ�T��Ɯ�ܞ�r\q              @/D��s��Y7��$.��r�q �|؁��'   ����K$���b��oё��}<ߏ�&��r^�G���+���#�$�˻H�T�̊)yz              �-J���>�g� s�s�qc   ���Qr�0  ��t?��#~.������*��$��]�����*O�P�b�L\               ��H�=�N���0!O`�@9�@  ʇ��  �r���O ��꫻���JB1S��@=�ۻɺyH���V���N�               za��3��R� ��/(� @�0MS   ʅ��>>��V�K(��Uxk��:oe�@��4�              �nf�qɚYqz_a��U�+�0Uފ�R��5��  (�tZ   ʅ��>�@`�ꫯ�G�c�	�JpD�7�F����/m_Z�r��$�              ��\(!��7(P��W� �4�k�JM�c�P  (�l6w´ǣ��a   �$�Iё��2}>��T=��P�G4�����U���	�c�              ��d:J(F��@���9����?9(���{.�W��f��� @���bRUU%   �,�J�y:
����k~���,�ٵa�4�0�:��5;�v�m{�U;��Jw���XD              ��T�}��֗���aݽO�7P�q�睨�w  ʏ}Ҵ����  �R��f%��n쵮����_s�5��|%���i��f�R�� R%��#��ԟYw�!����6���D               -KpF�Sq���I�t��c� �<١�4%
  @)I��233������񘕕���ꪫ����R��S���zB�B18	*Z�M�              ��g4��[8	��3�M�c  �S<�d2)�@@�^��\.1C   ����d2�H$r�7���������\q�?q����b�R�2��N�VC |� o���_���
�O�               �3����0X�@���(P?O��x�� �rf�T��  P����̟?�=]tQĩ�U�����p�@�E�����JO�JJ����               �3���W�{��u�Y����x����Y�r����     @�؁�P(t�����|�?w����b�,�;��W����;�q�#���@��#�               @O�q�y:%쪺޺!��T�����q     ���cVTT�X]]�\~��{
��P���q��Ni�U�w�P^��P�
�r���2I              �~���y��x�����L0�     �Y^�����]��WZ[[?��w�k�п'e��j�Y�;W�װs����������wd              �k81)Y3+.�%PkE�y;�v�m{$*������W�k(gZ_C�I     �s����xb����������Vcc�#�\rIB4�,Aq�9�+��]���k���W���ڛ� �              �������4��jU����9�	����:��S��(7��ʍ}      ��0�t(z޺�{����v'��;b�f��r�X�������D^���R�9e�{1)cf�Mm]9�ϸ�*�����e���� ���淄e���T��}_�d�r�}D���.zo��*.I�˥�g|�S��5-i>Sj�z���J �]��9�1*���m;g��٤=1]u�IgOLLS���u-�����#	9r|L�f�u|>�l��"n��?t�+��cD���
����-�;#^��s���H��H�j��qd��>��1C����PR��=�4���[��e�дtt�H"�q�JK�Is�_뵧d*-��cȑ1旪��V3-��"��c����R�u��$\钀���h,%G�Ge|�cH�����������@��O](~���ˉɸ���ǐ*���~u�����!ۿ�#�G�o��'��9c�5�����C#3r�{Z�q��ί�-A��i{o�56�0�T��g�{����̞�	9�ɭIB�5+����e���/c��u�0*cz�{JAQ�/���e/���3'���z{;�����	a�y      ��0��Ν;�JQ��#1v,�9P#Poq�����]�߻���/p�`bB�����q�j���i��ʎ���,;g���A��c266�e,Ǝ�$�Q�z�G���R���-c1v$��XL��r������>I&bZ�b�HL6���N�d��fٻ�S�X��LBF���'�{�*�ϧk����cH��.9��&$�M�r�X��'�ّ���)�u��B9�=�\e�/k����Ǻ���268a��ZI��284�e,Ǝ�Dcɚ��y���s�Z�O�r�Ɏ�t�Z����v�|���h$�e,Ǝ�d2���M����R�ɖM����ů��|v$�w`�z������N_&O?�n��yB��k6�������.���G{��_ڑ���	֥`/C�����_�2c���uq��-5�r��?0�e,fp$"3�1���VK��ކ_��4�_ڑ���!��Zp��-�?8.3�-c1����L�~��kB%��-gnY.�<w���_ڑ����9㴥�܋bf��_�w��z��t2��tb�:�p��n�8����pJ�ߺ�m5�*,8��       ��<�&���@EY(��!��y���u�������V����鋎
^����23�q{��v�`;fͪ9xؔ�I�b1}�Db�V���3V����*3����[*[Nm��^��.�I$�qu�!�pJ�v�;38<n��c,&����c2B
�9�sKrG�����ĸ���p�1\.-c1v$�h�u�)�NZ��)w�[,f6chxQ��YǍ:�bf#1�)	�S6��H^�߭],��w<��s��*d����k����0�t��y�����b�HP8������B�b1����qY�:�b�����a�}"k;�lIc�V�X���L.���9�ކ�k��#1ǻ���i�-��z�����"1Q"1
}rƖ��bf#1�/��uˉ���:��n�'�7�~O��������u�o�����o��kC��<     P��<�ȳ�"��{ll̓�dr�UVVf���S'q�b�;�L4�4�>3([jV�s.ir�}κ{� �+�8%���cڣ��7�[,Ǝ��7Ry�4SkW͓��E��'ť�����)�'��BE�/�y�٣��P��KDb
K�X����)�b1��W�+eI�X̫#1p޼����%cGb&����n��WGb�<�b1��3Db
D�X̫#1p��y��N����_��MJ&C.��U�b1Db
K�X��.�$N�+�b1Db
G�X��"1�=�n�;35C$�t���.S�q���b��g���`Gb����t���)��[�j�ig~9'��tֲ����P^eYռ+�i�     @��?-���2����Dno��{ �����I}}�=f�hLi(�#�"���U/ڶ�m�gO�>遄�U�����#`��&�e2�]b1l�҃.�;��)$;s�酏��у.�"1��K,�H�t������N"1�f�b�Y����޳7����"1��/]b1Db��K,fpdFf���WH��bR�,�l�تE,Ǝ�$�1A����DS�7H$��r��g�����X�D$F�`M��%31��s��wʖ.��\$�c�z�`~YH��bG��%�����6���˧�4��=���韐D2F$��t���у.�;c2���	�Z^�x�����ͻ%({���U����!�     ��������v@&�L���b�4�>�"���՞�͡O��UP���Z�8���9+t,��H��F*m:�78%��:�H����H�&
����,�-:3!��B�bf#1�A$F���n��#1c������X��~uX��ؑ�c���/5Q�XL.�$>:cGb�{X{�E�c1�}�J��W�XL.3D$Fg�����"1�(t,&�%����b�������W$�E$F����ч����b~�kk~p�@�H�^
�!��B�b���б��n"1o�PbR"�����z��� T�9���e�����.���DӉܘ     P����������������QNY\�q!S�v����5����oN�b1٬�F**C$F?���ؑ��^����B�b���P��H4)��l��L!b1�HLǈ."1:)T,�H�~�X�;���ĸ9��J�b1���2�06h�P�"1z*T,�H�~
��ƒҗ{oh�P�"1�)T,�H�~N�bV:�!��B�b�F#Db4c�b�~�*�c1Db�T�XLO�$���b1�-�g�?�h,�H��
���6�&��7�4M��)�V�3N�Yv·������w	����ְ�f��Ǵ�sc     @9z�u�b_3Q�Ie����P����뮽�����ǿ!([K-�gS���#��7��X��9�9�F*M9��'�-�c1Db��t,��w�H������D���I|�r2���t�єӱ;3:a�
4�t,&kf�X��M9�!�/�c1v$��{X<�9�����Lq��fc1Ͽ�n7��HL� R]ٱ�_=}�:�wf�G$F_N�b&��22F$FGN�b�����X��xD�g��_j��XL�H���X̾}25=��ކށ)旚
����b����D,渘g�|\ �k'�Jw��lT}ɺ�A�Z`��S�	rP���     �$��[{t�P�Ö[�޺!S��j��-k��8�#��
�b1'��N$Fw�X�!��	��;#�5�b1�TZ�zFģ��o�S�;��$�r*C$�88���H�A$Fgv,&wտ���"1�s*���t؛�9�OgN�b���ϩX�l$�M$FkN�b��'%ɕ޵f�bN۴Ty,&�HI��'�i+�Ŵ�ўS�;3<6A$FcN�b���b1�c��&�3;�6{]��#P8�$S֯�/���XL���$��mЙS�"1�a�e��b���tކ���]�����W���ζ�M5K�#pTG�=�      �H}(&2(�7���zɒ��_t��ѣ���<������NʘY��ձ���A��^$֮V����h<�&�"0�y��c�l�#1��#�&ST�b:{�%�%ST�b��������Î]Uo����[U�"1��b1�yX�����).�c1C#3Db���X���:s"%ST�b�HLw�('�	ձ;c�)
�c1�3q�c��T�bNDb���	ձ"1����X�˕�b1���6ձ;�8EAu,&�$SLT�b:���M��5j���5wXw�����]��jv�9�xd@      Pz�/���8�e�dyx�.�n���\�낳6W/?E�(���T6-x��X�9g����u�������HUd�X��/�%���|�4%#SL�X̺5��;��3z�F��;��s�bJ~ǆH4A$��ر��E-242����� Sd�X�S����xot4B$��ر���D"��8?<6%6`;��sV�s/��c��M�)2v,fz&&�T�7�O�̈�ㆢa�b6m\"G���s�ޞ1"1EƎ�<�B�d�O���&F$��ر��K��0���ށaN�+2v,�ik~i�{~9%Sd�X��d�LLM�����'����K���|��^.֞�����IJ"��cONN�*"v,f˩K��ូ?vW�8{���yd��=��f�Db���Y�r������{���\,���b��<az���@$&_�E$mf��3:���u���>���{fecgێ��e���Q�EP�      �&�ž2ݓ[`��%p���%�w~�ݗ���������_�8��i����c�b���_��3�������d�l�$S�<^5c����ɽ_�S*E�����M���Wܮ�n�wO�j(F�IA���旼��Ϛ_zU�x=���%~ǎ�\��A6����Q26�&��(������i>+/Fn����؟3�Q{���ؐ��8��uY�
����Q����P�|^���>f&C����n�!�_��y���DH�)�I��YU�@��z_س�]{�u�hH	��h�W���aǣ��p�4     �R�|��^Xj����y��׆�%�Xw	Ŕ������͵�V	��S               P<Lw�)�3�V�;���7����k�8�ukݪ��w     ���H�y�t��XY9��cw���ۯ�ӂ��!��n������S              {��{�-pV�7�Zh�w���(��*o��`�d�      �49�90�%U��kW~��۶�Ӄ������~�m+*��7���}              �x�CEa�Y��o�p��?��nAɺ��^rz��͂����     @ir,��h��xV�<j�=WP���s���jWTP��               ��hbJ��~k��<�[N�]���m�ַ��e%��{u���?d�]�y��6��      �&GB1C�I�����]��k�|����oJ��ݵ�*V��P              @q���65�)���j��=��u�
Aəny顳*7�

�=�      �͑P�m�t�l�o8�m������v|�޶G���qÝ�~bK��5��90�":              @1�c
�j�((�s������_z��'�����ؾ�܆����`�      �6�B1/N�m�b
�5��^8�ۺ�6AI���Z�mX���a
c2��3              �����1A������'"muM�=��mm�<����0h��

�q�6     �R�X(�ٱ#b���(�s�ם{�]�ܲ���n�U��?��U9�3�?���Q1�/               ��ب���d^�NP+*�W����u�RA�;{~�VU.��@|\z�     ���Xdb$9%�!Yj�a}�[w��f�H<�՛�<,(Z����=��z�bAA=;~D               P��?"UP8okXw�G��껯��Ek��\{nú���8��      �:�B16;�@(���}U�ӫW<k�ky��ᤠ�\��K��ָ�C��2��&�	               �׳c�b
�c��u�5~[��oy�EAѹ���ok<�n�����C     (u��b�����&(�U�j�N�̺{���\���k�Ѵ�_�.Gt�'�TD               P�^�l�������B��U��4,��<����U{₢q���z����WE%��Rٴ�<�!      (m��f��H&.!w@PX�֭=�{�{�m�}�:AQ��m5g4�x��f]v�
               �-�Mɾ�N9�f���VVί���h�]#(���YY��FPp{�:%�I
      J��������&������2C�oܴ3qg�Ȯ��@kmmm.M��C-a��%              P�}��b�pz���}��?���_&����w�cg֮� �{�     ʃ����c��h�c������Kޑ>r�M?��@[��C��\�v�@����               ?{��Υ��a[��Kw'��_>������]v�;��_,��o�      J�㡘�=(]�#)A�<ƅM��C���q��O<&�Χ���'ή_{�@��/Y3+               (~��Q9�e�A���M�o���N��_�ܸ�O_ؼ����`�a=�     @�s<3��ɋ���ڕ=T{��w�l�~���/���_
��{��[�lZ�@+?�'               (?�G(F#��i/j��?�wH�Λ~�wm�p祟�������?��g��q     (Y���	���v��r�O�;�w��O

�w��7�k�x�@+��?�%               (?�+��|1C�;��e�K2w������.����S?�#��_��     (Y����A���BAZ/����¦�v�w~���+(�����Ƕ�o�X�;t�5�              ������~YY9_���+�l�{�.W�n����Mw^ֶ���������^鋍	      �CAV�f�qy~�l�[-�K�7�:��w�������Q�ڶy�-���Y�k������              ��c_P�P�~<�[.j��)�=��ۮ��u��r�{�9�q�N�����({�     �I�R��":�=U{��w���U�.��;n��g�����7����Z�l�@K#�)90�%P+�HI4�����^I&E&�LK&���C�1\.1�YA�'�JƆ��_b񔠸$�3���̚.럆�m
�GR��೎ҩ��x��I���B~�=���`24���Z���^�d�7Uǐ�O�񨠸$)I���zp�ݒ����j%��旑(�O��~=�{��^�2��H��Ȣ�L�Y�������x�fV���/����5.���G2�T��d�/��/�I*��^)�������׋Q�z=$����!k��q�N<�n�ɾ��=��f����n��PL������+�$���w������/֞����^���B���%�7��W�j_�����x�tȧ�~��׸�}�\��~_���     @�(خ��FI�L��`㋎n�\�r������~n翿O���r�Ƴ��ri��J������Ǖ��R��9,-���Qhn���G\261.(�_���
%��-�W�vI�XLQ�����䌒����R^>�+3�iAqػ�GZ�J��vI{W��)�SbfRJƆ������SIb1���d���Z���cۯ/��-���b�DG稄*������
�����d���Lf���~%��c�r�%#cc���ʑA����a���v����.b1Ebz&!#���֞���#S��/������\R��~�K�t�p�N���T"�dlh�Y��.�ŉ�{~��^%�K�^_^�[:{�9ɬHt��Y�!!cCM�B^>�e�[X{*v$�C}2�I����1��^4*(G�Im�W��/�����W�$�%Pf�	S6���������8�;�'Muj�6�=9t���Ebd,"�XL���XW)/�h,"�߉�������'��%���=)4���C3���j�@?���;ֿ�yϱ�W޶��o�3!P��3�YU���i5˗�e�Y�q~   �B�d�=�G���C��1���:����}��+*Ԭ# �W�*-�L\~5zP�5l�ɾ"�y���[�@�c_��̯]�{H�w�����/����&i�ɡ�ؑ�c�����:���z��9xD��;ST7,��TȚ����n1���tfGbF%X�U��.kpظn��t�G"����HLu���	ۂ�p�X���H��tD|>��Ƿ� �Ni�Ɔ.I$�j��Nl�������?k��Z1�Y�"�9;cf��v�9�2�ʆ���� ��ّ��G�$\�W�kV4ˡc����btgGb*|���p@֭ZL,�ؑ���a	խ=�_�@^>�#3�/�gGb��Ԭ5ؚr����b������_�Z���t�by9w2_T���HLm��c�����F,Fv$&�L�ǣf��s6��Ɔ��d~���HLuX�ذzyS�Xrh�X���H��c*�Õ~9e�bb1E IHWװT��/�, S$�HL8�noC}]PV�"b1E��Č���K5ǐ�g��-"Sf#1��*�6T�a}�w����Џ�^$�9;\���������v�\�wW�y�[���di�YAY����   �0����������~/3��o����G  ����)��PL�T���>Z��C�s�M���E[[�+:�7��p��=����?�gz�Xd@���H̬�X́#Y�����+}RY��%�Y�P^9�C,FS'"1c�"1��X̦u��hNu$f����/�w�ѕ�H̬\,f�bb1s"3k��z���詣Km$f�}\b�b^>�!�4'��Ȏ�:��$�Y��5K&+26N,FW�H��P���Y�r��r�;we�Gu$f��e�Ƶ�ek~9e~�+Ց�Yv,�4��vb1��(��̲c1���wK,N,FG���~g�v,ƚ^JW�]�􍟈ĸծ=�b1�X��bt�D$f֪eM�@��(�]���̲c1��,����$�a�IGv$�Sa$f���:3ˎŬ�Er�X��TGbf��b^<�%1b�Zr"3k~K8����X�2?zY�]�]n��x�+j��?��~���'A�ܸ�ҿ�ְ�﫼.��ٔ��+    �w����7�yR{����������햚��\8f���A���	 �+h(楩v鍏ʂ@�@o����;������M�\���k��zV��AQ�a��5r����rf�bo�Z�r�<l���@/�K��#N폯�����Qb1��]$ƙ���X����e&�շt���^��rnak~s8������U�q*3�w��nI$b}8�����.wK,F?�HLF}$f��ٸv	�9���b�+������M0�ԍ�	8��U[]!kV�ёS��Y�X�:b1��kCV���_67T�a.�#�btcGbF�&�Gbfٱ���|��$��R+��f.vn~ٺ�6wK,F?v$&��+���
<�~m��=�%�tR��t:#_�מV/o���яS��YU�~ٰ�X������"�7�"1���?��cݒ5���dԡH�,���S�-&�!'#1��b1�t�b1�<�d���ra�f����e-g�c��5<{��?�C�ނ�m;�*{{�)�4���b���}�1   ��&&&����v^��{GGGs�JEE��c^����  �SAC1�ƻ</W/�P�?��+�7o|_������=x�Gsv���Ϸ7���xC֋D,��=#��O8���;�o�<9`�b�̧�W�K0��禹U�b�29���	�"1��XL���{$�d>]��Ĩ���Z�R��%���!g#1�r�����@,F���̲c1�aJ���@NGbfٱ�k���W�$��|Z�Eb�8����_��'��%�}8��e�b֮\l����h��H̬\,攅��@�L3�Ԇӑ�YM��bʉXg����H�,����)�]�k>{4��c1��R:{�����H̬��r�bb1�#1:��e�b�a�X�6���̲c1�����N�d�_� KJGװT����@,F?�_q63��ې�.���=��JPx�1������g��O!"1��T���/����R���%S$���ֺ՛��*�������	��;��8�f���8����    �{��G%�H8�\�X,�����G���zsјW�c����v�3p �s
��=1�\�z�x�l����%���5�S��/\��Nʇ��}�P�׬X�r��g�{%�q栽�ؑ��G���̲׭l�}��2���w'�q�g���*�lm�e��歽t�$!�sg��d2� 	�;���\Ba0!��Y +�,$���ֱ,��h�w��U�JK-���9B-�ݒU�9U��>o�Jǖ���S�=�}��2��MCb\i���肪���UѤ!1S����h�b�����D�Bb,��q�L�-���)Z!1����+�v�loQ�M�YND���r��P��C��4a1�v?$f[����Ú��a1U����NHLvdCb,�� K�����NH�%/'݄�t����E��Č��IVFt�=i鹆
��9!�k+��VH���8+�_�b� Z!1�����t���a1�d����F�RUU�K AJ�qh��h��Xv�b����m��͐˙S%~��/�+Z!1���4�?s��А���i�VXL[��2k�NCb�3��䲴(St~IXL�-��eff1�!1������0���h��X*���<wd�0�P�Z���9�Y"p���bW���e�Ͽ>�q��_�'P�s���|"��S�^^�C��I��    �������;��ޖ��i3��r�v�ctX�2��Œ��-  ����ŭUi^�'
Α��Jx]ɥ7���m�c��o����
���w�3q���_�����s�3�S��#��4I����o:[&��	�^q����d�G/$�RX�!g����(�vH��t~�+�;]c��N��h�vH���X��LXL��ĤD7\4-5I.֟��]#��D�?��D���r�D�$H@&�g�����4�UJ[����y���ݐ����c�����%At���Ԅ�/��S)]}c��D����ep_<�PNXL��uD7$Ƣa1-�#,&j��c1a1���D���'���g�b�'�!1����.�b��!1���J�1an���h��nH�E�b�TIa�Q��lG5$Ƣ�⹳��D[�Cb,�(7a�ܿ�����^H�E�b.4����D�Bb,U:��a��M
a1������5?(pm^�=E���X��y_����}�O/���C�ו���/wF�b�K�Z9'   ���ݻ�9�x<fLNN>�mw����������: �\��\�^��IP�C��T�f�?s�Ew�7f����"�w��?����$w��_�u�h=�^���qA��%$�b�b�4,& �TE����D�˼Q�b�H��qv	��h����J��9&a1�v�cL���@�b��0a1g��KZZ2a1Qb�">K͉��!A��g�e��KVF����������Ґ�����Xt^SW{\��daiQYv	���纤�T�t0��4��~H��
���9.kk���2!16���iX��\F&�Ϙ_F�	���~H�E�b��Wʝ����D�����&��qh�0���X2ҿ�9"��mA��)$�Rw�T��	���II
�f~���n�b:	��8��AH�e',�[d��g��K��/*����H�KH�%Y�6v
��T���221|f�s�X����'_/�	�y���������I퇏�������_���;��篽z6���sO�$P��Hހ/x��#    "ohhHb��Bd���$''g'D&//o'D���HRS�s] �-�Z�\�Iς��
Σ����pv�b�诲?5���3O�җ�zE�[��?P�y��.䜬�⹳}~� t�cїiS]��w'8nAd�-$�RT��o��h��-#���UH�E��/6T���QY][D��Bb,��r�g�Ad�-$�b����g��c��ԉB���Ԭ 2F����6��$+3̈́Ŵ�豁 �H�[H�E�7��Ǥ�Odj�b�H����T��/�3��t�t�뱁�e$�-$Ƣa1*�Ŭ�"�n!1�������(��H�[H�E�O����旑�����"�|��'����%[��X�Ŝ�����3��"���tO�*$Ƣa1="���_F��Bb,y��bD#��
��ל����Y���!R�c)-ʒ�@��� +R4$��6Xa1w;�dy��a�_޳UH��*8�$�=5旡�����g������Ԑ]Uz:�칲�.�1�1��?��_�8��?{�jWɇ��~<5�^�i8��϶�{��~    ���%��|>Y\\4cpp���YYY;!2V���X� ��w0��OO>/�x�Ε����ڒ?>����U��G�����o.�Z����^��S�eu1���{������WgnBû퓶�	�t���=� VW�{E�:�qn�sR��&k{-��������b��`'�<�208m���zl8u�T�n]\�!����&L̮�Bn�K

dd|F^K��woIRS�dk۞��k���삆��s����ֈdf���PZ�++k[2A�N��̮JR��$��2p!!QNT��Y��������i�cCUy�,�n��nã�R\��=痩��R~�4�>1!z%᳹�ޞ)I��SU%����uAxu����4������HƧ�qh�յM�3��U�^{:&�}GB�zi�����,Y]͗��9Ax-,��+5A���~�=_{'+��̼�/������r뎽����Ž��Aqݫ'"�&��0C��9�LNN���R�7��2�4���k\2l|]ڬmXfmC$��kD�m����49V\,SB������HZ�}�'�J��K�6D­;㶞_��k�/C�S����J.
�#�+51Y�Ya��K��.z~la�?|�W��8�~��OU�<y%���i����i>5�m   y[[[��rwuuՌ����%''Kvv�NxL^^�N�Lqq���\
 �`�����[������f'���қ����]��K�9�8��X���s��w2��o�ϭ�I" &f|~�l��y3׉��Ve�q���x�ƈ jxt�@=��� ��g�@��p�m"mȢ{C��-�����1������w�P=��f �k�@�n�dum��%v4�0.��7�b��y���o`x�@1��?�k���Ҁ\�?-p6Hyea�y[�����k�3��~����e�a?�ǯ{eEF��_̯y<#)����Ǥ�5�  �h���<��,..�18��kiě���"c�X���� p0�	���o���OV�J�R3����U�}�?P�1�1���~��?&1��������,��S��r1Eb4(               ��S�&(&��'�������y��T�d�����_ṱ���w>-�_��W'7�d�JuF��r��i�{>=�    �YZZ2ch���.��E�1yyy;�2�X�f  ��&(F��T��h���`�?�H�ׯ�i�*g>z�����[������o~��)��w�3�^�-O/�ņܪ�L��c��ӷŽ�&               �_�܃2�vOj2�	bGbB��˭.����������|{z������,��?�K��Ն��W��P���֦���    ��J����199�����$���1�1��1V�LQQ����
 �[] \�Z�g����,�M'2J2�����s�çF=3_����ч����bSo�����3�XZ�O�f�^zE�+�1-���$I�               �N�]z�y���-�M�����W�����W��g=�kSߚ�v����+������gAr�/�d��*W�K�>5�msL   �D�����E3��r�v�cth���X���kl��"�J��4��LvyAp�)��M��T����읅��/������ۿ2�?������yNZֿ=����S���3���!�������               ��L��T��0-G�*]E��x}���_��󾡵��٭�/��?��_x�V4�lo���]�J�xsqj���,�-L͡j��\6�"    ��<����lKNN���l��1cʔ���� �4�;r�������gu��Q�Q��>��o=�T�ƽͅ�����+��oz�/|��	��}�;_�\S����I�o�Jr]-J�n��()�Nq%
��'ƾ)               ��|�����N�� ~hKpha�����O\�ύ/m�u�z=�^���ғ��Wo��g�彯���������ߓ���X�^TY��k��D���X    8��+���f>���r���a�ʤ�� ؑ-/���3򊂳��@�����4���������ѻ����_�z�6�����z�|	�Y����߿��$JRVR�d$$$&$&%O$�$&��&��RRJ��\�rS�r�Rs�Rm�2@��X��1               ,�{�E~��	)L�ħ�Ԝ��>��C���ɫ���Ս孵�U�gzÿ=���No������>�V�7��N�%���yRrbqb �8-1�XJbrizb��dWiNJF~aZvzfR:��1��b�A    �+8����c�����v������32�c�	 �b˄���{�N�ޢF,y�����%�|zB��g               �m˿-������	`�@�LW�K\E��Ӳ�$@�}<x��c   ��"$�<,D&))IrrrLh���hp�(STT$��� �bˠ�����Da�$&$
 D�w��wuB               ���x�U~��	)M� ���M�|y��     ����������lw�\;�1:4HFe��8
��Lx�幹v���� ��#��
               �o�'������ ����>'�~�     ����199�����d���6�1��1V�LII�� c��GF��W5IRB� @8}c�C��	               �R�2}K~��{�xz� @8Mo,�Wgn    {HII �^�,..�188��m������cdtX2V�Lzz� ���b&=���myC�c ���婱g               xo�'{N�s� 'm���    ����l�b�����/KKKf��Q.�k'<F���X�2�8!!A �>[Ũ�F������DR� �������
               �r�6sG~��{�:�T  ��g�ٻ   �^���eaaA�h�x<fLNN>�MÌv���Bdt�v �����M���ķ单� 5�oS>4�5               ���_~I�}�- ����/�/x�   `/�������^���Κ���������� }���  ���A1�cߔח\���\�P����eakE               ������,t�?+� �����R�    ��'Nȝ;wp"��c�����RSSMh��Ck�����D`����o˓�_�_9�c �2��(���.               �a���/ɕ�Ӓ��e� �����"    쩡�A���/��֖ �D��{����l)..�	��&���. "�1W���k�:~UsN ��ޜ��{ũ6S6%m;M�����)Y*`õ!�[ɒ�s�)�%Aĝ���|IHHķ���Y͑� ɽ�Ο��ՌU�Y�`)gI
�o�O�;_�O�S�%}���r��h�H O���-S|)�8<UX�^��bV]�������~�3ݒ��/�r���/�KB��e��%�d3mS2<赧�E�s�I�A�l3�����/�����5�$� ��������sq*mZ�����c� ��L|G&6�   �=i ���祵�U�x���b�����222vd������=�T���/ʟ^�y�� �m��|g�[���|�\m�*�-� ~��蕩�)Y�^����k-}MZ�Z$5�*�گI��1�y1]Hu��]Y�]�ӣ��b�B����Ι;���)��.K��b�x�O�Kk}�Yx{�����k�hҜG�~p���Y�7�+7�n�V�\�*��LA�(��ccR�Yn�#96�/�iil����^{J�T�4���d����ɩ�SR9S)�_Z��B����n�(�_Bz��-Y�\���z)],įقY�^���+{.�4����E6�7�J��Z�į��2X6(��R7T��2�m�l�kO���%m��e�
zN��T�TOUK�d� ~�\�f�MI��ʵ�6�3�������]?\/%s%
�1���K'{j������ 5[ �(�����c�    ���׾V:::��� ���u3���ؖ��$999;�1&c�Ijj� 8<G�e�_���g���K.
 <*_�/9�%q:���r�E��_��M:�ŝ���.�.�6O�K���ڱZ[ơ5ך�4���[����S��v/�R�U��k�ŧ��9i?�nk�ԍ�r��$���7���f�MYO[7�k�A
݅��������M�Z�]��go˅�& �E�9774�7�k���䕮+��N1_<�;�'E��D�	��/>����F�ѷ�������r��e��B�*ė죘/NY!�j#mÄI��a1�&��[u�dŵb�w�tI`( ����!�ׂo��tKk]�\�,���fw��}A���V��E�=��R5]0m��0ܠg�R1W����ҵI#�x��=o�ɛ1χ��7�K#�8e��*=w�s�ħ�!�������,�-ğ{E�������)�oS><������R �(>8�UY�m    {s�\��?����O~Rn����dqqь���m�5G���&@�
���d�sF���Kq���}Y���Jn
�<��L|G�צ%h��.���yE�<�ŋ�ݜw�,�4;�ŗ��,���b���w!��b��dus�M��4,�b������nm�����Ǝ��nλ���r�����	�ij6獻�ַʥ�K���+���9�F1_|ZM_�ֆ�}M���M�N�f� >�!�P��v��Z6R7̹�^{J��y���z�����}�[��~)���/�����@�������f�j/w]�D?a1�bo�E�i����w� ~�qA�[�6S0c4�����cw�E�6�s�Ϋ��a�W�0kNw�\��6X�pΌ�ď��%�]{�E_�J�N<�Bj��5sϊ�
A��*������x���1� ���^��L�    ����(KKK���O<"}�,//�1<<�����������͕�D֨ ~9.(fy{]�z�+�k�� �aMo,�Sc�J��"�˝�%ۓ-�q	"�\He�)�jľ�Bb,�ŗ�ZHe�b>-�;9qR�vwsދb��b�97�S7���?�vs��t~��n�w��b���h����y�[gnQ�'L7�]2�?��v����rFp~Y����
*��qU\t~�u/Bj��/����JGMǾ�t�a��ۘ_��;�l�)���n��5מʧ��M�!un�s������k׺�I���e��J�2�{CH-wO�5�Bw� ��T?BjY�]��3����DPq�/�t�����uE��i������CH-4/���Zh�_^*���_�/��T߫�6}�?6.�K���}���=�6IMp�} Q����>k�%    ��'�0a����essS �����ݻg�^III������� +P&55U�X�ȫ�_��%�.>'���Z	�p�����ےX�])�m/��y/����|޼��j{诡�/>��B*�ȱ�%���(�бl�x�tZ{��O������� ^���^�3_�_*f������ךkMn��4����b�Fچ)�|���)��;'����*��YCH���봘����r��"�|1�a!�����Y�v]��u:�Ǫ�!�P�Bj���VPq�67�c�^O���V����U��vҶTOVb��C���c�;��t�?I�^.���v�M��d�D8o�E&���CH-���r�lp~���2�d~���֥�K���+�M���v�mqg������
Į���Zh�^.�Ԣ��g�F8��a!�N7������5 ��ѯ����    p���&�����^:;;eaaA ����3�7��^o���|Qx��XGvv6��x��
԰�����Jb�)��ѐ��K�˴������rݜ��b��ڶ�a1,��9s�s�^�.A1_l;�B*�x�l'lK��|���9��|��]��/F�n�7^6$��_�o�ҙ/6=���^��{���I1_,�ߖ��� �|�b���rݜ�҂��b��w��9���ȕ�+��F��Xs�R����a�A{Bjѹ�����x�㒶E��X���D���1||�NNR���*�d�d�@�VCD��5˵��c�ACb,]'�L�o�\)��s�R�;�-�u�r����XtА˭3�X����!�8���_j�����z`A�9H��F8�MCH[�Zd#y�@�~�lD|)4Ez��t}C,���7�E�R�Q" pc25�-   �\�׽Ό��UY\\���%q��|��:�: G���f����Mw�������yyyf;`w��K�7��#���Ϟ|� ��Y�^������ij��bAl8h7�r�����b�Xr��t��>�/�v!�e�h��ә/v���^Z�g[�_��m��b�au,t�A�ӿΓ�/��y/����<o�"�~�^6�8y����)�~��S�+�XoBb�c1�|��r��b�Xr��ݴ�S���V�����6ܔ�����Xf
fL��	*&�4&���1�8\7g�h ��/]���
����ACH-#�GėL1_��ꑩ⃅�Z�>�t�;Bj��6�3��`BHO痹��_�e��sO3��3���!��'�hH�^����ah#�h�[Bj�Nl:l�E��>Q;Z˵�2P1 ����������?#�	��x8�c�Q�ge��k�    �+++ˌ���}�{<&���"&@F�e��}��������Y3��r�^ ��1V��>fm=���+�>3�yUQ���. x�?�������:NvHCB��s��p��漗;�-/�}A�y�U1@���GE1_�xԅT�̧A3MMt�CC2Zz�n�{iXL��f��vU\[�9�'�c>c�3_�0ݜ�s x&p��:�ǈ�vsޫ��w��f)�s��vs�k�u�����$)�$p.����Z���n��M1_�x�R��նQ�#4�TC$�)�k
�/;�J��b>��L�4ř�:��b>��h1.xh��Å�X�������&,&u;U�l:'hihy���_�/�$�TMU	��QCH-8t��\�&�>�f��QCH-R?X/���g{�R���B�I�N��!���'v<j�E���U�Pa11��Dp~Y�h�K'�Y��߻!���+ ����c���~   p&��Q\\,555l� �����P�X�F�~�crr�m��ɒ��mBc4<F_�:�ynn�$&r����j�/�����Ʌ�()���_F�Y薯ϵI���3Ig�l�L�LG]HeY�\�ֆV:�9�.�?6.�G�^�9�QRY�r��w�����蓉��#}-�k9�"WگH�f������^t�s>S�s��ݜ���-�� �4o����r��v��#���~�oU�T
��Q�9�e�o[L@�����W|�,�?*��w��P�LG!�P����ر�#��uE��)�s�ʹMinx���D�9�P��\G!�hP���\m�/��_:�QCH-�e���R=Q-p&Bz����xi&,�j�K�2!����}��CH-]5]
H�|)�pJ��Z�Z9�Ԣ�p���1�O#u���c�=��h��|�)�f.�s���F8:?in��C鿟�3h�y�yr�i��V��� �gjc1x���    �nB��:����|����&c���ssss��u�5a ^��9Y�����IJJ����������׳>OOO T��2�6-O�|M~�� �Z�^�?���W������|�\�,G�漗�ַ�"�b�G�tˏ���B1�s���^���,�|����n[��鶥� �H�J���P��4�������Gg>�2!1�we1�h!1]��AR�:�I��ߝFC��O?z7�*ė���j��������~�R�����(�s��<Pq�RK��6�������Fu4�!����-!���u�K=�$w5W�,�u�QwCBu�H��t~�4�D1����:̼"t~�|�ل���\gY�^2�p�2|lX�	^9=~Z�,�Āܪ�%+����X6R7��\�	�J��%T!����&l�b�B�,&���!�w���).w�ǉBBj��s���6�	�چ���>�k]��,&����!�N��m��v���ᅟ��� x1_�/�����bS    �04�";;ی���}����	�X]]}Q���ll��f��i��K��(�˵�C�d4@�z�Z\��bԧ'���y5r5�V ������Y�Z�x�W�'ۉ�R=U-p�Pus�K�u���CKh@L(RYL1�P���S������|Σ��9�7�����*��.K�z��B��y/:�9O��9屢����.�گI�&��N����:C�}���}�b>��'��f�MYOMH���5Q��$���RKWu�	$*�-8�	�	�����y/S���9�|����ܔb>g	uH�E�FK1���:�ԢA�Fz���dlf�a>o^�N��������kg���A�MhpC�BH-z?��_�doL,a�y:�?6n� B���_h�� ��ۦ�E�BH-k�5||�38�0�t�P��Zh��<6��tJ�&��bk���/O痹��_:M��||��� �����K��    @8h���
��z�;�1���d��t�s��Z�crr�m���cBc4<F�c�@���"IM��/^,&VY���}V����%'�Ee ����w�e�W 2\6ln���<)��Pws����w��ŖN�]�u�t�t��2})泿p�X����ۖvs�_�-]xK1�3�+$�Bg>�u7�t!�.���A����N�{�C��y/���c��sjhCH-V1��6�b�N�!�ˇe��H�~FoU�96T�����B��y���53���y�b>�3!�'�d&?�!�-�c~�8y��fؾ?�|��ҝ������Ody��6�?'�5�a���%��K�I�PמlN�!o6�>�Բ���T����6�W��4�Iږ��j��m�l�kO�Z۠�K�4�p�O�I�#��B#�Р�����}w�[n��M#W�Si�cy��!�J @i@�     Z���w(jjjؾ;HfuuU���Mx������n����Y��+��g^_:�'��O��V��h����'f*��V��?'�^�� #k3�����d���Ylyz���v�n�{i1�.��3���n�E�[He����vR�������X�c�`��i��3�YHE1������^Z��~�]���XliS������	~hgث�W%ӓ)����Is~����|�>���Ϯ���y/-�k>�L1��U�hI���W��k����d�97�/$Ƣ�%��[$BH-:������R�=�;��B1�������������*�;/K�'[`O���I������i��0� �'m8���"�a�9&�T�!ۯJ�v��~���1n�Ǉ�ϣ�}m�l��l��v���"W:�H���vdBHk�BjѰS�(�+%,Ʀ�Bj�i��u��b�
w��~���O��.�M2�9��Ƿ%����96    �]��y)�g'�B��h�����9��
O�C ^�kN������5���m^�%%%RTT�"���+��\O�E1u���.���M���� ~m���޿�-����Ƌ��"����^���y/:�ٗ�Fu��t�t�~&�|���T�̧�-5�b>{1ݶ4$&+rݶ���q�Q����n�{�g�S�gS��漟����}E����n'z9~l\�"�3��j��.���pws�K�כ����K�����G���Bj.6�'�(�3߫�E�u5�k�k�M$CH-Z4
H�<�|v����3w"��(泯H���v�ᦹ֐��'�=���H�)�o�W�������迋Ah������R�H5,Ƶ�؋�����?$�B#��z���H�m0k)��`~iC�!�tWw��'��O�BH-�N�p�(��[u�	!u�{��/�/��k��t��2�1/    �t.�ˌ���}�[A2������l�dv��v ���zw^[���/ږ��$999&4F�c���v��
%-���NswO�j�Kr.�T��@|z��?��Z��f�x�,����]D:$�Bg>�1�j:L @�i1�$�TOT�!��,�a��|�b�m�B���/��8�!	R<WL1�MD���^����U.wS�g����(泗��c2X6(����u_lhғY�@��9�?O!(泑�[Ou�LD.$�2R6b���)泋H��Z��X�ITL1�=D#���}��|��مs���\��b>�1!�����ȅ�X4��|�y)p�/!����i�m�CP�-�s��ȅ�Z����f��yM263��s"8�,���R�l'lK�k�"�!�=&i#��mW%���;0!��������/i�c?K9Kr��v�.�p�'!�N���m��W+�.>' ��3�w噙ȅw   @4YA2/E�-VVVL���	������y �e�|>�K��(}�Z�1:4HFe��ԓ�W̭���m�;;?*r�?JF27��x��l�|~�Y�p��G�RYv:�]��|�d
uNEg!�e�ذx���@��9�eu��B�_� z4$F:�2֢�g��3Ig�l�L]��漗�Z8f:��	���Hws��|��|c�"��y���9Sp������n�{��u]�����Iu�j�d&o&j���q�/֎�rl��h��Z��(泋h��Z����5�ʙJAt�̚p�h���>�Bj��D�P�/�K疃�!�,�,��3��B�I�=E�vʶ�����"�ϯ?�J���d	�(8�����5�1?;�O���k5}UZ[������r�E�u\�ԭTA�D3��B#��{�#Bj������e4E3��i���sr2�TNd���2晓?��     �KNN�	����y`��hX����������Y3���c������uj���WUUIZkB�-�bԸgN�����ku?AJG�צ��?'8S�w����|�D�vNmih����邪+�W��%f!U�]m��/�/�c�EK��9��zl�b>�b��,���i�n[�����P1M��h�f7罴��F����(Zݜ�c�A��Bw� :�N��D�D������R�M�!ݡ�|��E��7t��0�}�m�x�����=Z���L�u�Y�|F��͍�h�C�e�r@|�>���D�Tє���^��b��C�E����d����Q���R�;�-w���Ş��`_�$��E+�t�ֆV��sIrWs�g����\~��4�h��Zt~�a��گI�f� �L��[���R�p�O��;OuF��a�_���i�Ev!u�oK~��c�'���d&�~��oS~;��_�n
    �`4����Ȍ�hH���	���c��h��G�����3vKJJ�ӧO�k^�9v� :b2(F=?�%��x^~��	�V��[��_��:�B���|�XlivYHeѰ:�E��RY&K&M��|��n�{i�����t���~�����X�+����jAdE���^�EOԻ9��t���[2O1_D����w�pJ�b��v7��P�Z�g�9� �Ԣ�|��jjDV��9��/f~I1_��)��2||���E�X�TD?��B1_�������!����.s�*�-D�4D�.ܙni�o��ݗ%��4����7�o��2`�����R�.DP�H�){��ZL#��N��um��C�6]��	$��Y{��Zh�=z��:�!��D��BH�7ZQ�  ��IDATdbc^~����u?�=V yO�gdt}V     ����(yyyf���������������IOO����ʫ_�j����>�uFA�Ũ�����*��y,4b�^@�þ�ȤgApx�l���N1_�إ��~���r�e��d�ORݪ�%+.���X(�<�ts��t�k�.�:)��;��pC�R�j�l�NN�����9�E1_�٩��^]'�L�@��"C��w>�?#vC1_�٭Pg7��"+��۵��u��)�1���)��ts�k'����dlf�ώ!������A��9��BH-�E�	�	���Bj��5�ފ�
Ad��"���Z�\k&�L�Y%�_F����Ե�*$Ƣ� �/#G�wk�BjY�Y0k.�\�6�Yc�|޼��j�����G�yU2=���c��F8�7Y4)�'z�nv�_��m�D�CH���|�|b�����' b��ǿ!ߚ��}    ����f����]�b������b��?�N����g�5����DVL��~��ݟ�?���R��' b�Gǿ.��w	�N1_�-�ͮ�v��[��.v�םRY(��us�K�W:�E�v�47�{!�Hو�R|rz�@�p������X(�;vs���%��b�b�p�_��9�>ݜ���/r�c��/2��kBH3�{Cr!wA�ϴKS_A�af�n�{��t^�,O� |4�Ou�Bj��/2�r�|XF���]Q�9v!��W����jA�]U]2]4-v���v��t�UI�'	�g%sEn��;��e�P�/���/��2��]���r���p"`.N�k���ZZ�JWp~���2�LHL�=CH-4�;?6.��]�`�4]��;���4A��9��I>4�59�u\���
��t{iP�v�Y    �Szz�����n�z�;�1V��5� ��'@�{����@^��W
"'��bԲw]~���������&���.wZ��##\@S��pS�|L�,�',��P�^NXHe�b��ڶ�a1,�9;wsދ�|᧡Z��u@����q�OԎ�R�&=U=2Ul�n�{Q�~v��W�w���UBO�g7�L1_�=M�(��ŜE�S{G��b��rB�e>{�t~��/|���y?��&T,ۓ-=�W�{��3�N��T�P� <4�t�dT�b��sBH�e�l�́NN���	!=�a�[ٝ�-�-r��$�Y�N!��~[�(�/����H�!u�7$Ʋ����$�p�ԁ�ݓ����/赆�U�ȅ�BH-4�	���c2X怵�9O�fᄑ��v�����Q�5��$���;��    �L���RXXh�K�x<����3VWWM��>������M��3�<#���/��Ћ��4�+��=��w��87�2�6#������2����bK��B�I�,�.�jij���q�������	ݜ�Cg���H�0�q���j�x����b�漗�Yݝ)�-'ts�K��	������,���X6�(�'��Z(�B�pS���c�b�ξ ��<��2����y?��R�zN
!�hX�v�6�|a��R�|�c���;#��2R6"���=-3�<�_�:h~�E��nȵ�k��e~JK9Kr���8I��n�'��l�L:N
!��F8�7M eb�Aop��z�$z/�F8��R�p�C�=i�m��4�	��s��!1!�Q��o����d%s=���M�����k    �\.�ee���\[[���%Y^^��md��>֡A3@,������O���FAd��*�o̵K�H�������-l���c�^�-8�|��n�{i1_CB��S�ڽJ靴��B1_�9���~t���K���+8�ʹM�.��b>]�0� d����9�a1󅖓�9�E1_h����9gؿ��^�V ���iǅ�Z(�-�_�6�:*�ԢAh��r�����n����/�6S7���ّ�K��B,�W�S�#S�	��P�z:��Bz'/7�D�h-AR!`Bbj��b�sBb,z_����r��y	*���9i?�RKoe�ٟ˧�G��R��i��pBé!�m���Bw���Bj�N�T�x�8�pBˉ!�N1�>+���1yW�%%�{j��y>�����s�D    �'33ӌ����oz�^YYY12���j�>�Bet1�}}}2;;+��ł�����������& ���ے_����l��a�i�o�/E�h�����Y�)g�H�,�|G��T��B�iݜ�s��-��B`ݵ.7�n8z!�L��)T�����:Nu�\��Bb,����Y�u]�����sb7�(���YwS�2�ĩ(��{���焳�9�E1_h��g��Z�����U�t^�D��O��̉ݜ���|�C�R������R=�;���)�;s[.�\N�96<*=6t�t�Lތ8�|���R�d���|R7T���L��[�:�SiPq˹s�2m���Q���JGM�8Y_E�l'nK�T����񵥩ő!�ᄎ�-u��dm�ۤ~�^J�Kh�sN!��'t���T���6�'4t.���>m�ayO�g�W���c��i���}Nn-9{�0     r���%??ߌ����k����	�q��f�c�n��|��ݻw嵯}� ����_~I��
�r]�'���{=���Ug߀v-6�[�x	�yN��WoU�YT1]!8���M�z�E�NG1�9���~Lg��sR�Lg�GaBbnH,���Z�w���|���ݜ|k�`4}���P��(4,���3�9�E1�јn��7e=�yݜ�����u\�ԭT���J���%mK�d��𶓷M���CH-��χ�v���Q9���^';�>�^J�(�{�Bjqg��N�:�?"=o�8����L1_�%�]���Q,e/��5�`�`���������UwKV\�������|�\k�&����Bo���Z�ˆ͵Փ�'�gBH��Bj����J���d�96�Ε2�|�Bj��_>�';e&��!��M,��:�s�mR�Q,o�|� p��ƞ�����59    �=h�LAA�/��������������|aaA66��8�344$�����|��u}B�s��R�yL 8��=}g�[[I[�|��b�C���T���~� ��|�c&6ވ��T��M�tsޫ��M��d�b��X�X��ck!�;�-��ަ��b���~t�-�|�����:%�P��h�I~��pӜw�
�K\?w�b�Gݜ�>>l���Vʖ���BH�E��ֵ�do�ݮ8�X��WWu�	J+�-\,��X��;�|���w��H�.:g����b)��2S0cB���#���ބ�.�B����p�G��p	NC}�9D,9>"�d���Y�al�l� �X�_����R����ۜ7T���0bq~i�υ�t]a~y&��d����F��F8�&�BH��#��Jij����� p����LP     ��r��(+������,--�����l=֡A3@�LMM��瓤���;��"��\y��m�ot>%��R��# ���ǿ%�0�,�,S��x�,�H�J<��$�������H;�颠ʩJ���y���5�RY��O[>���$�b�=��S���Y�Y�X�8ڙ�x�X�򖳖�N��EZ�����|�yI���/�L7�3�d͵&�H��.�^��5���o���y/��´��:��@tn�ߌ�n�{Y�|W:���M���*�Bj�b�@R@NL��<����X
!���NV5�����s}�E�p9x������V3W͜"i1��i)�|/O�m��̼<Y�|y�y���Ŝ��r��L�4Fz&���M�H���`:�l�o�+=W�9�����!������S�$���r�R��y���5V#����MX�A��藩��
!��W��cC�a��!17�nJ,�����V��}��� �~�]sc+�Ԣ�pt>AX���~�^[!�N����9)Jϑ��5�n/��|�y)    ��222�x� ��++++���(���j�>֯i�s^��Ĭ��IN��k�����o.����M�����\x��d	 {���-����
�C���`P�ǆ� 6�7������Ov�~ +�+���@�9��H8���9�֥o	`�b�_�ђQ3 ��ι��z+{� 4,���_�>-��|��|��7А���V�D��i��t] 5P9`�������<�)��y>�����w��,M9�v׽2.���1��    �����%??ߌ��Ë5�cyy�Ƹ��>��_X���	�����Q������)�I� ����yo�gM�                Vm��MX̻ϽEj���=�M˯u��x|�    @�JJJ�	�y)�G�X]]���������!�1� 6�A1jxmڄ��Ϧ����t`/��w�{�>CH               �oC�{Ǉ�νU�2���Lx��u|HV�     ޹\.3���=�z�;�1���d��t��@�:r�0�>(F�Nɯw~D���fIOJ ���Ҁ�n�ߋ/�                ^,o�˯�P~��OK��H ��̦[����,n�
     xy��ɒ��oFMM��wɬ�����	��P������Zs`7�b��syT~��c�o���Z�h���o_��~�                �F�(���!y���JIZ� ����e����1a1      4v���������N�����:���dkkK�xB"�.����������� ,����!��Ώʆ�7e               į�M����'��M?%%i� :4�mOʽ�E     ����$���f�����k<�	�Y]]���e$c��,,,��Ɔ ��4�=n,��o���V�ŕ�& "�e�O~�����                �Mz�����Hyz� �,�yG��2EH     ��r��x)^�WVVVv�c4HF�[_��@@ � (fm�a�ն'�w��,��.�z�]]����W                �7��_������ ՙ� 2F�g����e     Δ��,���f����|��_�����KFF��5>�O�~�lnn��ښ	�� ��m��A1/�wuB�k����7KnJ� �gg���~Z|�$              ���V���F~������
^�kS���?$���     b�ì�������B���0�2��鲽�-�G���eiiɄ�蘛����-"����X�2���nz�������T������@�               ��V��o���jz�4fW	���X�_�xJ�|     ���5cIMM���"3TBB�$%%Ibb�x����h���������"@��2�<s�_�5u��r<�@ ��'ƿ)O�<MH               p \�?�?,���'�r�iZ-�}�;ݟ���    ��c�И��,3��ʤ��фɨ��M����۽&��5�Ff��"(� &=���_��?)M9'��g�>࣪����{$��&M�M������Dľ�UWwuWײ�������
� "�TtA��&@$��>ɼ��?�H�B&	�7��r�̝�D'w�������ޅ�"a�                �/�0_�m���Z����@�����zy��r�
     PLL����W�V�J\����Wa!�G�=�bܔ���#����vWiH��p�����>GkRv
               @ř7����I��/����Ԙ/l}p`�f�-      P�����"���s��$��C���3��-3�;+A                N��������ڏ���� T������kI�F      ���
2�hS�N�K�=mG���G ܳ?��:SG���               P9�'mQb^���t�����{2�9zr�ڜ+  �������
]&�-   �P�)����r�g��\�P�@(�j��c�\��	               @�ڞq@l|KOt�^͂��lqىzb���q  ��5Mk����+t���p   �bN�O)�t�7�X�k�*�� ���r��C+���o�:�               ��8���{��G��R�:@�V%o׿v�SVa�      ���P�i2�����G�������d;����y�!y�                �y9�y���9�"��nmu�|���E�"������)*      P����.��߮O�-��js�|�|���d�߶�RBn�                T�����d%��sƩ����]zA����֥�      PS��D�(6;Q�0N��������Q/�Z���               ��Mi�u��7����!����ծ�x=�m���
     ��	WJJ� w��d[�cu��7�P�1��F��$�0_�ٻH���                �K�O����-�/Ѩ�}���%�l�r�4?a��ٿXEN     TG����b�6B1g�#?C�n��+�Ӕ�����Ì�o��c��ڟ}T                ��|�S���R������c�&��K-��;?՚��     �΂������b���?j]����5j�@@md^�^�7�~-��P                ���S��u���vW�_�s�VkSv����R�)     ��.  @��Ŝa�YGu���hJ�5�a_yyy	�-̇��o秊I�%                �_ZA�����.j�Mw��\�>�j�|�S��[�	��NQ     �چPL04��g�~N٣߷�Bu�C�t˓��ݟ)Ù#                5˷G�kWf�n�ڄ4P���J�s;�*.;Q      @mE(�
�v�Э?���[^�z���K@M�R����|iC1                j�ج��w�ը�nj1L�>�j����9�B�,��U(      �6#S�2��zi�gZ��Q����AQj�˥�{ݾ�w�2�9               P���4?�G�cT��{���j��鱚�k��$	      8��Mi�u׺�uC�!�d�|��TW	����3�O�+                ���f��-�5�~W���R�����N|����Ykw�
      �-�xP~Q��ٿX˓����T������P\�Yq�+��               ���7�=�^�R��wm.���T7˒6������)      �lC(�ؕ��׽�a�ꖖ�(�/D���Kݣ7�-Rl�Q               8{$�g�m��-���h5B-C�9I��w�~J�%      �lE(��p�������t��j�_~�<=�z�r������&e�   J��u
���|k��$�           @M�>u�~��u]Ҡ�&��:�����qK�y�j��      ��(�T3��\����>��njy�FuP2�9�sp���ANW�   ��>�=��M�           ��L�c��-KڢqM/И&����G��f�k���:�����      �PL�u(7Y�l�H��ӭ�.U��hg���|����D�N><               p2�cJ�S��7趖��gݶΔ5);��ޯt 'I       ��PL5�S�.Ť��Q�tS���$(R@ep�Y��U��.V|�C                P�ج�����\7��P��PY�d�i���1m�       ��PL`�˓�ب�	�Ln1\���	8Ł���� uu                �`kz����=uo��ZӹuZ
8U��4#�Z��W       JG(�)����]C꟫�U�����r��&e�f�~�=Y�                �kKz���G����}h�ڞqP�|�U�      P>B15��U�o��ײ��uq���|5�'�$��"-Kڬ���^1                ΀u�{�~�^��w��i2@��[(�ƴ}���J���)       �#S�廜�"a��L�I}�����
;`��뛣?듃?�h^�                �Lr�\Z��ݎ�!�tU��5$�\�xyp�Y�ةY�i{�      �8B1����t�c��B�����0�,�R�i�A��W)ә#  ����v���M�-L^���            ��;+A����ޏ���j�_���@��cv��$q�>9�R�r�      ����eve���?8�DW4�a�]�$�~�2苄5�>q���B  xRN�:�=�\E           @����=53v�F6�{�a`]����qhё-:�Lg�       �>B1���@�|��־oԯ�9ٰ���i-///��0�/Kڬ/�hO�a               @u����G�i�����Z�女Q����'�EN�r����1Z��W.�K       *��Z�|Ⱥ<i�M#uI���AE��5׮�x[U����                jױ�u�{�x}�B��э��eH��:����G���#?+� K       �B1g�C��zg�b͈���E�����w�v�k��9IZ��Y�&�W|�C                P�e:s��p�Y��a�ua��� �������/%?S+����n�8        g�����U�I[�0���50��.�� �1��ѼT��خe�[�%=V                P۸\.mN���=_�cX3���Q�*�/D�>2�9Z�ة�I����~?      @�!s��/*�*�;^���GuР�.��F�^>B�;����ɛ�}�f�ʌ                �-�\Ev'�f���k�m��ƽ_d��
U��a~Hަe���>m�
�=G       <�P��*�շG����N���=���GvT��(��0�o�<���;�.u�vg%�">                �͜�B�I�i��no�	i���α�mH#yyy	gF\v�V9�k]�^mJ�o�       �G(%�+*��3�ٿX��{D��z��m���K�t�M������Mݭlg�                 %+riWf�3㖨�_�Ϋ�R��uP�z��$��tg�6��۸�v�Pr~�       T?�>����%���c#��O�Ú�Kxu
k�����(��u�'6;Q[�b�%#N[��l(                pj�
��<i��^�j�@��6�����؈Jw4/U���5�l���YG��      �zN�S��Š��
�)m��ױ����T��:�5WǰfjXW^^^:��iwf�0̶c���\  �j����I�&j�\M�4Uh@�|���c�]�S����tJ;���x�Oٯ¢B�f0���Md5�h� � ��ٹ��ed�@��IڣC��r��
           @mW�*��;$������������)�������Gg#��P����(�֌8�I�K      ����l�"��f�����ڱ0�'{�� �Ip�څ6V�h�����MT�?T��#?C�2��=v��r��HI  �
������jH�!�Ӭ��5�&�/���Ӷ��s F��.Ӓ�Kt0�����v�V]w=���;󕖛fGjN�����7y�bSbu&<4�!E�D�8��w�#q��B���{�Xl=PZPx�{{{2�ӊ}+�����O�'y�            pv8����&��ў���V���۷�mݏ6��U;I5۸o�n�s�:jG���R     TW�E(g�)���kQ���C���u� 0�À_�����1��H^����pn��Ä<���ˋ
  ��g6��v��<�N��0BA~A�|]��ָ����E.�K?�Y�n�T3bf�@�J�ݣ:����ʖ��nc(���Fo�X�3W�����v��lS�Yߙ����������R�f�O�:���e/��#��Uq����W5{�l
            g�BW��mܗk����|��2��ݦݎ s�ǎG���K�+"St�~$�g�Hn��m�S�?6b��(ә+      �,����E(U*)?ݎ����xL���+�7�~�^��a��_N�������K7���/�z~�/a�g����������,9�3����r�  @�1���z��'չa�3r�&BӳiO;�z���_����Y��*<0\�w�܎����n��g�{F�6��1��Ğ��%O�E��z��[��㉋�У��Q            ���6�����[�^>vǨ�#��p������m�Ͷ����c���������ۭu��������3
����:v��m�������Yv'��yi�r      �=�����P��wq���������z���"���"�\.eRD  �:6��Ƽ�!m�T�:}�}tY���X�o���a����3s��wo�:/-�Q�y�	L�qo�v�����j�9����O�PBz�            ��2A�C��vT�����}�� o_��R������e��       N	��
��Lg�=^|  ��cr��z������pA����z��7t׼�T��z�������k��������lX�a�h�G����u��<Z������c�*v�            ��R�*��6�      ��A(   @�e��3�����{*t���tmHؠ����K�SF^��yv.�/PQ!QjZ��ZG�V��]����zyyix��I����n�N�_���UG7��Qo�{��m�q4�V�[��;��S��5�yl^��:��Z^����r��qxc-�s�ƿ?^�,                    ��    Ւ������&�����1b4w�\}��sm?����~>~�ٴ�.l{��>�juo�]����/�m/O��"�"t^��4�� �b(�6:W3����߹\.�K��=o�;�ޱ�wYLfF����m��)�~��O�f}4���
�,u� � ͹q���~�[�                    �@(   @��ҕ/��1a�g�}F��V��z

�*v�����P���p�&���ЀPU���jڪi����\��b=<�a�)�Ȏ#uc�5=f�����]dc@�EbL ��E��P�!��ۄd�k�-���y�?5�ۄR���񷱘��֚�5j3��֢nPrd;t0�}/,�yo1���<߆�2�2���:��4O�7�WZn�P�� ����j`��j�F�"��9���M���u�h��/W7���7T�_�]&>=^�E�                 �g�   P��?�~�u�]e.c�!S�L��;���uo?�]wz���1=2��s�=6�P����f����/(�7����6�o��n����i�#[k�����.�KM�⦏n�'?9�uť��ڙ���m_j����T�r�y�d�'�=��gP��	���/�[W�w��5�vyOؔ�I�w.�g[>ӏ�?�e��z{��'E�L8�YD3��<Z��\���}���Em9�E�3�~˼���6���z7�}Ҽy���/}ZZ�'���k
�Օ]�ԥ.�sM�4=�2�}���yk�[�j�W              ��쐼*v�z��   �   P�to�]���e.�|�r]=�j�<z�nGJN���a���U�>�u��0Bՙ���y<�L�c�%1_�{�X��$o/o͸v�"�#K]&13Q#���1��ޙkg*��ϧ|n�%1�Ѵk�i�;���zM�!�z�%�q���_=����O�I��v+:4��'�L��־��>����7W�)�c?��H�Z�Sӈ�v����g>\��?���S�(���������n�`�`���ϱO���_-߻\��֔>SU����ꕫ^ѝ��T��V���Z��1c鞥�q֍:�z@              �b���"5  ��|||�t:���,�á���FQߵ���    �6L��D�|�J]f��%��(e�gU�m�M��ȷFjr��z�ʗT���8W�^�o=0��R��u��C1w���P�|vA�}�+3S�82�𖅥��Fu�	�&h���jt�n�:��`/&���v�p�a���\���Qm+���Sj=Ȏ�4k�+�\i��#[u�����o��	��#>��<h<�V?��}���˜��;Wh�!m�h�����~s���g�Y�ھ�                �V���6cFaa���󕓓���,����0̑#G�q��%�2�   Pm���vuiإ��]I�4f��*���ڻ?�k�����ϩ:{�����~�*, ��y����QaQ�<�nP]=}��e.s����c}��@�>��^���R�y~��y�r���+�yv䳺���
�PMЩA'-�}�>�����ߕ������լN3�)(,�χ~��Û=�>�)���߲��G4��s
r��=,�y���15��DՉ	M�bj��v둅�ؐ                 5I@@�BBB���`(;;[������PZZ������A�"   �Z՟����yg�S�̸F�9��G����Ru����y��iR�I%Λ�L��m����"�"J���~�f��y�o��+_��.����K�71.zqy�1����ײ�-�9��&2�3Jc��^]���.������Чy��ϼ'y{y�6i�V������I=��                �:���1���@��������UVV��<xP111�`P��   P-L�=Y��:o��7��

T�}��RC1���'B1&t���:����?{�Jn��`����j����W�2}؆*L��j��W�^jQ�������3�2l8eJ�)56㎨�(���jr�ɚ��D-ۻL��������0��.�[�4����U'����srV��d���۵��z��                �ʖ��c�/fdff*##CyyyJHH���q��    �Z���m�Ι0�߿����M	�ʜoR��<a\�q
/u��/و@U1a��b�ӭ}o-q�qxc��0B�o�\@Uh�\S�N�=nP����/����kҬI��~�j� � ͙8G�w�\g���u���=���oi��5"�                �~�1#55��`�HJJR~>;6E�A(   ���m�W]v)u�|iܑ�ܓ��T�|��<��7�:�_��WV�����e��-}n���W��7���Pθ��=w�s���������u�\.{X�k�$��Z{p������������Y�f�������uq��=��]I��cڢn�
]μf*�z��@�@]r�%vH=��?�_�l�D                ��[aa���ӕ��i�C0��OKKSQQ����    7�Ө2����=�}&�P??U���hh9���/�~���xU�mG�i����zP��&X����g�9����[�T��6U�^���|���Y��m�q^�����]�e����+q����0��u�|���%s�f\;C���Z�e�j*�xͺa�G"1?��A�/}^���>az�˛X��{�ײ��l���Q�+�?DU�YD3ͽq�^^�~���*r�=                �VN�S6�b�/&cFq�Da�w��P   �j�N��:���VmL�(��^p�2�==1Q��o�X�2gÜRC1&c�����<���ܹD��yd���{9�6�aDE��WhR�I6Sҿٛ�ܬ�������_=�W�zE�v���u,ݳT���:�ѹ�}{Md壉�����̣����������_���c���j�=��̵�s̹ctU��*m��[�s��w_�2��v�w�~g�3�-m��[Iv&�Ԍ�34k�,�M�k��~�L^`���=�c#5��                j���~111��1Üg�� �#   ����U�F]K��v׷B�4
+;:a�UmX�a���_�Sn[(��m��텄bpZ�F�U�f}�>����y�Y�{��J��ħ�ku�juj�Im"�ظJY���){��⧕����1��hQ��n�}�u��˯M�b��o��=�{4���m��}ſ�0��I�߳iO5y�������|�N����8�o=<�aM�h�b����cnn������L��q����͸vF��&��ܒ��̷��P���������s9����������N��H$�P�!m?�]u��G��,w�����+�?؞����mG�i������                �sL�8�R�)>m�0���Py�    �nM���˫�����
3�Հ2��PU�ޤ{�s6�@���s�����jZ�i��=�V^� go/oM�5I~@]v���6o����;}����Թag���|�k�Ͼ7����˘X����Z�e���bSb��7O��_������N`;g���a�1f����;��?�%�\r�u�(���O|�B͛4��8���%�f�a����?���A/�xI�bn���h`���u=G3��~h��L ��yw���o�ߟ�Z:i�3}��Zw��Z���C��H����\��v'�>�:�E4����I�I�Q�c��?�Yi�i6~4󺙪l&4T��d�'z�gl8                P�
m�%--M���6�b��6�f����Q-�R5F(   �G�1�ǯ*fD�e�o>�YU���_�t*u�����i?���PL���TDdp�>��������	h<��Q
1�Օ�ڹ���5��H��8RC�����=��ן�)�����?e/����m�&!#A����\rv�.{�2�y��GN���ﳱU���kj/���k��u���m{{��)�os��|Q}��є9S���SU2���RC8�Z�w��.��y7�;i��t��~�V�_iO{�1��_�f�7�n�u�9��5qkԢn��w���O
����Σ~����rۗZ�m�VŭRaщ�_��R}t�G��u}�k������ݯ�x]                 �9�N�1���L���� ���8�)**����`�^^^պ~D(   �G��l[�\V~�bSb��o�_�Z*u~o�^�J�굲���l=�U����]���B�l�����[A~AZ|��r#X�S�c_��|y{y��dh@h�����?i���Z�}�	��L�i���S����6^�u���E�b�?��ɚ3݆_�EΓ�1�?/��6&l��	���M	�l��X|z���>T����������;�^%f%�˞;!6S&�0���L���tUs_>��q��Ky>��&̜Pb�k�c���1�3���~zOw��=��m0��b�-�O���^o��F��3���;4w�\}��m;���e�7֬�g���/�WZN���O��z
���2���Ƽf�ӴU�                �Enn���������Ogee	�>>>
	9��T�b    ��"��:g"1�K�pO�o��^1��e�����Zӈ�e��s쓧�J�U漹�b���^��J�Ę���ݬU��t4��I�u��MT�k�O}��U���6��-Y1�߆b~-)+I��|�w-ݳ��e>Z���d�G?�mso;)H����U�]uR,�8���留�i����n����]<��3��y���8׆ON�y�n���	�?��]R$��c_=f�2�����[�\��HHOp��6�����ֲ�1��8�<��2���q��0A.*���u�Ѥ��y�?էy���|�F�Jz�                �6���QJJ�233���n�/�v U�Q�F6SK�T��   �QM�4)u�|��1��wƿS��g��PU+�96RsR�i���~�5��T�7(�	^�s�=�r]���������֒�N)9)�9c�++_��5o��;]n�&������)&(���66�R��X̷w|�-��~�z��7lx�ّϞ�m0�/�|�K�]��l�	��Xs&�9�H�	��8�F�1�R�ϙ�ʅo\Xj��D������q��Ӂ���̳��,��ۍ	ݺ���m"ۨw�ާ};L0��A����	             Ps���m�  ��\.��������94!�_a�N���E�B�    ��L�4���(_ۨ��q��oѿ������\��V7�n��i�i򴣙G˜�\�} 1��,{NTv~��w��p�<���j�A~A�)ȑ'��)fb1WO�Z1�����ݟ�=a�������CC:��0��@�;�]M�9��ǰ":5褹��*�7മg����q�/�?~ފ}+�:n�z6�q�;!�SOFb�%��He�gU���M�������*嶌�4�P             ��ٙ����U��G�z{����Bw p�),,Tvv�����& �p8�y�xAA����[�nB�    ��}K��-ȭ�u��J˺-+�b�(5'U�b�	Z�=o��s���ۧ��
t����	e=�FuŔ����`����J�����n�~�`�.��H��g֕�]�<g��:i��_�Q������2�q'�2��8�;�Άg*���͟<_aan-o"0�>�'����v�z{�I�A��u���%���&8�H��Σm謼�aѲ^K��d�e              ��6^��H7|x��)]urc����7�m� ��e"/&����f�9^<�i��읢�вeKEGGU�P    �
�*u.�0�R�uK�[�ǡ�����`-ۻL�ebω�j@���z��@�M������苇���fyBYϱ���N��D���/s��@���ˌ#*=/���˴��`�`5�h��T��)u�|�}�Ƿ�y���z�	s�.�p�FtQ�:��6�oТ�N����ɬ�g�]T;��7��fߤŷ/>����D]��eJ�I)�r��ɚ�i�j+�8^����<����������a��P��]X�o�P             ��жC�����q���j�W��9�XGӮ�fwg����  ��N��������p� �9n�3Ü&���l�?|�p���   �j�udk;΄�A/.Q��R�hU$xTg&�Rٙ�Sp_�3Oc����A��?��_��o�۾��V˼o/o}x���5���$�9����%O�@�;Lf����vd����������^���{u�2Q$��(���}L��"1             p���h-��P/�|Y��vgv�лYo;a��v �ʔ��ic/iiiv��ŧ�a^^��$�����&M�U�P    ��)�QDPD�s>©s9���G����=z;rr˜7{H�I�'��9o^�@yv'�.s>�/X�'L��W��p_rv����xϏ�
�ҡ�Cڑ���]��Zu�*��jW�u��5o�{K�q�)��6�?��[˚�͕�]i#1��{��=o��4k�~��Q���/}Z]v)u�H���             p2���{/�W�w�u\g�ǫ�u?w�s���  �f�����8)����N'��eiݺ��.T-B1    <*�YzD��xJ�&n��w��\��R�sl�P������9O(�X�e���k�O��_�Z�/�bL����ҷ����g?ߑ�Ш�G�XLi�bC�ѭ}oմU�*�~�Gi����qk���ަ��p���sl(�ϋ�l���L������̊}+             (۠փ�����i�M�rۗg|}f'qfg{#;�  U���P�����̴�)))6 �p8�qs�Y���ر�ƌ#ooo�j�   �Q)9)ju�$�!т�

��������CS6��s\����Z�����`��ɺC�ԽI�2�{|��6tr ��P1&2��qZ���(ώ�v�&_L�B�^e�h�D�p�BL;X�u?2�ui�ŭe_��͈�q�y��̹Eo�y[�8�yu̫�>�Dx             �=&���͟��/��R~a�Y��6�����qxc P���󕖖f�/���)>4������6����СCu�y����K�z�b    xԡ�C�ѤG�s�V��ĭѴU��^~\�q��Pu���.G�C�oV���t�'��]eϫn��c�\W�V�k��� {e�+z{\�!�ЀP�0�]3���>��Y��/ھH�Z�/�q�˼��S�2�]��n��C�ztأn-�:n����O'�_�*"sn�w�z6�Y�2�)�o�/             �{�{��^�i�GfNPlJl�]��A�c=��\�{�,��\ �[999ǣ/��3�����UݺuU�^��͛7W��x�    u �@�s-교����r}e��i���zP��b^Z�^\�b�˥d�(57�F���Yi]��<�}t�2�˻@1�p��s��F�ic�F���e�_4��@����2�����=~��en]�#�����˥��?��'�7�n(P���$9��             ��>�>��qY_��ע��=�N7ts�찫qxc}p��fH��nJؤ�3� p�1����;233���q����Pn.!1�L

���q<c�����    ��I�K��V�z��'y�j;�ٛ�W����R�3�~ѿ$�v��unعԹ��G��v(�����u���Z�|P�А�4q�D��H��^�MnRh@h�˚�����o�m�׆e�q��{�߱_�\�zMR��F�.׵qWM�3Eo�~S             �_�Z7K����y�L5kP�ru���ӛ>մU���pf��S1��0���a�]����뎹w(� [ ����!3RSSmƌ��$�����gb0��Ѫ_����GaL&00P�y�    ��\�|�&�ϊPLmVPX��G���$&��i���.un}�z�:�ѹn/?��x�yџ�'Tj��W��+���\��}l ��=��kԿ�*`��K�\;S�\�^�zp��n/�̈g4g���	             ��ow}�^S{��>��V�\��~��W�^���2w
�[f�{��/zl�cvۯ�d�e����ۈ �f*,,Tzz�233�aq��p��iii***�3���Waaa��/����8��G��3
   ���Z/��U�������
5ۺC�J�ti�E���ɑ�'��j���K���`�1#��h�����ӄ��ܒ����uM�k4��2��ۥӂ-���0��?�&Jb�h��gbb�ۻ�|th�&����V�$             ��L;����c=Vn̥G�����ݎ�4�h�Y7�*w�=��h�� @�s:���Ȱ�1s��<s���T������3L�Da�����\��b    x��r����gӞ%�_|��B��ݮ�ts��K�3d�q�f��)O����eΛ���w��jY�e�/wE�+ŜE�"�n����k���S�r�v��#��/K�h�Cn���o��@G��yt�/3��8B1             P�¢B=���~�����(�Q�ˆ����?�;]3;S�.�.q9�-�;�߱;�,ϴU�t��{��� ��rrr���i�/�!�1�8�����(<<܆_L ��_��0QQQ���P�P    �3_�/-�.���[{p�Ps}��k���҂㺎�X(�J�������(O�&�N�r�Z�S��:�q�Rn�����7VlJ��v�7���o��w����(1ӭq7m;���l;�M��|E��B���3�*�Bf���ޤ�����             (ْ�K��n�q�]r�%e.;��D�=����k�������s�?�{�c��*�ٹ�ߪ�7|, @�0!���Kq��trr���vU���Waaa�_�����m�DaL�N�:����B1    <�-���Ꮧ:?��dB15\rv�V�[��m�8o�4�<���R��vum�U�[�/u~��E� n	�,w��1������h5kh��q8��TV(���@)9)����6���Ou0��V�}���w��AuK]�¶�(����'�o2������~�
��1�z^�g�v'�����̣vc�^������D���ƞ7*4 ����D$             �a����=<�a=3�Rwitj�Ik�[����gw�ֲ^K;a��6�[�z�ĭф��ϱO ��QXX�����/���r8����4���@�

������@e    ��L�|A�|Q�$��L�S����@���O������}�Ӄ�?X���Ae� �Y� w�8Ky�{��_<|�oKzn�f���F�l��U�V�p݇��i�2�2u6I�Jҿ��[O]�T���s�=�2g����C���Ly��Y��w|�����ˠփl��D��������J_OV~���>��Gu��ο���9r             ����K���q����؝ߕ��Xl�5�4��(i3��`�,E�"=��9��7g�S  �9������L������L���H ��������m��`L�8%g�    ��~��^�z�s�~��������N���n���WLUDPD��w�K/�xI�)�Ur{�kt���q}��q�q�f�7ܱ|��r�11��~xM��U�t�'w�C�zv�z��W���Om��N�w�/-�F�J{�1��z�����v�V�>�8���u6i�Z�{O�Ğ����G>�[T�m0��?.�G�ˬطB              ���
��������xg�5�C�b@Bpw���-P �-Z(�B��o[�@q� ���S,��	�A������/���$�����z�Րyff�;�3�y淜��yj�m+�}E����h��-6��""���A0�"!0���ɿ���D�����C��#�0Q?K�D	�A1DDDDDd��ÐC4S軖銀#8zd�$�a���*�GG;G�o4��42�k�Ib��M&���V���;~ǻ��@d�������c(���fY��-@�ɕ�g���Σ���(��F��]w����`���j��2��ɫ'*�jh���m�W߂��2_��]�v��W�Hv\�k'��zy��p��5q���<L%D/�������m���
Q�<x� ug�E��=1��(����j>:�ja+�zzDD��˗/U��������S�"��d<%��0OOO5D��H ���#���b������,��|�������Su��`����Q|\qu�,��=cѳBO�pJ�s|��ѹTg�84ä���*ߣB�
����a֡Y �		Z�z��6��:����G|�wm�M,����0��X����cꁩ������2 I�j�i[��
�)��
�+�<G�k��5-:�����3���!��`ܞq���H��� |W�;�m�=���i""""""""""""""""""����Wuy �zv;kʬO+4�����6��5Q�s��%�;waaa*�����>����I���?������D��A1DDDDDd6$��K�.(�����Sd��kQkF-U�N�G>��c���6O��Uo� A���Eo�>���ͻ7 ���V �z�g,��]���q��m���Na�ٵ�\�3~���K�WÑGT`L�@�x��DƖ�\�VE[i����<�=������?�������$I�UsTE�2]Up�����[L�7	öKР���*���5�3d�D��Şt>Wir%��w
n�nѶ���|���n%&
�j�*�����⟳��'0��8"kŠ"""""2R��6�-Bz� �]R�mJg.��]����&{�<�NC�"-Uѿ.�ٯj�
f7��+{����yj#�?�6ک�+O�TQLI�햴S�0G;G�m���B8F��� ��)��`�����O�^�;�e(��f`t�ј~p���擛��L�#�����0���<4Ӫz;���M�6�[�/r{����������8}�4R�\5���J8�;�m���*,8� DDDDDDDDDDDDDDDDDD7yR����K
�)�R��w�v��5Q�q�����ꤓȜ��������0���eppp QbĠ"""""2+R��wM_Lj2I����{߬�K�/1��Ib�B�����_�	l�ý���Sg�����f����e&I�Da�m0V��*�C]WtQl��sF����Go;Y'���һ�W���
	��@$�i\�q�������W�^z!�X ���S�O����_@.�\�m�)�
�+�w>��sx�A�d�Эl7�(���S��凗�om?������cf���rQ�s�6�[Q�H�c��LFr��O#�E�,�岔C���94""k���c�����\\\T�K�ԩ����!���666 �O1(�����������U!��h������UQ���~Ŗ[T�x\I��_?�2 �Se�Fhx(�/h�-]���F�����#f}5�7T�\�ղ�G�?���yj�m�2�%�i����(.Jf*ip[�)�5eV�-����ϑP��=��>���>�4��9�`뀶�ۢM�6���&��5;.�%����|�9�h�����ȍ#���:,Y�T�T�Q��?��/�����=c���k$$yh�?ah���gCڗ�X7��Ŝ���7�Υ:�z�C�>G�����bY#�]Y�|9Cb�$�zG�H LTLԿ���@D1à"""""2K߭������]�
Y+`S�M�p�V�Z��g���ͣ*��Pn�n���*�篏�y�"�sj�����������l� �"������}y7޼{�w�pQ9{et,�M��h��D�@�y�j�!���.(��l���p��_oG��5���S$��g�b�?�UP׏�T�a�RV�Ad�s��\�����Ҭ9�FoP�A�8��J�T�U�_o�O��r�j����an?���&�ܴ��b��A�\5U�L������Act�9m	��"���b��軦/^�}""kr��qܸqD�?vvv�_�`>���'"��EDDDDDf���w踴#�x��ڣ��3U���w�8w�B�C����<{�L����'C�T��͌��\|]w�S��m1W��h���G��-����s;��s������=s�t��H�ܠ��f�a��� ��9�:S%3���f����Hh�4j�(	���E��`��F�+����y;��p��6��.����R=�������3��X{f-,�����~>w0� z���`��>�ĪG��������������������(f�o�)�S����Hǌ�@�@�k1����۾[�n����4��;�ADd��ƽ{��(1rrr�$�����C ���Z
"���ْ/���돣7�b��T�.o	�T{�I������髧 㐛E����2�qIm{�Ψ����J���m�c7���� �/6���z�(����`�+�`ߵ}�Q����;������fbjө��S%�+�e W��[�cىe#�Q������%���퓰E�Q1���G�0p�@��i6�\��B�4�h爰�a��������?��H'�ӚNC�"-�m{��5�X�B=�%�̪���{bT�Q��m-���!�W0z���f����]�z�=�5�����>��DQ�vtt���ٓ ��0����['A^Æs0h� �
�$_����d��h��a�,S֫��z��� 2������}A��WFޑy���+X��P|\q����|�}�cH^��X�?T�öC�� ����Gcs��q���N�a5��q��:��G໵����{0G�N�R��Ib��=_�z��mK�?""""""""""""""""""�^��E�3YQ����J���㗏?�N��w<�T�fI�Esz'{'Lo6�U@������sY���D����...`���?�xzz���Dd�CDDDDD���+�;�.|r�`��p��T��ˌ|��'�c��q�֭���hN#l�k�_U �)H�������F[��p��{����l#7C�S�?軦/,��G��e'��Юz��}2^�IV�]�c7���?a�ٵ0WGo���Gn�9���O5~B�B�T���.ܿ�n+�aǥ�Q!1�
4�W����vߵ} """"""""""""""""""��o���SU��>�!�<s+�0Z�3��K`n���������.�%3�D��8q���,Qhh(�̝��Ӈ�$FBa�~��y'Y��E���f5��\��tC�����)���/���׃x,K�/��gw@�+�tV�Y�&�MЭl7T�^Yg�AL�{��/m��}�����9�ʂ��[�����]�7�\كU�W��\{t�gׇoA_�o8���2�H�"X�a�
�賺_?ss���XO+A+����#j�@�`kc����o_�������-��X3���m^�y��SA ��!�W>���.Z&��DDZ�!��u��m����:y�b��:�-=�4Na��H���O:�=x� �w�Y.WGWLo:�7���?��18�E�#ȳ�=����z#�`��6�gn�y0� ""s���%4[[[���}���@D֍A1DDDDDd��T���=*e���D$a�D�pwr7x>�_>���'�M	m�}e7�?�o��<+xv]ޥsܑG`n~����!�˩ۧL��������Ր�5h��v�g-�E0��On`�3]}z5C(�L=0�+�G�d)5�Hqj� jN���W��Ҭ8���oCЯR�/�I�e)�C=�m����7����/&ȴ� ���e�c��p�9��l#Ƕ�+����s�D�ΞX�q=<�{�m7y�d<{�D�8��ȉU�����Q���!w�ݵ��G;G� ÓWOT��O��UЯr?����=��b��%��GJx*�b����+��K�x��)������������X��#{��Ѷ8��+���6%�8J��t4��	��ʦ�V�c�k8N=�ii'���%x��޾}��`gg�!0���j�KH��M�:d&"�Ơ"""""�h��"���65DI��RdB&�Lp�w�KR������wx��)"�D���Oo���{��Z�_ܮK���b��[Oo�  ����M���7*A
�^E�R��^f` %	��}��W}�F���QaR��s�F
L�G	���|.����x	�iV���}�Α��L
Mڣ�Gꆴ���Lk.�l�ֱ�)��/�a�5}0/d��{-��7uބ\����{���8'u���}��!amrL%""2TTI\��G�C3r^+Z�2�wZou~(C����%��߾��%���c���`�!߱X:	�Hf�̠�����^�'s}D�L�Ó ���Z�@����Z���X�O��E3E�tEP$}�N�[^�9]��"߃�v =�9��K;���~�y�DDDDDDDDDdy�o�em����Ao;y��ە�b��9�^V��W���B����m����B�-�tDD����� 2y�G�`$F�_�a������%3�"J�CDDDDDVG^��ĭ �#��ʃ�2���{�·�/Je*����l�5�װȰ!7g��+��>�ѯR?���~2>�Cr5�S�N�q0]���%R�����O�_%�8	M
��6�
Y+h��t~:/�B�,�����E����7+�Qa1�B��Ս2/)J��=9��ܽs8|�0v_ލ;��(J���0����K�;#ǡ�On�ԝS�������?ypS�3�嬆J�+��%	T5��z$�P��=��W��b�e'�a⾉8}�4,�Q��j�Am�$�o�p��5ė?���e��V>�TCS��sy�evaLr\��9.��}B}y��Q��T)�y�x�D����J"U2�}���T�Z�H����
$�Y�n��F���t�T����WCkU��KT����'ADDDDDDDDD��@�ц��3�_|��w��yy�w��M�m�o1��hա��<r߷�����1~�xY[[[���~
�����b���������L�H��#�W��ފEZ״��mjͨ�#7���~��DЩ �m1yR���MF��h�n�v[�-���b#�w�"��#�D��ma��Fg)`�n�w�<+A�x�J���]63��\U�D�'�{�:/�H1��u�P�!,:�H�����u""�x"��;z��F�<������^��������ͻ7H��|��wcU�ml��u��ѥt�B�u�q��X3镩U�V�uۯ�<y�y�� "�u\J�^�k��S����ٌ��b˅-}n\���`ݨ@2�gBb&A/5s�D��T/���.�s�=��������GWADDDDDDDDD�/�H�z��؝�IG���Ò�K��#�f;���k�_CDD����C��#�0Q?�3*DD�Ơ""""""""���Z���NTq�>����vԝYW��TQtlQ��5}*��hR*S)�3v�X�<�������c?m\��ǟ��T�8k�~q;:.���PX�t������/ڶ����	��fU�̥�0�g8���ڞk�>�9������\sȦ!�A��V�_.k9���|L��M���v��賦��k�_�?ނb�=����	�mT��$W��hF�C��Zn�!F��Bu	rPe Zk��L%�|AB��[�
M""""""""""�$��=W���C3M��.���b��;Eu�@DDd�>�I�:5<<<T ���q:n "�	����*�(�ހ�(n�n��y�Ϯ�]�w�Rɍc�M8�T洘��;;����޾躢+�^�o����+�ӦvN���5eVus�'��f����u�cʁ)_(��=�
L��s��V�^�Wo_�N
������+ꇦ��⃋ ""2�L�0��<�,�����0�!��$a��TNW�}�w���I���~��˒�}"�>E��ή;1n�8u}���[�iJW��L})�gn�:0ޖ��>���h��*��Z������������ٻg�<�9N�9m�e={�L�ߕg*'7�l�2���b���...*F�_���?��xzz���DD�A1DDDDDDDD&"���9�3�wZ���b��m�d���C�1�1��t-�Ug�l��aK�-8��k����&]e2�I�icB�tzU��>���?v~�p��X��)2cG�j�0T�T�A�`ڂ8��|���K�5�����:�T�V�]����;�:�ӲNL�ſ����a$`�^�z "�$I����<s�M��RbӹTg��yX�����g��.Ȉx]��������%�N�""������!�E	��P�����/��`P����E��p�9��&������G����_�n�rYz�~q;f4���sti]�5j穭�b��)U�^9N�� S~.���W�2�l#��k~��#"�E�T�Qo޽��wҋ�lCQ���ث�y����]6������������I�\�	ep��]T8���T��\k�9��ȗ*��%�Һ��wodI���yv(�A�"8v�XX��[�5�����&[F�B͐�.)�Ⱥ��[�Z�C�-���/޼���'�yý���w3r�J�,�
�-��$�m�ѯ�.?���������������̗�?�z��<�`����s(�W)�^�w�,�DDD�bkkWWW�"0�
�*U*$M�g7��z0(���������D^EF߃��6��v]�����VYH���r���b��(����6�=0��|4/��v4I���V�^)���k,����:c��6��P�6H��E�v��Q�5�{x�$F���P�s�Θ�h��4�=fd��iH��>��R �GN��\�\��	�Y�z�
�1e�5Y������Ѷ��O��T�K����%�A�Ϛ2+�Z��j�����揝������aI޽��M�^݋�W����c5�}�s[߂�h_���9���S�?Xwv.>�k��95|r�`���&[��cQ�	���f����I��ʾ2�W>JW����W��R���N���k���vb��]j�^{���v ���|o������[��տADDDDDDDDD�G�'6hn�����^�z���'7��� ""2���\\\>	�I�:5<==���%�!"""""""2��U8�j���߼}��K�Ú{�����O,����!5��0
]���SߝRa1kϮ5�khX��*�v%ڡ���0�,)� �e�*��G
y$T���[�VR��2Jv�_��B�$I4۞�sd�'��ĺP�`ڂ�Q��*p����)����펿��DDDb�х���f��+���U�f����Vo۪9��cɎ� �9���a�$tGMV�^���ǿ�x������&�p�\�4�;�9��Z?�傖�To޽Q�%�<s}1ο��ɂb��ʆrY��w��iHS DdZ�^�sp��h�+�Ku��*~���_���(�=�����QF���/�+�`V�,���$�w婕j���f���U��|�7�w

�)dp���6f��~��$�H �Â�����ȁ�&[x6��H��H�DD����I�D#�0Q?�{���(�`P��09�{K��#�� �g���hV���6m��Q���uV=�Z+�ۆm��a1��<� OgO�n���O���W��ĕ��W�_��ӾD{���UXkm��ń����E�M������E�M�R�1��T�0�(���ŏ��O��Ӥ}����b��̭����1��4�{����,ˑGT(Ʉ,���R�wK����Z#�C��޾���[�ޗ�w�F����q � vtݡBM�4-�}]����۰T�.��>?����������}��E�u>����s�à"�p0������V���W�m�d)ѹtg��5?�?���`d������O�X�9�	�m�o�~q{��SZzb��mx{����Q��ךx7���ADDDDDDDDD��ĭ0W�����*�_j�����<_x�hW[WY:[[[�����	���P888����cPUR��������k����ňv%ک����Uo��l��M(�g�h�B�ȭ�R~[�[T�^E�JPE\H��Zˊ	)���O��#N�I�B�����G
���o�=W� 1Zc(��m���ۧr=���:����@���K�]Z״h\��*:'""���������8�� 2�Ȭ����-��Ĝ�s`�$��TB�CQ}Zu��wJ� �bgc_o_L�7�j��^s��N�N�o3���_�_��W�Z��7 "�"�W�Z{�ك�95�IH�bL�U�+캼�C0��]����������6���⃋�3����o�9�i��T��b���������(F$��ڸwGDdjvv,�7���Ӈ ��`�g�h�&""�xD""""""""2!	E����+G۶n޺��u�Ϯ�{�����zz��Tƴ��жx[�v���ǡ^�0h� ��{<����/+�sjLh4�ҽlwU����XM_){%�o9��3�m'�g�4TE��N��'5��.���~������(��G���
��؛A1DDd<w��A㹍���~8�9j��+�g�A1�v��U��:���]�M՜U-:(F��}���|��_��@c�?V�$p$ %2� Y9.uY�;���lS0mAbv��]�q=�*S������uδ���X}�f��wN��u߫���T�Y�N�x��1����������������#lll���{���`�wwwxyy���C�#""�aP��uZ�	�{F
�Ѷ-��$Bz�������_k���k�[�'o��Ⱥ#akc����m85rՀ�"��7x�X�f<�=���a����Q�R������I���C1��Ϳ5���{���X;	�Y�UrV�5;x66�� J8�_���Y*4IK�UADDdL�n���ѳ|O�6��U���+��z
����f�ڿ� ?]
�) K'-��b$�3�[�xr�h�j]�����|r;/�dP��P���vj^��w �2��+ū�/����;��z#�W^���{/9֮;�DDDDDDDDDDDD�D���������ogg��)S~�����-�0��� "����""""""""����bmǵHf�,���3bO�=賦��k���?q��i,n�Xo�N��u�+X��,�G���~���"�-�kZl�էU7�wp)Xh���m'�=�2#��0Y���l��X�z)һ�7���K;���o@	oҾIz�b<�{ K�,�������e��Q���b"��3W�;#b�����ЙSd��[vb�j���%����W�#w�4�r$��y��:�-:��޿Y��g��=͖2����]�_k��٦P�B�!"""""""""""��%K?~�����CLT ��a0�CDD�A1DDDDDDDD�@�U�̬�mW U�TѶ����M&�M	�x��l˅-(5��tX�<��h���z@�%���r�v.I]���"��W�R M��ug�ŕ�W4����.H��%��~�6�mt:�Nz��_�?~��Ytb͙5h��^�}Jxg���Uh���9M#7�X=�W>dI�E2�;��5�+""#�.w��������p����	M^��7E����\]�kvst��W��������w-��������9>L[P�3���N�Nx��9n>��sw��`�A�7�+9FNW���G:�tpN��K/޼@hx(��9�������0'�Z��z#{��*`K�o���e�Ku,���?8v�Z�̙l�r���ΞH�o߽Ž��p��URq���/W���B�4���%-�9$S���վ�ԝS�/Y/��8���Jj�)��0�b�H�.��bd�#�s�G�D��pU��[���q���6ZPL�<�5��Y s��3�:�ʚ*+R;�V��$����S=x�@c��;���ΛM�eT0�O$�P�%���r"��ze���X��U�Aʬ�;j[{����|��K���<��i�B����"Y
Y������aPY�ܹs[TP���-���>�HLT� ""�à"""""""�x���nW�zR�w�hQ�*e����:�kv��E��X�;�G�L�4�IA���K���?��U/��BA��+��_�
	����mUO�k��Z��t}$B��Cq���m1e2�1x����ۊn,�43�!븖n��<)X.��,�樊��+���J�l�]܆U�Waىe*X#������E�����-�}��޾��N�������ͱ�H�~���'A/���s\����u�Q+O-N����켴�LÚ�k��O'�$6hV��o�*9���k}��|�����:~'	�}��7>�}T@�!��ץ]Xxt!V�Za�0	=�_���qR�?~�x�㤈�[�nhT��:�3x�`���/~߽lwdJ�I�4c����gw����;�o��
}�
Y+�(;}�4�G{������`��:۝�u��-��eK�]Jw�?b�p��쾲[oPL&�L�G������s�l��l����m)�����~=�]�3(F�%$L����?�%�3��1���HHr\���:����f���r�2h����c�ŭ*�F�>b]�s��{�PP	��GΡv]ޅ�!�x,P��\��H�{��~��6�K���s���7�ux�?[x���$�N{ÂQ�\ȵ�.r}!��&�4�9N��~ݦ:B�G�X�� W""""""""""""k�'O�sagg�O�`��ԩS#U�T���Y�ţk�����қ����Pv}l:�	�LS�O��mW��9-R�;��@U����/��h�U`p��������)�tX��#跶�*��7��P�T�'��>�_����{�N�C�~�7F뿐B]@���/���0]��'S���P#W�h�=��p���al���w���B5L%�Cr��Vbj�9;;�PLR-A,R<;x6�N�h^)��Ā*t�;z��A1�i�1�w�
�1��%�D)���{��AB�B��M&"�gn����K�Ed�~q;z�ꉳw�">�qC��~��#
�+��e�����F>�W��j�b~)��Z�d�yP���'F���d]6�փ	�P:si���8�q��� t+�M�=��4���S�WL��9	����w:�IhTb��^�;ސ���V�!��7`I�\˘S�Flm8�Am�~�9�_�5(F�$�D	�H(r��c���y����O��2$ `Ķ*�L�LM��6����<�w�<@9'뵪�΀��$糝Ku��U�GF��1�^��$DN�S�Oa��*��������S�	R�k	]$�)>�bU���=<dY$|�髧����=�5�{�>>>X�xq�.���I��D#�0Q?G��2Y�Q�5��v��� 2Dhx(�>]Q��Ɍ�5
�޾R=*K���nSE������QV}��"F}j婅ýc����]�w�
�E��h�1�Ǡh��h��A�Ӝ�w>�}�8���'7���,(�� 2��פ�p�wT��rVӜ.��G���Wdn)��[�o�V�H���>?�cɎh���]�g�eH���fӑ9Ef��[�X��\�y1��	)$]t�·d{��m'���?�e���J!�c�A���t\�OG���+�Ŭ�Y0�\��0��tT�^�(�K�OD�bm�:��*�O���������#F�%A�Z�r�²6�P!k�X/w����p��_|N�%䘿�������:��"AQ�������.�	��"!��@��_��>ײHKX? NǬf�����y.:�	A�If4�����A�Y-СDt\�W]���(�B�WI�_leM�U|ʱ�ۊn�|��V1[E�w�$�N	�j���V���ў���Ix�>�_>����*��Y7%HƔ�M��`�ܵ4�'d�Ş�P_	�!"""""""""""�Vy��A���b�y�������C���sԿe<Q�����(ƶ]�""��ӷO�p�㳤̂�i�GP��L
7[.h�
ݺ�骷��,?���)\Vs�AmC���ά:*(1�B�Ca�� Zm����9u���$�O�w|ě�8Ϳ|��&	���L����v¼�yF���Oh4�6��T#j����4ʼ$�E�%�����0�����y��F����#f~5S����8���$T`N�9&	�(��$�<��ͱ��ćv%ک@�,b*.�>r^���dK�-N˕���#�U��ζJv0iPL�����9��q�g�e���H�Ǘجs�?���RNs��k�a-d���5�����V�ӎK;p��-�7	�Z�ne���Q%G��A��M���N�Ͽ�����F��L�ӻ�G㹍վ>>�kTu�:���"ck����B�Y�T)ş�r��!}����#�䟓�ү�~��ɖ/A�����'7M�� Ӓk$WGW��#��Y��u���������������C L�������]]]�vo������$"""""""�g�o�1�m���,)������H�$$Gzz������= ��>x��+	�^s8W�����q��q�������ǰ(0��l^��آ8�Ϸ�/&6�h�"��"]�
����ʾ�o���7�ckL�1F����Paf?o�٨����wUo�Io��;�cM�5h0����b�歋��f�:,)	b�>�L�;o�UH��|��qh�fPL��Ց�=���$�F��K�9D
�z��W���*��һ��oM����҃K���eЃ\��v_)� ��	��o��Z�q��%5�2d����&�����ͷw��Yo$��V�Z���բV059�Ȳ�ok��HP��n;Qir%�
'�v>�}4��yﱛ�`N]��}t��J��)�bd�Z�:,�%[2��z�{/?�""""""""""]�\������߿���ŉȢȳ^�k�F�p��!���!22�`>���"""c`PQ<�p~��z7G7���䭃#}�����~q;�~���9�3���k �'uf�I��R<;��T�Q5ڶ��M(A��;un���>�k���zq����s�_>V�4�����]��PT�FG��f~5�S1gZ״j�6$$�ڣk8q��<���+	y�����5�+<�=�7u^U|��!9�K���W��4ǟ�sZ�G�_�����"Y
�Q M�P,ڠ��[�����e8LE�ѳ|O�� 58,X}��7�G���$�D�ȓ:O��Vs��$��䵎�?ڠ���=���P<�x�g��� �Je*��)2�^BV�[������0���F����{~O}&��q0Els�Z��9�����P�ܣ�Gj��3���A�re����~��R����vޮD;���t��T���Y����ET��ϱ�J��?���9���[X}f5���KHh���?׸@cu�}��E���_�_�~L�t:�I�ͫگ2($F�1��V�(�(�wM��)3�dƒ��C����,G���T0f\�����ǋ.����'7�k�c����^:Si�Ǥ�EZ�P�!���r�ihH���#��%45U�T�)�C���Ҹ���ΛQ|\q5=����7�n�9^�s;&-8�@���G��|�t�M�*�dD�%!B�(�j䪡w��GADDDDDDDDD	C�.��<�窮��d�Ȯ�3�}n�G��\xp�Ba�ŭ����b��X���g.�~��`gY��3����(>1(��������(�I��;����'ڶYSfŶ��aىe農�*�Nl���ۊn*,Ư�,�0֞Q[������)�~����<�#��o;~����R�`ڂzۘ��PBJd���^Ut&�[ё��f��u/�W>�vN�N������x��]�^��~P�Z�Pt⾉�{x..ܿ`�<�!�9����
4R�ȶd
2_	������~x�хj{<{����r����w�Z��ސ�!Շ`ۅm�wm�M���7����}��1v�X�xrCsz)����hZ��fy�jz��*�%�qX�^���m8Voy�%dN֝=����-��B�2�ЩT'��@�$,�ȟELR�<��d�$u���R����b�=�_���"?/�N��U�~l�)�Fm'���H���m��p^��"鋨�Z�j_L?���A1�}���e�/�A:c�@�����s*D 1��}$�b�?�|���G��Ŷk���&��	r��ػ�
U�)�b�:t*�_?G|���em�E8'�*r��������l#���12�[�y����6K�1&.׮��Scn�ц��9�#�����yH([�h��ɸ_k����7�TT����6%ｄ�I؍�"�E��e1�� ��[Ws~YRf���3�7MH�6�S�u��󛛫���sp�}}���Lr'��
<q�N�>�<_�Js�뷯�FDDDDDDDDD1#���[��}�3Z��|^��h��!���Ig9�L¬C����+��cPQ�w�*��N�mP�f���p�����bFc$�;�{�-ngg4�� �(4<զVÝgw���\O����c�H��H����W�h� ����eY�0y�dT	1u��}L�?SLQ&��F2�d:�M_����UQ��J��������ƪ;&d�'�22L�{�
��^z�ؼ�xQ��(���a�?���^
O��V;/o�\��\
�紘��
� c����å��;�'o��vz)�m6��x7��su�7G7Lk:�g֎�k��g��B�ےζ_��n3h�Ҿ늮j���Gʞ*;~��z�2�z��+�
���|����S����_�#�t�lb�ly��s;/�D�U=p����@_
�eеܥǗb\�q�3���W�Q�.n����۾�v��	$v��W�;���+���p��F��/-�����_�6r��Bv]�P�Ӡ9���S�Gc:b��`1?d>�	�&� ?��T�7Lj<	m���l+�79�o��bkB�	*�O��&�qiG,9�$�yIP٠�0/dV�]�z�"!:r^k
����L}֝]�Ν�Z1:d(a�{g�U�h#=�R+O-u^j�A%�@�ee�jQX{���]s$۱VP�|O5p��Xgj��}��,���$�R��pɾ�����������ܧ��bry��yR�Q�wU��O�N`HODDDDd�CDDDDDDD� ^F�T��{V=t����[�W��7Ɔs��H!w��0�2�g��i8�!�?���F
1��+�o�ك�.R?��t�����Ǡj���Yyje��s��=4e�<{�,��Xd^{����n;5kV�
�c��K��5TX�.���L�QAq%�-#w�T���W�1}��Ja���\��|�B�)U���~��Y��-�-���'���AB�*O��Y�����y�fh�a˰���X��IM&���]s��c��yigDDF�x��SqRE���2���曲ߨ���0i����d�;�.v_����&@��e˺��Z��C�+ￄ�u/�]�4Jv0jP�j�L�� ��L�y2�g��&�F��Y�� 5-���F�T�4��>��F0R�+(�z��H�V�J�t�ys_y�]�vz�H��=�z�h��vq[�zzK�3ii^��:��qib�L�2hV���x�.�k���h��f�)�p���%&�(�r�s����U��.r�9|�p��:"V!��WqrEl�Y�����`ىej0"YW�d��Q�G��I-��JP]l��⃄��o8^�*���n���h��U�L%5��b��:�_tAXs���o=�w���cJ�'^�j���%��ɳ;DDDDDd�CDDDDDDD�@.?���j`s��H�,���I���;�W=�\?{��Ab���t��`�rx���['�Xdpˀ!5���lb�5��K�mE7�y]4��̪�͂#q��o��Iz':}�4jϬ�=�������=s�\�r����1��@j�e�QBb>&�[.l��H�f�-c�⃋�-��z�*��Ez���	O3������̺1�����Nt^�Y����g��c���7�t:���U�x��Qgf����'N��������s�MH�1��;>�!1�H؁VPLc��H�,�
q2�%:h�[{fm����?�/����i
�,�N����a�y�C����Nױ�cv&�,W^���Єq�}&���[`잱�G���]��k�ΰ�����q���ޱ����T@I���4��\�g��a>�_�\'�4$&����ձQ��brS=+���[�����a\HЛg�{�<�J�]�tŘ�c@��}�9�+�9$�KRu��}�|S?_}dN�9�i�_�=֝]s%�%�ϭG�&:��vm̠}�		���)�,-��D���5���ɜ�"""""""""kӶx[�l6Ө�����Ʃ~�T��<������L�A1DDDDDDDD	�ȍ#�:�*�tXcP��Ǥ����wc����a�8s��]��4{e7w�޾Xqr��\�6ߔ�F3B����۠o㵐�#��6=����n�?�q���8/�!1Q$�D�����E��c��5��8)ƶ4��ga�ٵq�����w��v�H�����qhLa��8y�d��1?d>�k ߂�:Ǘ�XB-컶/F����O���5�5$&���H̎�;`����_�
}��5I�Ȉ�#$$����跶�Q�)Ao�a�:��X�W��M��r$ģi����e�L�zW�*9��m#Eɉ�bu��Ȗ*�����J�e� $s%C�mP������f��G� �NWX�i����2��J�]Q5GU�s 9>���?M~��YCs��3k�/�p������g���:��������?eY�n�����_���9^�����Iϫ-E���`J��jځi0w�#�ﾲ�Q�%4V�4_�Ѹ�R������m���r-CDDDDDDDDDѫ��f}5˨!1Q��@����aؖax��-������|0(��������(�IAx�qű�o�ނ>-�7D����cUL�?�L�V,Uݼu��.)^�}kU*S)l�	�N�1�V��z�L�E���;�7F��>J
鿮?,�;�P�7R����9��x~^�^:���3�+������`�>w,�Q���C�&	����ю��@�|��>\���:ƨ^��d��kU/�x��"a-*��8���^����;�t��i��=�MB�,�b��d=�#d=6FPL�"-��>��q7����[�XI�ר���m7��LP���6ÎK;�XH�����"鋨�CB9%TF�'J�U|iW����6��WO㼜篟c�����|�f�?��پD{��#�E�c�1����{����d=�0<]�5Ϫ�Fn��2zU�쩲1.kʬ���v]�2�7��`���m�
"��oP�()���b��5�� K�/��rj殩
	t��]	$#�!���Z̃���f9w��JDDDDDDDD?��ׅ~M��|/�C�P m4hn�ϽY���/�����V��*��*R����^E������7��A�f9=r�J�*�TRl%E��C��Z
;�>��ܷ���ܜ���e}�
X���M`�)��v�v�*�G��ҙK�N�:����A��Y��n��%��m��,
ϓ:�z����{�/y��:�����&후;��e^RD����1���^�%`*s���1��:B��凗1;x6���s��C]�w5xy�K������&)��k�ΠQ?}��H@���7	R9|��I���b���O�$u�b�M_Go��2:��9n���0����p��*�+:F��տA�#�פ��0��T��{���s��2)�R|1ο��
W�G��P1]�Z-��úr͡E�ӌy="��[��
�ŷ�/���n�C�Ӵ`S���.��{�a��}����bm��0�v��i�����zz˨˓mw잱��Xw`Y�|�c"�%er�v��]X�&��X��e��/�=cŴ*�Js�ʵY9'�����x�����������(~�Q�����{,�1��g�U�����e(�3�^��N�4��ب�Q�1(���������L�MX�����X�j�f;)���
~��޾��bH�!���쯳�T�EGY���6am>�[
U�7��s��M��X�i]N�`ǣ��m�d車bbc��1��o",����uňi
�������I���/a#�bѱEF��l�i0F�>\�iF$�5cy����iR��#� e����˻��������9^�LA4�>���)�~1�\�rjۗ���@t�ɕH�B�l�R�x,]Jw�9�C�8�����TR�8	4����"�C���婃N�:�����{$ae{����7*�hىe�<+Q=�)�	�w���%����?��LK�B�t���4r�/��F�4�����;bJ�%����G���膲Y�b祝��+�W>����'�!���=�6O9�j���zߘ�;�k̿����>W=Wu�iH8�G2�M�W��]|�DB���b|r�������z�r$�ZdD��A����z��X�C]s����ʋ6���m#�bM;0���f�]ґR���u���}}j䪁-]����F"""""JX�]YCDDDDDDDd�v_٭�Ȥx^)�\m������1
2�T�=sï�,]�h]�5��k'���0L칲�!1�@�fa
��"�wM_����9塚��_��.��Y�'z��Kp��9��}ʨ����*���t����Q�7�۠B=�i�~��dtϨs���Ŕ�X)���9N^��[a*��t�H�A�t�p0��Q����*DDF ������j�.cơ�A1~E��om?�z�*V�-��Xr�m��
���6�-R%O��/g/����h#�����Aq#a1峖W��4��5Z�%�s5	-е�˾�R�Jz�N�_�]�w�Ɠ�/UsV�'�.�fl2ϑ�F�)Q�)GU��b*e��9N�*�GL�9��S+5��!�Z��<���P�B��pu�&�����ʏd���؜�5�}+�U�IC6��gwa	�����+Ȗ*���8�U��0iߤXϿ��c�.������������5� �5@ ��`c!Bd!hwwwwwww��=w�����������٧��p������nu�����L��#�\����
�C�9et�і�S�ɻ&�譣      @����G��ͨ�7OKPH�쾰��r^>(���L~^����g~�r�]����2�=�v���   DA1      >�ܭs���V)�����
�)`~x]r����w��gF�,���5pDW���j}e
o=�%QQ���䃊Hろ%F���~�@��E���?0�"��Y�Kڄi�Z֦S���o;l�V��l;��/
�����Z��q��u�M�4�FG�r���P%{˶�G������S��оD{�m��-(f�i{�㮝�w�;��U[�l��vH�tE^i�0�FɄ�^n��X�!*ds���
Y*xt��vN�o�|#�W��ɥoݾ�0Ci5��_��j��u��	m���*���e.�M�g"��kH�8�/�~�tz���T��m�;g�R�sz�Zw�����h(��9��'�y�QP�^G�w��s�\\*X��/�&��Ň�������L0�#z܋HPL�bm,�4`��3c�A��e���$�疮S�
      ��7f\iZ��e�ѫG�ʠ*nfp��Uyk�[淭�M�¬MWTV��Jj�a~'   ��      � -v��NG��IG'�~�)P�QA��w˾+u�ԕ�"c�2�� SpU$��@�o`�+�QGtqOL�~Ϟ?�!��ЍCM0��iQf�TyMA{���$0V��4Ò.Q:�6-�sǊc+,۴@wT�Q�X��%������
k4���u~�e[�$�%~��r��][���p��9�K�ϥeN[ز��������"���xCd�W�}zwDâ�S?_}ss����&���2B�L�b�MN�7�:# �$��X��Of�E%3�4Ǯ��Kg*-���$�U����KT�,4AC����0�K���x��=��{�D&g�#O'���ny�?u~����9+�蟄�����}�݃b^�# Z�$��P��K&�S�b鋙�Ύ��������~�6v�Xˠoʞ<�)(pW��i�Z�j���6V��4qQ�Ef?�r���R��      9j�i��v�ᓇ�ttS�Bb�N�)�k�j���J�TydM�5Rmp��b�	   �     ��Fn)�V�ԭ��LI2Iߺ}�:?ȆS��SwO��/��ґ�	�E���EZʂ��(,�J��5��E�R'Oˢdg�_���b[���Ѣ��|퉵^	�ɐ8��2YZ��+E.����h،;��Ro������<�
53��v����B�>������r��>g����?}�T�]�'�����s�s��:��y���+�œ�ܽbٖ6aZ[֡!�^'O������M�DÍ^V%{ɒ4��7�u,�ѲMC+<y �_7�ߔO�~"m�K�֝\����֩T'�\����@�����R)�gy9~�DeV�	��$27�N�9镶6��8\֬�����;Y�|�#E�v�CQ\]��gگ
}�t�R�l��1^V�x�8n�/+^�xN�]>$�t9��e�]�yv����kJ���>Qzs�~��;���z�4�����-��$�j���¼L�)�������r�{�@�vv���i_w��s�`�����O���eυ=       �T�i}_�w˾��<��V����Z�H�j��������VK�AU���#    r     ��tt�6�ۘScDw�+�qVt����f��{gȌ=3�j���a�ĉG���M˩�d����/��R�a�o$�s�vX$�*��sݟ����Z����jJ�`y����ש�0�Wx_�f�jy���~���o�Z�jan_�,���c��ܭs���BYvd�	��"Voy����|�#˾~�	.K�0��v-`�#(������w�:�F�s-�<��+"����hȁ���۲�{�����^��p��m�(�E�ۗh/_.����i����f%ds�����5l�0黼�\�sQ1z� �_W�*?����X����=���8��	努��&�)�敠�ҙJK���Y4t&2�<V@,�vO���|�i��#�o� ��X�k������\�r^�^��y��Ǖ?6����,d6Y�d{���,�F� �(�7w8����l1R���.Ǯ_6v�X��<ޠ� ��o�sɴ�����<y�D��in�a      D��K;�������umY��?�ga�ua��h>��1��{M�5R}Hu�{q�    �<�      ���6H��-d|��N���B������'s?�_V�"�NQ�u]fF��t�y����Z��u�T0�Ì�^ֺ�����D��o�ЍCÜOtS�O!���lɲ9-vUoK��M"�G56�b��'U�t�-����}}͉5ft�>�����t����%�6�Ҡ�Yvt����*�Eo�d���X�hȊ]��[n�p-�u$�����: ����xKx���o��0��=l�0�A1J�b����s��o�Om=�Uv��%�;=6�9�F��.SvO���o
쥣v��՜�F�e�Oj��{�ߓ�V�&Q�UhB�\�$E`��	�j[���e\�sIZ,�)�s��{W=��ºtۜ�$�*0���{��nײ�O����Ů�<���7�}��5d�����jC������WM�5I~����k}���h�J�ߊ�+�M�G㶏�.��m5֜������s��       �K}ț:��6�=�ڽk��oʮ)r��y��i���4����]�   D2�b      |ش�ӤFh32���]1��<�sݟ��4�bN�9� )��P���ሆ���J�eZ8�ӊ��W�^榃��b"+�h�G�����ݫ�s^O�����H�U�H��On9_�|���7��.S���t{-�����/}i�v��	��!q��~f֟Z/#��47�h!�'iP�'9���<�����'���a{X�!Y�d�bǈm�r"3��uGbH��Seυ=R M�W�2&�(5r֐E���=�v(���=ds�Dڇ+�JC�4 �Lnʍ{7�쭳���>�wi�<~�X�yZ���\=�Z�Y��\?У�b�6q�D��	���5�����0�慛[.�S!zVc:m���s�Ȱ�����o��s��=�'�b��#Y|>��s�ǫޝ���O��i9R%{y#�2��|�U����B	��]�	�	�iS��e����yZ���o:��`iZ����>����F      �4�E��Yqt�G֩�UTUu^dy���Ŭ�Zj�iD   �y�      ����WK�~��*�J�r�%i��.?VG	Yvd���6����;�N�:f��$q���B�_�e�)��uկ���,�#3�͔�R�R3gMɜ4�ˏ�"q���M	����]�W�l"C�qZ,ֹtgYr���:ʶ��~��o0���q�봮���v���O�#*�B�{�����G�?d���������	�qR�'f[�a7VA1a=���'D{>g��oy��A��oئa���v�ֱdG��b�d�b��vL����ؖr��9��k�_� _��������)�E����}��Y�&�-���A1�`6f��la�~y2�+���81���m{�P��)vń�������D��z/�-+ޱ���V��O�(���*(F�>���K�m���*�ʲ��F��Ǻ?J�R����oU?�y��      �;��WP[�z.�E>��,�DR�p8���(x�	��vv�    �,�b      ���GwMȆc����P)k%	���q:r��;e��=>7f\���&'z���=���'�3��3{ȥ;��W�r�L�s�s�ˡ�eƞ2r�H�xj��?ݸCZ�ma�I���b9߀Fd��Ur�����R�J2��@��Z5dér��A9}㴜�y�l�7=}d�+�$��'�;�O�q���;��44�jD'W�����<��H�o.v{��x����q�������za�ÿhA��j�e������L�=Mn=�%�7h �8Z���Z$*�(3p�P2cIə"��kh�#�/���ͯa��<y��>�^oZ�31�o��m�����=��<��Zyl�쾰[
�)�]���$L#n__5g���pr�7�kP����|�򖁲zM6u�T�o�Y��|R����2R>��|       ��l�+�W<��]�wIŁei���.Q:��� x˺.���js�   �a�      ��Ї�2x�`3%��܌Z�?u~��c�{�ߓ������eѡE���9p逜�yZ|A�<u����%iy�i�m��5̈���B���`�7U^)�����UK*d��(�e���̌4�#�����}Fwɞ<�T�Q��<z��x���#"�Ĉ#ÛwZ0�E�Z�=l�0�qn�<y�$\�J'�x�ބ�cF�nQ���.�Z�f.�P*�Y���TZޝ�n���#��œ�N`�fW��������<�ｂ�i�֔]S�]�v��iX@�bm�5X>^?�oxӲ=ds� �r���rf���X�a���4�QFԜ}s����Ge����V�&���s�X���Cz�T�J�X�~��^ga-���$g�w��'��Y~t�eP�~6�e.��!)����vɷ�k�ƕ��ϊW	��M���;�GC;M�$ϟ?       ��(�����Vq�2��	�ɐ8��yt/�:Ցu'�	    � (     �O]�{�(;�yA��g(n�4tF�btTk��޻j�y��e9{�칰����J�*I�j�����?Z���J�ҝ��eߛb-O�jQd���LH���20��R�OaF~�I��]Z$�)���(F��c[ȾO�Y�&T'O�`~��\:X�&�jٮ#5�D��:'� �=��a����8�L������	ܩ���)(���2�Kˣ'�L��]�*���5����C�8	-��zZ��L�&1���6s�:���4(�e����kұ��j�i����A1$�#y9t�DUzL�~x�R�^i��s�ϙP��i�}��q���V��îݻ�u'���i����ϑ΂d�ƈk�J��������<��)��]fAԵ���G�X���TƧ�b��\Y���W�|V�<�c�x=&j����{'D�i���7J�h�,����V�Z�      �=}d٦��u_�����ʛ�p��]jq��Rx}Yvd�    �A1      ~l���ҧz�������yS�5�����К��h�PP� �G���aM\&��d
p]��L�9�֑_����	�	Ͼ�9��x�ޥaR��XF�m9��D����p7�-��e��k����N��ݡ��M�+�3��ґ�*d� ��V2Z��3�^��V��l8����tO�8Y�vמc�'���ǋϲ=���1<s�̲��N���cҁK$O�<��i��m=���c�
���������x��+����N�:J�(5p��v_����c4�I�8�����N۝��#*Q�DNۯ�w�m�Ρ^�76{*L-��W9;�k g��1L�"��ˡ���[�(�K^�2&��J����,��:���urױ�����|K�<u͵���O��9�M��'       "ύ�7,�t�������~�\��
���Rɗ:��y����gK�e��%   �^�      ���W������
�{d�@ѐ-��ѳu��EZJ�xI�˕"�i2D~o�L�3�B�8�B<y��n;��+������s^OAԥE�p��&�hȑ~��^��
�S�vئ�|�Im�Q��y���?�L*M�4� _i[����\6��S���k���ET�q$y�䦐�nZ|�6aZ���w.ڲ��ҋ�貵X�JX�Ao���WC�ɜ4��<OP���i��Z�W�mz�t��I�rDC�a��R�%��I�F�>��&��qJ2%��J[��>f춱�-n_pڞ!q�u~�G���5����Mϑz�iV�A+�
�I�؞�Ù�g,���K�s��IA�VP�?|������KϪ����k㴏��V4�֎�اr��2�������m�z!����{      �7ܸg�20������,z�D��UeI�%�~G4,fN�9�lL3��o�    �A1      ~���^R*c))������"_.����iq_�Ty����Y�L�����ƌ+���6��hX�e������n�G�����?�}S�nW`�����i���+�Q��Ͻ��u��YΣ�%SvMq{�q��5o�<9r���)K�,�k��z���f� 	��V�Z�r��ɲJ����m�i
������hٮ��v���x�ҝKb7}m��|?̑���V�ȳ'��=g���3z�h����44�������:��h����� D����j�4��>�����˥���>u�T񖻏���{�-)4��E0�ݬn�U�뼬�2z��@���h���z��`N;h_F��P���s�Y���/߉��6�2(�J�*&������󫛧��r5l�C�C�Q|���\: ���6��       |���o/�b��V��'�}�W�ŝK�tEΣ��Ln;Y��nj�W   `�b      ������+�L��9kFxyZ����Oe��N��?2%�$��7���'el�0NB���k�EX/
�t�vv�)�<x��)�9s댜�q��Z鿶�l9�E�7�/�3��6=x�@ޛ�	BԧEfP'O��^ҡd�a�[�u�1s�L���[v��u�A�����{�߳�O�l�I홠g�ZX��	�֥��A1Ξ�{5&,;����������'����nBa^�(N"i\�������z���Y�<
_��[΄>
�ׁ�&��7�z��~ߥ}R!K�m��c�!4V]>�R���K�-�b��/��;en�Ӗe�>�c׎Y��sV�Ň��d�9mw����s���v)���+m�L�ߪ~��5)��ah�Ұύ�6
|���w�/	b'��G��j�!WB�       ����cs_���f�g)/#����m�z��	�Y�PJf,�p�y�[S�Ř2c�   q�      D:r��ސ.e�H��}�(��u���Q���6�����($��M ��8���ΊJ�48FB���y��5Ġ�27��4�_�$��3����oƈ����'=�����
^_-��2(F}V�3�y��I�U��d�l;r��)z��7��=0�)���	�r�b֊���D��	�^k=v�Y<��a鑥b7g�aυ=.-c뙭��֑
Y+����_�m�0(F�]���	�i���e1���L��$L��ƽ�:� 0=v����2ަ�#���RKI�h�L��N��2��X�ﾰۥ��k��#�곕�`�r���jS;WmȊ�)m"����S���[�(�s�,��� x��<먾I�%������RcH9w�       �M:@�UP��ܸCj�)�X�n��Ni7E�Oj/�<    CP     @�E�����GH���]�vR%{�Q��xj�vo����l;�M���.�n�2Ӆ;���[�����Η0��p2&�(��d�lɲ��}]�m>2i��'B}��<#��L���!.$ j�rf�,>�Xj��=K�,�`Нъ4��ʥ�Kb'W��+�������j1�a{D��^V/o=sް���p���Z[�ո`c�a��.S���rղlw�98��#�Y�g����V��+�M���*e�d�Ǯ3�ݱdG���:����*l��׏��B`�
��zEZ$ަ�w˾�M�mJg,-Nm�u��L��9�&W�|V��a�K5d�ڽkb�&�����^*-
�pئדY�e���^����DC���g1a����O�d��+"�R�}�����آ���h0ո��ާ���.K%U�T���1V9^�[      ��]�w9����s�� /ݱ��W�y��֒���[��D���Gr_   `�b      ��O����Ǌ/�rT��%�K����u���#Y}|���?O^$/4EJ�z��R�50�v��f*���D�M^':�K��}e������~���A1�󪟛��Ϟ�+��1D;YQ�*gE�bbW�K⸉�{:g��K���${����;����a����
q��s��쭳�>Qz��V������/����)�~��:�� }�1��sT�\�����z>����e��	��>/���;'J����&�}��O���8��O��SZia{PL�����/?�ܥ�9������>�a�z��K��R5{U���sM�_�h�_i����ʟJ�i]Q���V��4P�_\�sф����)�F>�����U�V�y��BG�/u�Բ��ɐ8��<�ܖ��j�O       ߴ��:����W��S׫�;�yxG�����q�T�V��<�[����    ���     �(���{f�u��u�E��O��Q[F��]��H%v� -^ԩ��ޒ1qFi]���tD��A��I�J�*��|h���H@9S䔦���iW\�wݲ-e`Jۊ5��a���O�޽�]���Q�Ju�5(�s�Ζmz���Ë�n����缞�-��s��#W���=O��>N>����ҙJ��O�&�Q[Gɷo|+�b���V�����_��>�Bj�_����! �ﳢ�~w�����&��\�r���6Z|�<h0C��e��˗�����oڲ>���eZ�{q�����ca�l���
���!��{Ktt�:B��K�V�Z��<���oMh���y�;ET�O�2v�Xˠ���D4I9;�r�]z�^�y��H��r����K��e뙭      ���wy����G�2�-����>�:Ց�fJ��5   �g     EiȐ&C�J�*�i8� �[�O\:)�<}����3i����7���]l�k�Xl��{�E_�k���Ϟ
^o�-�NtZ`�ޫZ/��k�KE���P�e)g
��0��&Xş$��ܲ���Gr��]��U?_}�����>�:��ʛ*�t,�Ѳ}��Y�0�n�O�\����y&��j���T�R��]��1d����'��!?�,��Xe[�"�ވ��s�BM_i�p�7r�!틷�|�� �@b����t�y���݄v�/4��*(F�Y���ќ�lY�W��r*4v�{!�vN��)���	 �#�R�U=��(�w�����#����O��i.��ƌ+���/��h?ݎ~ud��w���?0v�+m�[!kZ$]��\�F��4�'a��� x�HS�r}���nb�O       �A���Y*���z�M�mȝ2��|P�I�$S�M�zy�	    �E�     �א�hz��}L�RT�-Zp�wy_9��׶c��ufʔ$�	��P��߅P�#~���/���� xJ��8�C��Zxp�l;�M��/�]��4hC��r��i˶&��/+����V���X|�cW����_�~����ʓgO½�hѢ�c�� �?��)����� mƷ��r�Ĉ#?��Ѳ���n|��~B�o/m�9޶�i
J�F�����2l�0�A1����9if�m�ܒ���
`%i��r��u��G����Mv8��b5e���� ���|/��$r�޽|ws������e�Z���÷�7b���hP�ն��N�C澩��$��X<A�o����|�H�B�L ����MC�F��4�C�u�����A�w���Ү�㐬�E[��X�Z�`~����U�R��C��w�Ή�^���gw�-%2���G�ێok�+       �eѡE�bT�bm�����m��b�Q�eJ�)f�"    �"(      
ɟ:��k=β(-*����.Ǯ_q��)�2�����'3�x��-LPBT�� ���,?.�Q�Z�U�%�߾_��L{k�e{�j�]
�Yyl�|Z�S�m�2�2/���
�vV�ZQ�4"vK?����wZ���^ۗ=@���nپ��z�ש���ӺJx}]�k����e�lm<�Q<EW���"��#\����Q-GI��,��m�\�������ҤPD�Hp�`�y��|6�3�C�^Ȗ,�|V�3S�z��aA�-;�L�_;.Y�e}��*$FM�1�* V�Y㟦���/e�I���*Y�d2��$������4���v��m�~�����a{��X��Vn@9s�	��3Ȝ��8��"WB����;� P������z�ɨ&f����X���p��������N,��w�K�P�u�ǶC��W�X��n*��~B��H��5�Χ���W�,�HC���b�l*���iY�����Zڄi-�VU��½���J�*YΣ��~5y�d      ���gX��_�vɷ廥���oк���4��m'   ،�     �(@�H�-����e�yD�H��o���o�����U��I���H���$s�̒&a۷C�Xޙ��,8�@|��״�J�nj���'Q�������������!0�/헼��:l/�������0?�������E�4���+Ԣz��2��L�+��ME4�DGk�������tz�-����u~0žVf�!�ХLs��f�7�z�X���O�~*��k�_�❋2i�$���{����Y�f���}tW�Z�U�������gAs޶�I�O${��<9X�ݻ&v)���)�o^��	!
o�^�� ���߹�8}=����b�y��=0WB�Fx�z{��[�S��L�3@��p�}?�����L�]�l�;/�z!��<�p���%}�����⿖�K�C�=�t��/_�(#�ߨ��������A2��`��y.<�P�n+m��qخ�ߑ�G��W�SGԴ�>��٫��U?7�gگ���=��S����GXFn)������rs-����%������)=��?W�����Zz��̇�?�
      �1��`����0�W�4�����H�U���� MF7��m&ʛ���cI��لg�zL�x)����   ^o�      ���qʨ���^�ߗu'�Ɏs;d��}����������5Y�e1�1E�1�ڻRLe�M��?��(62�<�R��VD���y�Z�^O�=�37Ϙp��w���+��O��'�'Q�D��2i��毎r�Q��Q:Si���i?������
�.-���񱭬G��@���b4xc��i�#�'��L�t[#oM|��B?���^:��l���Ϊ�1��8�A�f�c�ĝe	r���p-O��YZ���C��r����7�9���׵���)s�{3�3Ǟ��1^�m����t���������n`�����Lh=����^��9��ECδ�<�Ѭ�]��ه��տI�ܵM��-�����X7����8�#yi^�����/�[F�ύ��B�Ƿ��*��j�i&=��͟P���v9x���/�B��d��Qm�����3���O�}*�n��>=�<�c�r��<%2���l7!�s��qi�z^�x��N���|=���+�W$<�\�aj����<��ט]�v���¾q6v��&<�O�>�\���w�K��=�l沒5YV���o���GҴPS�y��&���~�#%3�4�v:�5 ^�-Y6s=��o�o���T,}1��%G��������P`����ԑ�e�Z>vʮ)� Y����J��=nXɖ<����׭����p��=�W�^Ҥ`��yZR'L����z0      �^c����_P�S�q���c���ci6��	ҷ
�]��
5�;bō%    A1      ~,g��2��Lɓ*O���A�0��|YulU����N�e\:`&]��w/�����zp�N�9I�����ga�!��dr�qϟ?��+���C��䍓r��Y���.y��f�s-.���T�V�x��M{k�|��;�rї&<��|j8�a:R.s9�����8���r���_���*XItZ ˎ,37����r����GC�*f�hF"jR��	�y����c�?dr���	ZL�M�o̴��N�xj�	��zv�9&>z���h��#�p[o��������Uxw��q�pr�+!/�S'O֥�[�}�5C�oろ�K�.aTiA��xsM��U��o��~V�3iS���0Hf�!�����M���+j�k���5�pj�����m�#��n*뺯3����q���*~ K�,5��5�ט� =?���/I�%1�C-f�I�'�A�p��	\�0Wh0 qc�5�]����5����&$D��W��I 	c'��)$O�<�O?V|��7j�(�a�����5r֐���ZΓ.Q:��q�l>��]�9F^\j����r:��(�3s�SwO���Fh��|ݨ@#�aj�79��A�u�	��|f��S��u�.G-]�i�F�=߯��M?uC�� j�ߨ�|Q�Yth�ٞ�'�ʹ��^�y[?��,��8ϗ�Tʄ�9�w]��������+=�X�83v�X�4��C��v�Ϣ����sA1i�	s��<���b��T�      <a���r��5����w��y'��5�I��h?���W�]�v    b�     �SZ�7��I'Q��q��=ST7h� �vv�x�����OH��z���~�gZ�W�&H�|��aο��n�5�W�׫EKˏ.7�ٓg�7r�!urב��+�D�d�@�BiI˱-M^d���ehS�����z��!*HҥL��U�Q�L�❋r��u��#�;�	��t�w��+Ǯ��P8ma3I���7-���Q�n-d��_8��W��4s�L[��ׂ^���Ad��-�I_�K���ҝK&t U`*�`��i�y�Q�M�'�O	�-�oy�([�῭���t���cd�����;i6��-=�:�ZKw^f��#�50��<�ݽfn�Ҁ;���a����㶏����`(��6k�,�<����t����h`�3%3�4�zS����ԝs˖3[�㤎Qz>o=��l|o�dI��r>=7�S�3)�~�n���5�Ί^���^Zm-�r��Ay�7d~��a�O�O�#h�}M}������1b
|��1k�-{/��aJB�c�:y���=�V        ����oxV���(�F��8���>
�RK��n��v   �날      ?��lÛ�X�����׎K���e�֑+�Y��	̨���BC�т��@�G���$�Y�� :�����v;z��y�u҂��%�K�2]_	�����A���2������Q[G�5����;l�`�2��ȆS�.��Y�ҙJ��^-��U�,�FFo-E�o	�h��3����a7v����^�f'����<��k�?}l��7��,����c�˂�������;4�'hx���uV�˪8��Lo?]*d���c�y�r�ȱ��b9}�dL���|3���ɛ��a�����S��hJݿ�����.��TX�&�l=�Մc�yxG��Nz-���r��u)S�),D�ab�y~�G�b��{*�YQ�t�cB{�;FlI�0��,=�T�Mhg������ʏuty~���       ���.�F�b�M�&    "��      ?�A��_P?S��.���%����ͨ"���
�PWm:�Ij�%�ܒ�D_��&�e�v,��r>`�P�%��xt{4��տ��k~�j٫I��=�~���,[G~Y�}��R��#���������~���O�>R7����<|�P�j,�;/�|��ٶ}Z��������:�}��g豢�CWI�!�e~��.[���rlK���D-�m2��Ll;Q�Ĉc�2��W���v��4P�꠪�Uͯ䳪�Y��M��4����B6��׵�v:_��|ե;����2e����*��HH�iU��G֡�I���M0���_�/�U6A7��d�e�z��4��L�5Y"�>�"����K�"-#m�ڧF�8v��Y�G&��BR�o/?���ٺB�e            �Y�      ������n?N�4X໥ߙ`�Ȗ9if����.Ͽ��n�9���~p[�"-��,�bI�bm,����&� 2
�t�.��e.'���3A/�+E.Y��r�4����uN��8LzU�e0�F�7�h�����v��9����_ZB��H�B�"�]��u��E��'v}*wN�Z�j����W���ޗ���m;�M�('c[���`�Ž�|LsS$�f�e�Wƴ#ْe�в���v|[�x�x���Y�G&� ���Mj��u�v\Fn)���"��C�o._��B�8l?q���8�B WL�5U�&L+urב�؁]���Z?H~X�C�틿�<y �ǵ�Y{g��0��v�zE>�����>N<���R���2���Z��yF:L� ˎ,�Ȧ��V�Z��^�HS�c��~܈-#L�<G�gYpp���:��;�:?*:{��h�mX���b>�            �,�b      �Ļeߕ~A��~���҄�x�HkQ_���\�_���B��|a���H�Y�e1�,�迿U�-�ed�nۺ��L�2&��o��&�'"4�ay��RyPe�p�� j�������73�#ѢE���{K�Q��\����B&� ��������=Z�<x�`鷪�)~�}�z��=�T�ZA��+U�W��i
����Ϟ���Q[G���S����Y�^=*����e��'U>���3��x�����'�s��������)�ka���ҭ\7I/�[�?t�|��+Y�]�g�Ҋ�/&�Wx_�o(	b'��25lׅ]���b���ĚH	!{�iQ��k�$g��۵�?���~�7�)N�8&D*(_�T�RAr��m��u_\r�9ߎ�6F�<�#��&�l��}G����~��\?Є�j�Ӯ߻.F40A1���/��r�^[jP�n޿)ޤ��B��ڹjK�rݥz��&@4"�����Fs���o�׮��*���F��z̄ jS��wݕ����c]
��m�            ���     �M5����w�0Č�~��}�j~%��Uvi^-R�Q�O�<-��\�2�|�GR�p8��6���*9q�D�n�L�9���o�_ڗh��i���N����#���u�hd#�=�ö�#�e�/��c幸P���̽3ͤǒڹkK�lUL��Q�LC[]>$Om�Ȓ�K������I��88��3��M�<{"+��0��+���PB�d*c���s�#EI/��2t[w��-��m��g������ܭs�-���|��!&��~��R.K9ɕ"�����M߫�7N���M���s<��������W�M�9_,�B~Z��	�	�$�2��,I�����=r�,?�\f�a�z+Pe��m�nB;�#�T�^Մ��X��K�����k�!?w��A�sq��<�R.ݹd�v��������x��X�/�~�[s���� ����$=����O�vO�t��~���a_��s�[uR��`��鋛���y�Y@�#��>���Å=&�`퉵r9��Df0}�t���&���_r�[��VC�t�����T�ZQ��+��'w�j9p���.Y|x��9��+��_���f�7Mp��>�n���'e�٭����cy,�>��˾w��=i?U�Dq��m��eM�DC6��������iߥ}�ߨ�y���u��y>����M��{ߙ8�����üEC�f��|�4���V�jd����������l�����x���{Ao����           @�     ��Jf,)�Z�r+$F�ޚ��L�=M��fΚҫZ/���c��Xx]h��{3ߓ	m&8lO7�Ln;��h�LdӀ��:ȢC�dp����1�
�-$�[�7�&Z${�R ��mܸ���j�N/$����&�����ޣ{r)�����zb;_�c��۬4@&0v��
��q��NC.nݿ�@O�`���IiA����k'F���9�y����m	�����`�t�S'Lm�����	��bF=��(&A�c�$L#�b�}��>�Ź�>hѴ'?7�Df�qDu(���MC��<#Q���Xr�*o��v�z�aj�0NBsl�c�#�8����c�2}���3��7??�_Ґ �^о~���̾��znѐ���o�/�P:���I�'Jo�Y�u�<x��E��Ru>o�j����'J����2}��1�y����aOo���z����4*��uSx��6��S�=���5%           �A1      >L�f��i��\��|uC���Sśt�Ǵ#ѣEwi~��-���;'J�R��Z�jۋg(.��"=f�o�m�tz�Lo?]
�-������hF�"J�:�S�������Ұ���̓�O�?����A��XҦh����!x�J��KIt�'�'9q��D%�O<~�             �#�      ����2��XI�0�ˏ9w��VK�]�'ޤ#���4_R�t�1�^�o�+J�ӷK���Q��u�u'֙�o��*���쎳�B�
�^·?�U�Vɜ�s ���y��"0�ö�w����s               �b      |TϪ=�R�J.���I�2����M�bɴ��I�4�z��mc�u���J�}a�LS�r�-F��[ge퉵�-7�ߔZCkɔvS�n���ZF�h�dx��R�_!9��  ��(�òmĖ���C               �      T<Cq���W.���-�7���Cb4 �fI���z܅��صc򺛳o�Ӡ�81���3�\�rr��!����K���d|��Ҥ`�p-#y��2��(�9��<�\  �
�d*#%2�pئ�a�	               ^�      ����2��`�ݵ�n�<{"��4�}���}[�[i[��ۏ�x�@d�������ϙd���N�L�2r9��x�㧏�����.Q:S�sT�VEZɸ�� ���G��m�-�#W�               ^�      ���e�J���\���Y��co���gҫZ�p=6a�����κ4_�dYeN�9RmH5	}*����i8��lzo�dN�9\��%�����zpK  �gE��f��Y�\?P               �� (     ���L!������'�$�o�Q�����7܏O�(�Ď[>y(�3w�RJf,i�b��UW�=�'�r9���u�ׅ+�'u���u�����!  ��x1��_������w_�-s�                "�     �!W�X�M�ҼW�^��f�'�֡D����ZF�q�t�Ҳ��*y��L�����U�YgIPH�<x�@�e�Ž�cf�bT��N�w�տɩ�  ��w�[��"�X��͒o����               DA1      >"E`
y��.ϯ!1�C/�7�)�F�j��D�=��jU��k�+E.�S=Gu��n�4�X?},�2z�hiQ������+ �|Z�S�6��  ��l�?���1bK��TR&S�����o+;���{�               Q�      ���+},��]�w���2a��&��|�-!1/��{Ao�z������������K˱-�ɳ'�-]�v�=q��طK�-?,�A��:+  �=�j����>{*��v��ϟ               Q�      ��x1�I�2]\�W�?��xSp�`�d�m!1J_��� �S��u�!AM6��l"�[?���[�㧏�N�<-=����ot���cĖn����?  ��~����3[               �A1      >�y��(N"�杰c��zD��G��G�?$Z�h�/�cɎ2q�DYvd��n:��,��&��2�j*qbƑ�����'��n*�Wx_r����c;�� _.�R=}$  ��9��H��               �A1      >�k��.����S�n�w�-�T�D~���ǖ=Zt��v������v\^i��/j|a˲������4<HB�Jd�}��e�˨��~l���~��2u�T ����2B�M�&O�=               �.�      xY�4�dƒ.�;e�9x��x�W5��/k~���$��T�w�/UU��/HT+ �Lh=A�Id�2+g�,s;Εz��y%,f��qҧzɑ<�ۏ.LP �/=�\�].?��YZ$               ���     ���<ﯫ~��=Zt�w�K�r�"m��R�﬐ZCkɩ�$���vhӡR)[%ۗ��\�y�����ܸC"��gO��e�ˈ�#�~l��UMX��{����<�#SvMq�v��	�ش��$F�WV��յ{�dυ=���Z9{�                �BP     ��5�����]9$[�l��;Fl�r�4-�T"���l~�4�D֜X#QM̀�2��HiU����Q&SY�m��1�H/\�}��T�'I�­�i~���d����~n_�fc�	 ����5               �*�b      �(S�LR8ma�����Ȕ0NB��~�T�^U�%e`JY�u�|��[�~������
�%J'�[���Y+z|]�S�u=�I�a����Y?},�wM�n庹���                 ��b      ��^�z.����s�}�D�T	RɂN�H�"�m1b�׵�����K��e㩍��Zn!�����G�:3&�(k���z!�"���c|��bj�%�bɣ��                  �AP     �U�R���6��$Ǯ�Ȑ;en���<ɚ,���b�����eҮI�υ���W��?)�����T�Q�+�O/�,�L��n*�̏�un8�A�_;���?V|)���߇                 ؉�      /*���K�-9�D"���Li7E��M"�(Z�hҢpiZ��L�3M~^��l=�U|Y��e�g՞R/O=���/f<��a��;�]�i������s��s������ǖ�\��                 ��!(     �K2&�(��wi�u'׉�u*�I�9Pb�_=@�jf��v��-#e���r��U���2�\*X
�) �$F�2��Pə"�|6�3y���G׷�Ȳp�h�N�U�                  �AP     ��h�+�>{*Om��vD�]���+�T�D�Q�tE��k�_M����se������~y��y�l���6T�VE�o e2�1��/���ǒ=yvi3���}t�c��tz�<y��Ը���                 �날      /)���K��Wn=��m�(cZ������Ӱ��Y+��z?ɍ�7d���&dg��}�u<~��	މ����K�d�$��R0mA)���	�I'��}�W��J��/�o���:4�f繝R<Cq��:AjI�B��^            ���w�Q\o��oHB������]�\K�ҖiK�O�8(��N^�	\B<�{��
dg}�@��\!{Μ�����<��b��������M�t���`���N����R�'"OgO4*�HM�D�D�v�m�"?�x�ШP�F�":6��������ƑI�K�{fW�%�RYJ�Ч���f8v��M��/h��A1B�#�!"""""""""""""""""""""""��b��������I~��F����՗ݰ@C��0_�$'������USR���K<	����O�m�j�ӥN�~�B�,��z/���̷���`P�A&�'�}���������������������������CDDDDDDD�(�R�!w��F����Ֆ�"E
�5?��)S�%	����?�~y;N�9���N���K�����_��l�ِ'm�)���UՔ�5�U�������C�,�1x�`����Z�~�#_�| """""""""""""""""""""""�1(��������(d��
G{G��Z+(���s��A��-�¢�p5�*��?AdL$��=���<�=Ք�-#�\��;|�0f������γ;F��2A��Դ��6L�7A��P-��D��7]^����*��x��h3��>�5��66L������������������������(9`PQ"H�����)��4�-F.�\H
�?h?v_ٍAp��%�
�ep���U�I�,�а@C��Vv)�𾋍�ŲS�0�<^?h�q_�|��wO�釭?��O�>�T���AD�T�UGE��[�`KI8г�g*�����>!"""�j2
_T�Bg[��}0��ti���?ޭ�m�ɥh;�-�������������������6CDDDDDDD�|\}��'��a�)R೪�adÑHe�
�$���j,:�;/�DTl��c����-��;����ӢI�&����(���G������q��q�/��ͣj�eV�~����JV������7ǘ�cT(�%$�H�"&�c���������$�4�wn�T�d���'<�=�d�>���4�)�>��s�����k�{��J�&P(}!�P�}��5�������q'䎺�y58,DDDDDDDDDDDD���\���쥾�x������b�����������^<2{�\�aN�9hX�!l�䝓�gV�Z���p��-����j���>��9>*�*vK�xPb��oqȊ��hq��a�w,~��z��
M%�B���B�<��eq<}h�:1(�(�8�9 �guR���R�H��KR�,!_AO�&�����}u���I��S��G�����E�oDD����ʧ(������~&$<!�Nb"! �لtsvpFUߪ������)�Y\\��_�Uv�R��2��z���t���[�/h�o����ᛇ���R�u�/u��T��k�,�P:Ki�z�j���?v��`�U%g���CB���<HKDDDDDDDDDD�����;y5�j����
�Whd(��9��w`��E���������:CDDDDDDD�����3�p�A���f&2�e��칲���?l��-A�P\?���F��0��xU(�T�ym�Q����A��Y���OƟ-�D圕�G^O'??	��~��Ӭ1̹:}�4�H3,:Dd<)4����*z.��rx��~"�&A��p��q칺G����?��g��*$�V.>���W��B�헶#*6
DDD�Y7o]����Y�ܡ�=%`"�e�3��e�bmЬP3T�UM�Ř������R���M=0���N�+d�Tc��E�\�M�O�E%(G������o;CDL���;Jf)�:F~���eTX���2(�@��]�7����A1DDDDDDDDDD�X�zd�/~A��m�_��誂�e�����x~#���5N�9"""""��b���������wjo��Eǚ#oc��E�ҝa+r��/����C@P ʎ/���>��h8�;!)�qh��ȘH$'�D�)��e�/�C��
A����lèݣ����n�����_��tX�b���h��]�W��22i^	�ɝ6��Zk�n;s���3s��Ž��@֑/]>5�*�K=��&a��xUXNDDd+rl ���q%��
����_f����3���g�������ː�K��%�!#6��Ā�	�*R�H�����5���K������R�Zmu��,GBKg-�:&O�<F����l�ФP�7]^|/�%�źB"B�E��<�����γ;F�+���$����	�����?�m?%��Y�A1DDDDDDDD��ؠ�����lY�%&���i2��J��o�c��ETl�|I<y�d���R��vR0f�^?8��M�_w����bA�����1䄁�j|�f����Ҟ&]���"T'��D����ʩޗ��t�j�s���k�_�}��U!��=Y�����U쇁�b��� ""��\޹0���*4F��\?��`V�Y�+� ˒���$�z���o���?���\\���R4*�Ȫ�J�`�� �-�ê3��:v�l��~���������������X�b�<��@���%@�g������7`��a8��ޱe�ojc�:�Ō$���O�=�)�G�CDDDDDDD���1&\CBR���E���SwO�ゎ8s����wN����X�X]q$1I�|i���}�'�ǒNKT�9�ˇ=��`R�$u�_D�08Ot�yA1ƾW��'{'�5\��
����..?������i�Sf�"E
x8y���GgvϬ�	2�^�;~��;F�����z2�eĲ��0�>_�y�#"�O���1��5�T��.�]�/S>���u��U�a� ǁ���Bݼum2����gǖs[���Z���Cb������������D���uF� cI�f���~���0���.?��_���Զx[�E�����H��<΃���M��3�'�����CDDDDDDD�R�~��&����n��=T������EpdL$�����bN,�[��EZ&�:�92��y%$"�f5�c0��@�Ɛ����I�&�i8�X�7����#]`%Ge��łT��.�����S˱���_�GpX��1=�=Q9ge��S����#�1���P����ӡ�@�5�� 8�;� ""J�9rR�IputU�pߣ��$�nNn*d�������f,��=7�ꤪFl�jZ�iF���}�~y�
~���2�gB���Q)G%��-�:Y�i)*L���Z�����������(鐿����/t)���1��,9�,�c���Ƿ��Bdr!#[�V�^?���#�r�r�g�i�/n��@DDDDĠ"""""""�D��θ���>������H0@�
}Ք:Uj[��
�齼7�>�7����(����;�WWIH�e��X�/!D���������/
��;.���1t�Pl��Mg���qf�Ϡ����$�I޳��#3z�hl��UoИ.O`ݹuj�b����&>���o������~�C���}��D}h�=���7��WN��p�@��UQ���T�SwOa��� ""����ta�Q}�󡧋'
�P�!c���W\�����<�9�����6�}u���_��ޫ{p- 7��DL\L�~�޾��[�KwF�\��[2sILn9]���.r·���o��R��KN,�������=����qvpƒNKPz\i��$��?��{[x��!�����������^���/�ļ���߫s��!�>�n;���F�Mj6�߀�!�ADDDDD�cPQ"�+�C�����c����t�D圕Q*K)�W�����bN�ڏ���I�]V�����b�,�a�C���R�꼯����
q�d�E�H����[�3p'&�O����_U��U�Ro�TƽW�>tv)�0��4�(�#^���3h� �q�*˒m�����T<Sq�m6��"h	��ۊf*���z�,������Ҟ&�#�?	}kY�%z���Q�H��s�q�����6�ژ4��
g(���~��+|�t������{g���}�����{�?v��
���vΑ9j�P8cH�L���F�l�0���XD�<*���b�C�q���f��������o��a����@�>��`ՙUX�D3�._�|����#!]	����d��%�/�[pl�X������������l�v��Rc��Ɠ���<��Q�r���n��#�>
TA�O��"�\����k�9�r!����K{�������Ǡ"""""""�&Wo�����%�C��"W�1�.?�����Hp��O#�G6�/ﳵ��xߍ�3/����&�-�f�j
Ʈ�]��$�F�����_�U%gN�NX�-
�x��Q/T����Չ7�p��	ԜZKv���U��+��t���7��o���pP|򼜻NM������_���)������F�ar(�+��9u���d�#W�Te�ޫ=�;���?'���˗/���jL�?;.��8J��ʎ/�)MA�2]����a���j����ѯo��K�Wӿ��j���f4����nWǟ��<�K�؂�
�9z�(��:�'�O^���Rއ�"""""""""""[���l����̑�3�:?E.l�Y��4�`��q�;�B��TྜoҽlwuQ"-~�����o>��������
�b���������Ȇ#�~��J�5��|/Cb^���>Z�����]J;�-G�/W	�P��3�d��տ��xѪh+��iV���V�ޫ{A�ɉ=�;-V(��`  ��IDAT�7Iq�l�lU��&)f���|\��NKP&k��mM5��NK�bN��ŀ�������U�󪮫�������C���#YB��>_�9��<���#e���};���|��?DrL����?>y��ƍ��PW�tvpF��m5���\�rT¾k�,Z^.�\�\��f�<��7)$�9����_`R�I:��n	�밠,u��5�y�u0�Lo���6�N"_�|��E�����9u�F��iU(��h�R����}&�L:�뺸+��\�w�ѱ��;�����u^�y�<9��k��s$������8�!"""""""J@r���E[#)�b�Sj �Q �w�o�8�q���6_��?>4J�'m4/�I���@���Ua'Qr"W}��zz���]���|Ns<�x���#żU'U�B����Q�4.�3��D�%��>5��s�U����4�8�;�m��C3ADDd��/R'�Jp�9	W��������'9	����6?�e�,��YK� -�K��8(F>��E�n0�>4{�)��Р����loS�������f/C����������������#a.��9��7Ǻ��T@̻�d,�a5��]�v���7U�YW��ěGƩ7����u�w
�'W�ƞ�غ�.֚A1DDDDD&`PQ�B�QMF��b5)x�M�j�A�ļ2b�Ud��H�\s�α�(.���F��~���_]�>�(��,:����(9\m0�����mkϮE�ymi�X)S�����]���ԩR#:.����Q�Bn5������֘�z�[�&' �����d����ѯb?��ɯ٧n޺�!""�� ��~(���f��!��84��ː�!�`y��}j�e�2��s�Κ�������!�C7��w�l��m�*��6%���Q3wM���7���V:b^9}�4:,��C��a�S�Wf����|�ݖ����\��vz�i�qL��x���q���� """""�CDDDDDDD� rz�T_�V�Q	I���t\��fWVO,a�a�rݗX�u�UǍ����v�*	j;�-�}v���H*f���^9���_�]��K�_޺mg�N�Cb$�Z�jhR���SьE�h��_c.=���k��������:��{�ײ^pwrG�"-_��s���?h?�������p¾	��r�f�r�ˁ��Ț�����"�E�}Je)'{'�'���gV�a�C�sM��=oڼ*�E>w�C�|d~-c��QA/��se��<��YK�l�P�����zMQ�$�]�wNࣹ}��'��5&4�����7&U�g4,q��u��=
?��!^�\|Oέ\uf������0��X�R��g�?Օ6����b��5��>�Z}�-W��%'� �q>d�]Ơ5�0��L$v���Ϩ��.:-�Oo��C%ſ;.T��W�JN�g77x"�v����+�W!eƒ|Jf.��������쟂헷��/A'2���n���o��\]jA�(�GA<C�m��Mo{V��6/�wvpF~��j��I]�K&y=H�ZXT�?������R'~%..(��(
�P'��9�!�S�xI�QL\�E<SW��d�o<���ޒ�
��L_�2�5տ'���d}��?��7'鐆l�P<sq�x�x��(y|�G<ǵ�������cI*�MN�,��0�˫��^.^걗m��n������gq��$�`:��J X>�|ȝ6��ox:{�� �٫��b��������{fG��E�'m�O�^-[B)�=FГ �~\ %]�ϯGtl�[�oJe�
�3V!!d:�v�1T�2]u��Iι�s��9�o��&ۀ�V�Z���#��
�+  ( DDDDDDDDDDD����]�{�~+������ѽlw�������u���Qg�Π�b��1(������H�!"""""""��2sr���]�7��M6aԞQ�Pɗ��o�����ژs��Ar0��,4*�-
�@RRշ*N|qBf콺D�o�|�
�_�Е6�ڨ�_}$HiF��p�R���hY�%<�=t�	�h;�-�~\��Y�	=_��
�_�@� a�H!y�,����z��z���[�sVF�H�"����c�ŭXyz%֞]���+���S�{-��P�׺:�Y�㷏� ��A��1��!��ɺ�"�e'�Ż]�4z��%;�L�2w	��rq��&9�Il�ӯb?�.��22��I��>�Z�T�X��(�2m��A�**�4$���㋰��:>dMsTD��]t��ܩ�	�%ۄz��{����>�S����$`fR�I:���z���~��MB->��1�j�b������������7���+�
�[kR�	l���v�m���G$7r\q���:Ԓ�3����.}Q��m����NGrv��E��޿Z$ܧF����oDxt8�e����|����"�$�%<���.�Ё�LO`&L���������p��M�q�rT��&�!"""""�0(�������������o�j���A�t_�=I���skq%��*p���'ױ��n$}��U���2ڊRl�tTaD)����ۅ����\МG�w��3���Y�k+�]�x��X���m��¬C�I���C͠���f�2�d,�v�۩���is[4���7ڗh��{����]��PS�Ff��K`\�q*(���R�\�rjPy�Z�m��a��1&�U��iZA���fP��'�V苟���?c�8����$�f��*|!1Hp�7��Q�r�k,�_w+�MM���n0�=���������O�>*,�T2O�b��t5��
�����v�,aGZ�!	�z7(�f��|<
g(l�2t�$�Hk��nPLF���d�چ*�f?y�h-Og"(����.?l�ɕ����dH�A�����zn��\��b�?���]��(��<\]5����Ú�~�1h��t�KhՈ-#@DDDDDDDDDDD	G����}a���\�ά��VSu~/("���z��uLgP�|�KDDDDD�aP��IQ��t~����\�Sy褠wΑ9�@�R��/B��8$&$�c��ER�d�������z`*�>CkU'�����>�>2[���j3K1�#�-�/m�ᛇ���#5	w'wU^(C!�!��ԩR���hг\O��S[�.�?��0t]��ߓ�'z۝�,����&K�B^7c��QAt���ǭ:�����7���v)�`m2~ろUp���*$hmy�娕��E�H�Á����1jϨ���뺯S�K�,�R=���z+H��d�(�ɑG�crk���ŜvsнlwtZ�	7��@B������}25,,�����f����˕c����\�깪�p�K/�V*d��#WE�ux��Ga�����r����5,*̬q+���7��k���� ͠�RYJ��epEDDDDDDDDDDD	#m괚��o6{\9�D.�&|x��{��z���;'u���l�w�DDDDD��b���������(�cl�ML%eRԿ��:$�?��A�OL���V$7��OB��P0}A��'E�rR�����#�EωL�h�c��� z��{�cɎ��0�����0}!1�.l��[�7�d gg�Юx;�.���u�fN}q��{�C��n�w���:H��������-?�O~ؚ,c���h?�=V�Ym�1]]���FT�Y�+���ξ;-XyEC~o�;r�͍~+�����IȐ�J(�5H���%j[7f�X���f���Bil��oUt-�T!^�������V�N�:f͟2���X�4��x����\����.��]3^?	��U��\�%lEv�l��7��Dr���.�����������Z2sIͶg��I��&A1���$����# """"""""""��!�'j������������>��~���L��QrƠ""""""""+Ie�
+���($&�qn?�_/_dt�[���u����xz����r��f���Hn����cs���5��l�8��������VSQ=Wu�Ɲ�|�>��S�A�>�^��ڗ����z��sB���U��t�E�D����Xt|�I����֫I��%�r�К�kТp���(�#�� iK�:�����O�>p�w²���lv3l<�Ѣ�$<B�D��	\Z�m��Bb�$�#a1�$ǡzn�ZH�+���n2Z_L�7�j��U��َb����ҹ�S�Dg6�ޫ{m�	h��q��!1"���3G��mձ�<W�X��Suň.������ 2&����6��h�O;0ə����v��C�+���f�����+���f۱��l"v��!��N�!""""""""""J8Z���=,=��:o��zk���Q��v������?�!"""""""�)��~.j�m��R(6`� �;�N�.��-��ĴV�����V�-$7�.m�((&�Z�M�X�[.n���Q>{y���?�����.>���Sk�[�n�t���إ�������#쾲D�%:�������+A�ZL�Y�/�ݵ��Ɓ�,Z9hɉ%F��{��ѡd|��;�|�_V��*tB��s�}U�7=�|��wN�0�k��!$<!!��1WGWu�.		)���e/�,�Y�g���:.B��%p5�����q��U�!��î�]����>����^D�P�9y���S���P�3FьE��c�����g��{
�oP�-�1y��q��Y=��
5������?��1.=����� �ٯf���M��A�� �In>����(,#�i9�jT���F�#���G��ta���+� ;��D��E��������>�{~�/��ދ�<Hx�L��?u��*�܄r�y��a����=}��Ї8{���F�������z��z��>���T�}�cN�9�!1�X�}\-�዇j;%W,,�S E3Uag�.w���굮+Sw���O,����􃋃��6	��|�������'�O@��G�<�4�%T%&.��q%�/�WN�vٗ�����ն_k��7]^�69.)���
2��O���5"�#ن�zzKm�N�=�;������������~N9�RZc�F����J��{DDDDD�b���������`dÑhW����I��Ā��q�*n~���V�ʣ+���*H�	��w,��헷�z?�=��&g#w�TE�搢�����M^��{���"�E�H����X�m5�O(����7%2�x��V����߻|o��ʡ��ߊ~�ĘC�y%�
ry�R���RYJ��ͣ��j殩�]���`-�����?Xyz%֜]����#��5r�@���T��V��~Mo5����'�����N�}���<�O2u[/���WD�BMмps�I��P%g��ױ�����/��M��lѷb_|W�;�j�5�{����I�2�Q6[�x�K������;�9�x��*�pH�!Te�
6�E�	$):��E�H�����!1�oƯ;��sk����]�����Vs�
��En_�e%J�+e� ����O�>�n������S���Ru�^��_����j�ɚ�2��,8�;�k�zi+�����j��)'�6)�$^ Ltl4f��o�|�s>ٟ�"(F��"��u��_�������<m�����]L�!a\��i��s&�%aT���I�*嬄u�ס�o���$TK��$@x���V=$"""""""""��\�A�7�=4��Z�M����%G�!"""""""�P���e�/M��a�Ct[��o��s��	��2����5���7���/��V��67tG
�3)V��C�غ|��U$���KT��&6��>��R�'����I�\���}���!�ѿR�m�Ϭ�ܣs�d}��X�ᵆ��M��bt��}���	u�v`��SƙC�۝�;�� �h=��3��[+O-��_�/l6y9-
��,D��H��U��9$������l�:y�`P�Ax	��r�U:k�x�M
����~fp_(� ̞1X{v�*0��_g?9�OB=J�+m�������_�_B`��e֜Y�B�ҦN���<�㚍C����^W����[W�]��>^�
2�<3��l�W!��@�B
���ߪ�k��'~В\=�_38���n�w0���'*���m7��@����q�!��Yx|�ζ�f`X�a*��]�����K/�Z�9�:f���Q!�ə3��Ϲ��@�� ���k���T�}bH�z�o>�	[����VparW.[9�瑠-	���A��5z�h<
"""""""""""C��P��1���9��b��������,��=涟���M�ϭ�lv3��m������j�Uѐ%��Գ�Fr%E�R�(���H�Œr2���l3Ӥ��XY���!�}W�U����cT����f,����,7/l�(�T�����[/m��[:Ki�N�[g��%��w�#�k��Q��}T��xa�l����y���'�O`-�.lR�^{?ًl�t�Zc�YA14�l��sCb�%�4y�����[�@���|R^�@ԛ^����)�����Y�g������!1o���ƳcG��A}m��UǺ�#�P_��Z�]B�Ϩo�1��:֚Z+��PI�|Q���r�2��Lu\��Wջ�貺����1�x�y�����sT�r=U����*�K�M�Ø�`�/�}���j�URA��Q���6i�}�l�͑>Mz���d+2�� 4�!M��I0�7��Q���6S�[�8������������������>�!"""""""2�}J{,�[oo��[~j9�,ꂰ�0��G�Fa��i������\�:"&�ٙ{g������n�ɥ�|�f��.R�oja�}p��],� v��&z��;����/Jf)���/�^���#�}��4$�����HL�|�o��K�~/��$�mh�W��������ͣ/k�Α���O��������c�v	���Ua��*���ğ��=3�'I�����R��pfC����t��`�9G� 6.�0e���8��:bu��:�%$D
���Ģ�o�~{��y׳�g*��Ҡ���p����>;�^����_a�ꁰ������	 ��&WS?�Eutň����Mߨ���ܝ�Ѷx[����#9���"Zi����A���	#j�w�}��������Ko��[ي���YF�i���Y�f踰#��?�b���������$E�UrV1i�
t��}MΐpK�b��u��YH���;k�|�|={���y�s�ҹtg��Y~�Y�Zvr"�#���r�"p}�����?�<���N���gy��l��c�5���VN��w!�I�F�@L_P�.E�..6�x�|T�#�}rsr���u_ �������ÐC�I�G��-TH�)2�ɠ��c���}��D/��쇘���9u�F���k��]�K�x|�镰�{��a�ơ�����~Z����S�SB]*d���%z.�;k�Q�����W��w�q��C�������$xH�迪�UCbĶK�p%�
ry�ז�5Zia��?�R~j��K�� l���UV��X�eR�H���M'��6��H�%�~�Yl
��&Ǳ$*�nd;�ϓ�P��p��MQ�Ơ""""""""3��ʉojc�<�����U�)�Rؘ�+̱��*^y���
�e�|R ��ktP���q��e�;��u���������F���A�������k���z��)��v�k�H
���P	�8s��+;4���T�u��1�桙�se����×տԹ�����IA12F��iu�=z��	�p��%��5r�Ht)��@�7�~�A1�7ǳ�gVk����]�%ۉN�:a��aF��qŏ5��]ۧ�I��^ڪBm�%�M5�����L	�z�	m��6y=I���S�G�?t��.��*%2����g��������-��z���#�=D���ޏ����f��Ǿ��E�H�Fo���ڊ��e���|&�}��=�Y�38�9��OO�Q�/�}w�ꤪ*̍�����������������/��ab��pvp6�����ʁ����}x6~l�|�������^U����a����f��`����O0y�v��a֡Y�~y;��2o�~���f_��v��;,���kH
���
�x��XCj1�OOܝ�������K���e����d�'x_H���
��V.^[�leMK���Z^�����D��x��VO�����t���>ܜܬ�"$�`���VO�O�N�B����kctP���VE[i��ٴ0GcI𑮠� ��<}�姖#1L
�d���3�O�ҹM�����c0,M���˫m�.ѱ����_Hnd?�y��ѥtا4|j����s�6�~�5\�]��uqW�}vע�H�>1�CA1��|�$q�ŭ������8�<�b�t��m^�Q-W5�.����Ǘy�wY�Sj��%O�!"""""""2Q��-Ш@#��o��=���($F�qX��V)�����C��"~	^�W��J�@�,s⾉(��z��a����FCdL$���ԩR��{hd�޾Z��I%���������d-�&[Yqj�,�YL�T�}\gP���2�g���F�%��Ln���.���w���������$K-<�?��)R����h�*9�`��V[޲�ˬ^����B�cY_o_5]�jp	k�
l����
���=W�� <�xm5rװ�$d21 �u���V��/��'��s�����ݫ|/|��+���]��fۺs�,�H,�z�����~NN�t�T��B
�r����_�vC�Y�gaW�.��$nv��z�q�㬲}6�b(���b�wP̩��0���9�F퇌%�X2�=:�������6��WC+娄��|g�`4""""""""""""""""J�CDDDDDDDd)��l����_A���R�)c�c����{B"B̚���ۓ�M6cJ��!�W�G�L�Q*K)��˗.V�?v�����Ё��0;N�N�m�n�M�����M~~��&L�8T.1<}�����kRP̥��t�H8ҴV��bNX��-9���c�q���GP6[Y���rU�jP�ғKam��$��
�Х�oU��b�o�ٶ��J���$�)�Z ���-�GVU����#�,k���H�/lFl\�M�1��T�A1�k��f�7ff�;��m���L��J����l��2^?����x�_�m���W����nj��i�c��9CcZ��ћGQ~By�q�ⱞ�?U�Y[�y�f�z�Y�K�����؉�������������������y�������ٍ���sZ��Xk�rˬ�$ԃ��2EJ��sHɠ�7�è~������B?����M����_b���x�DIQdl�[���O��W_�*�F�"�I�ڛlY��>���������&Z�X��$t���fdL�f[F��&-sg�NT�U]g[ろ����[�^DRv �mƽ~@3(F�ԬE�B�8k����
Z�އr��i�����?����2+{,^���}�AB-lM^�'���|�sM�EZ`�	�Ö�J�ivH ����A��ڏ�3��m2���v�ݡ�b��}vm�1+�HCAir�h��P߱�xB�l���cV�γ;�3�����^�zi�Ke�
#�P������������������(�aP���0���W�q8N�=e��#EiƆz$�^�<u�Ԡ�\r�^<B��i���fP�������5�4c�|RtܷB_��3DIѻ!F��\����)R�k�r��Hl�hT��$5!!�w��n�rS�z��d�(��
g(����p��9�Ye�4Ų���}��5jj殉�_�U!xs��U�8I-dG�P$L�$\C�<��r��e�E���>h�s$$_�|���-���fq�b�e�mDbH��1e�Lk5Mg[���
���0��Ľ��M�'&ퟄ�������g��}�#O�<�}�ÂQgzRd-��$L�Y�3؂��N�Z�l�$/C�hR��f����b��aV��MDDDDDDDDDDDDDDDDI�b���������ԩT'���aT�=W�`��x�._�9�
�N�NF�#Ş�#���enP�̻:�"4�a��}\���s��o���b���4���1y�d�G��(�		; �[;R$,A�Ӥ�ז�-�
TJl>�>o��X�I��Ll1}*�A���p���Yn6�l�Q��*,��a-�
��%�ߥ'��]�v�}�Rڡq��j����ᛇ���Vl��GnQA-�����6�9y�f��;�;Z%�A�rl9vv��痀#y�Ck��T�����}��r�!�H`BXx|!~o�����F�*�C��U.[9�cCy?�>2��}��aȆ!��d<	@��{�
W�"a-�gԷ�����͔���`PL,�b�-&.~�py��x�֯��7�k�@T""""""""""R<�=0���ƨ�����Ke)e��o��[������2�!"""""""2���9̨�R��ɪO�~�z���������y��:���bTcevˌ�/��eLP�-B�$������o/R�Ha�|R�ݫ\/4C��\{|���ͫ�`p�Π����cW�.$��is������H`��	�pstC&�LFl�P������{u/lEN����O*h���4s�S��ٚ���gYܳ�+�w����]��T���`�����Q/���ܱ��r�E�����F�ǝg�s�90�������X$P�$d"�$Բ%|q�?�пR�xm�Z�Y��
11V��5�֜Y�����ݏ�8�s�����A��ϒ�{m�X�Ƴ��ͣV_���V������؉���������g�?5�4/ܜA1DDDDDDDDDD�H����~��د��'""""���A1DDDDDDDDFh��A��w-��O����_��JSH�4�'�{f��eP�.=�d���&�¾k����4.�ؤ��WU�QR�����5���`���P^�z��T�Q)��U}�b�ΑHLܑ7�A7����C����\�Ө�ƒ�'�嫇Υ:�-*���u�סƔ8v��o-
���63�Ia	͔@�W�=��泛ccύ�q�1i^)d����jfѱ�8t���\��'�A��ڳH��*��t��JP�-���-A+��������#a8I��Bd���q���H��M=0UgP��Z�+���-�b��#�ж��j�O?8�;	 5�u!a"Oß���S�����p������zn@��e4���圖��o�u0t<eN8����o�ݐ��ن�P�x�x�l/����}'}xCDDDDDDDd�ne��O�\~�����C
�Mq��q�2�e2{��`g�Nпn?�m����WS|��;4*�Ȥ�<i�p	�!JjN�;���k��K`L~��8��ξ;.���*���^3OMju;����V�g*�4�i^�~��i$G�%��2��;틷��5�Zܜܰ��R�[Ҫ!+��fc�2EJ�O$���RX�i	*�h�8v��cF7���7��4	[�	i�)Ɨ �Tv�t�[+�Ė��P���+v��}�k��^D�@bH����q�ս*��]ռps,=���8KvT!C�>
Ď�x�I�K�ƅ����vgm��:C�^��~����������S��L�*�P��� ۑ��[/nE��u��~�P�B6	$"""""""""""""""���A1DDDDDDDDH�U����;1`"�>�ٺDǙ�q%�
�?Y=��=o��%@�1&�A1R���v��[Ǥ����ΠJ��X�UP���k�l��!!pwr�v	����g�n0K��5��]�Wr���K,<�Pm�6�ڌ��u����[N��B?�,�m��l�Q�Z���]GWTح��T`MXtb�b��{4��]�t���
��ʓ*�M�6���O*���)�ѴPS4)��έC�U�q��MX[XTlI�O�;(&����M^F�����}��������\�;e��A1�w��F�H?-3�P�7"s9�;be���o��2ݗt���+m�.����۞�3�͖�u�"��ٖi�_o_�%��O��ʕ+���������	�۳������{""""""""�J�����`�ȘH��o�u1%xC
��G>��p��f�[2sI��>�k��-�bĄ}L�i]�5����P%%���+��&��+��Y�f��j��k��������8u�C������A1�����l����Mg��%;�b�y�̳hY�6��4�!1Q�QXrb�
b��������n�a+� ���2T�U]JwA����$�B	����":-��6Ú\R����/��,��v������]��!����G�4��I`Z�(Ps�r�ʡX�b:�d7���K������__����,�c�~�A����[�jH6��k��@�e( 8�{Q�x���lق�g��l�s�ҤI�:8F�W������ ""2�b���������Z��Q���Z
mɔ���!�Ao+������P������!�e�M�a������2�e2zWGWd��aJj����A������+�_o_\������cЧB�N����%�ay��(3�B"B�����lֲ�ƞ�{@�9w��,�U]Wi��l,֟[�'�O�^��~��"��Z���߃�R;���I8����j�Oi�RYJ��j�����4�iL3m�X�m-�j�m��Ym]��`+N�NHe�J�=":�*��
2���C���%�I����4�)�4�2��,�5<^��(ի\/�0Ds���{k��:�J�W��a���;�G�B�4�HH�'�>��C3d�n��BL\���/��rl)�L-�3(��m��3.%���`̝;W��h�]����x����*4���G����x$#��w�0""J�CDDDDDDD�G�(���Q}�:�lM
��u?Զ�5���_0�C
��窎M6���y7����� E��T�Ĥ��l Jr�=%�c�+�W����W��W���_��~��������̓��h>�9Z�^��4��~`�o}1���2�Β��gVc��hW���voo����/�_�3��~��R��gy��)��t�DB��ʡ��4r�HU�_4cQT�YU|����Ӥ7j,;,��F��'׭�~�����]o���VY�-���P��� �i2h�kQ�5��t�1D���յLW|��[��y-�-�Vs�i���)S��춳ѦX����)�� ��1����q�.9�r�d��7}'^|xd[���$H��������������VTT�͛�7$�111x���egg��b$4F�c^ȼ�)!3DD�|q/@DDDDDDD�Gݼu��'E����ak�oD�D��S.[9�Ǩ��>�b�?c�b\S����+N�09(�V�Z�Oio�} JH8�*(F�(����w������ݿ�n��*��]�2��O㇭?`���3z=�@Z�'T#A���68������{H�OW�������Cg{���1i�$=2y�VE[��M�ˏ.�e[+$Fx�x!1�������j��o�z���ZM5E�R���#���ݝ��}���mI7�����Jf7���C��߳�r��g��d�����0��ӛ�m�~��'�O@�	i�xa�
�{��[�n����ձdG��F�^��+�Ad*ه�l3S�?��07��$�c��iŔ�RR.�~њ}���/ٖ���+1 """""""""��c��-H18��(qm߾O�>�-���"88XM��I��uh̛22�Nm�=Q�cP��Ŭ9���Y��:�!W����W��1�o�O��v)��I������^<}�t�錞GB��1 ( DI���	=��WN�N���o輨�����i5��~����.�	㚍��Zñ��B켼S���=~�_�)��+'�e,��yj�"!�[Fն3p�Q��c�������m�����# �$`�]�adÑ:�����/踠��c��]C���}�d_/_$%�s��!5��2�7W�\޹4�@��7}�;��X���>��h�h���b��i�I�JTl�U�S4SQ؊lg�H`�!�_�۞�'^?z�L=0UgP��]��Π�]���Ux�)�xhj���VFp��/F��� Ǌm����&���f,j���J9+i�����;�-	��'42DDDDDDDDDDDDD�p^�x�cǎ%�j����j�~=�97���*H�U�������������2eJ���A1DDDDDDDD�j�R0o��V !��Ǡ�7��_��1���3f1���t�4�'���b$(c��Q��I���W�A1�$��������J�a�����Kg��`ԜZ뺯C��et����AU�IH�����$<I�-�%��U��[����g�~�'`@���Ig{����Ǯ?p��	�ƕ"q-+O��59�9�L�2H�d!�h��o���kQ+O-��䘯N�:�{t��˔Ǥ�O��7c���ػ����?2!H @(A� �	((ME�HQDDEŵ��E]�u˪k��� XTT�4�]�PB-��>����>a�̄��0I���dfν�N�{�^r���vn����4���?y:T��+�&?�W�ےf�W�󓠘����� Z�WW5��=�>���k�ԻD�"\��ce�	�?d����<�{a�zy��:_�����\�����b�\�`4��q��y�L8(          �g�����ʒ/3�/..Ζ������*W�l�cr�d�|  ��#(     �3�=,��a�i�Z�k��CA�b��>G�Z-U�J=��u{���ďO���Z��9�)��Z+��(xP�E�5v�X�f鞥��q�nlw�}n.9�K��O{���Ѥ���~�>�u���v���Pw�$e�f&��,�r��adƦZ�Dț	�0�@��������!_)P��6p�zZV����(����z������սQw��K\��2��t���m�'�g�s.��ۀ��2צ�vt[��P����VkP�A.��7�o�P�d����+?�+�_�Ug>M�S��:��ݝ�v��w[�S�������5T^L@�?��S�Ӫ��������Y�u����=��Z!��4������s�;3D��         ����S���9�N�����Jpp���S�T�r:L�<>W�D @� (     ��f�Lg��CA�7��QVk;�cm�r�-v�jV�o��m�*T;�2�����ӾN{������#|�c?<�~��)4(�>�[��c�v�rf;]���������n��W�yU�v+���M�=� ���~t� b3xټ��g�?�SW>eǮ�0�y��І|���6(�
y�mnPIa�#�Z��Fw�vhm�m�=��������ym�x�b�n�ƶ7z<(�o��y�0.�������_�Ř ��U2h���z�����6��n�x����ye83�qx��n�1�3@A�y�z��Cy.��oo���C�����l�r��z�e�L@�'m34�~s"��U�Qކ������?��!          ��СC*�RSSm����UW�|ysfx�)9�9 �A1      n���2_˭?�^���t5pҝ�y�f`��#=�^͐��߼�~���ʲ&՛�sO���֣[���f��KV�P��#����h�����2b���Lp̄!t�w����{W�	�mX�X?�� ����m�߯;h�����ϟ��Sw^���F�q�k&��PB��I�����W5�	.��9ll����|��W��m]A�!��D�ۥSI���j�u��=�������<��_��3�s�=��IC��虣=�xS�����٥��{��ά���1�j7�=��Y�9�N�d9�|L�n�V7_|s�:s�=�� }��[_1���6�ۮ%QK�	�{�G�w�.{WO���|���vS)���os�&���m���v�u���i����w����<C�Mhj^��          <�ԩSJI���%Qff��=j�+�����cL�Q���W�n�d����� pn�      �Ѫv�|-g����nT�X]�z^�S�6�h���x��Ŵ����\P�3�}��-�T�S��kY�%A1�Y_��J�v�=]�9��y���~���=���R�J=u����,�S��BC�2��I�H�����q|�`o�b��n��0�3}��SMZ;I(��V���z��g��uq����й��R2Sl1!.e�LX������.���Ԅbَ	+y���z��'<Ҟ	Ÿ���n�g�9[I�I�$8xk�[5q�D��רZ#i5�m�	>ȯÉ���m�+#;��+_��3(Y>\�ˠ�&(&�c���Y@~���1W��s�~�@��zD�d�����lCa\y�����~J�����׏�kU�7�TY�_�|�˘�4          �'==�{�yHMM�%:::W�	�1�19!2�q��;�  ��     p�e͖�Z���b��)��f�vx�pO>��lT�Qo�{���ڰ���Y��ʄ��Kq�[�l-TP��[�����f5�ف�9���)��j�G+�Tv��1�/��ɏ���k���=K�{B����W���Cƻ�77����A��W{�_?�~�������kގy**��R��T�DT�p[w��g��Fw��V|��1;����W>mC�ܙ��;M�������y}��6���yfʺ)j��1���S����J�JJsmm��Z�n����W��7�]D;�����k��������2An�����g�̾�����o_�����i�z���k^s[����OV}"x�9�M�yj���l�fl�!          ��!1�fd:d�_9������R���@��ի+  @ ��     ��	��\��e:3���.��<t�y��e:(����ݍ^i����Q�O��,2�]>G^��=�h�����0(�|1��M8�o��v����/�ߞ�n��6ŧ����PQ\��n�p�Y��A�'$��>]��r�um�k��n~��"�G��1���"Ŕw��ÿPH`�<�B�
v�7]���uێn���p�{�`�V�Z��x���֛ ����I�P+��^��r�C���{]������6��1�|-ܵPW6��e���.�GC?����V�nY����W����S|��[Ŧ�
8�����g��LZ;Iws��v�{s񛺷˽r�9\�_���\�c��
����?h?Gݙ�q����UYuI�K����|�6����sX��y���-ߕ��        �Ad�H��@�ԬPS��� �&N�Sqqq�DEE�>c�	�1�29��,"(     ���U�k��'���n���BK����z��v@�7�m�W��w��}+Uִ��Z5*�8�r���0� Tm ��%�%��'}5��jS���������׈�F��Pۈ��z�T{^9�G�P�O�k`Mi������������$�A��N���m͍����vY7��P]��*;x�0��뛑ߨ[�n�43������ͦo���J�F�տ���v�g���/�Z�Pw}sW���U��_��EA�An�7���&,�B7��a���2�m����4��B���G��56�Ǖ�G���{��G����ڡ��p���q���ƂgL^7Y�^��0*X��G+?p.�������s�i�iԌQ^�l-�=�{���/t�%w��7�O3n��~��Sjfj���yaO�>�u��ΌBn�&����\���,s�)���SFLQ�{乜	-~qދ        %[��̿��X�� ��IMM�%:::W����BBBT�F����"c��w P     �BX����v��¨[�n��1�s?\�ʢ�!55�Q^k��8�p�uz��O"�3�=?�W�n��e�fva�X�\E@Ip4�z��C?��ᬀj�����x��z��g���m��ڀ��]G����[
��.׵�]��E���TO]���`�k�_��u;j큵y��k�z��7\֙s�w�}�����������חÿ<���h_��$z���zo�{��q�%*r�&���w�9\�N<�y;��� ���=2�;�>���7լQ��][s`���m&0����{k�[
�1�W���}��S�OѪ��
��6ެ�}ކ��3����h�;g��P-�]��rBs�ŷ(�?P1'c�IJOҔuSt�e��{��G�jٞe��h�G����s�o7���Fʙ픯3�~׷����i������'ߘ��+j9Ȇ���6w�]���ۮ��������ž/�����W�w/.t�]�
�tO�{�x��U�B�s.o��&�          ʺ��,����yV���Phh��1�1&8�<6�z��
 �T�      �P9�r��;�|\�%"4�������ʪg{=����^���u.�a4fpYҧi�|-g	Vk�mG��ێ%"(&�������qPuG�;N��W�O�v�׆!�_>^o/}�#禰�0�p��]V�b��������*x�	�zu�zo�{.��g�	��ـ<�1�	?o�Y���wYo�q�>�T//xY�,}��[y1��/Pc��
�+�UgBC�D�Q�f}�I�6Л׾iJL �7����m�u"�@�ԫRO��x�#yz���+ә)O0�'��v��fxqY����OOj���y���������1�+�]��/&��au+��P��]N?7���}�k�O����phC�뛰>zd���L���<��cEz�����.�����v�5[h��v ���ߴ���|v���K�]�������e�.cӀ��s��;s�G��������s���bBȾ���ez^�S�ߤ澠Ik')%3��r&�ĜwL V^3�E���^������{h�����.b�v?��@�����v��Ra�
��.��)'�p�Bm��h�̶ޢ}q�\�g~��j4��c�u��m��u��	>{���       ��0�Pk��Vx���!�f���q��}��d  W�N������}ς��Oǘb�dL�L�����FP     ��f����'�/(�q��^���ixS;��,i]��^��gg�K�SYP�r]���|/ogGPLfv����8|�	65}��D-��!�U1���РP=s�3z��6�c���Z�s��$�w�5*����Ѝ�nT�f�]k��8������|.x�	3�֕k�_c��޿:�v��a���Fu�#���<��	���g-߳\{b�(6%ֆ���m�!���juk��m�Ǆ�'hw�n���0a+�v������s����z;��<7��|5ǃ`]�J];�ڼ����y���,���)�����6!Kgj�Vs�k��f�9�~�N��A=��]'��<1Ǟ9�����н�A%�%�
��դ��?�^k�Ѽ���z�=�d��^X=�ߚ�U尿�>����,���m�9S��j�rFL�_���"�ǅ=l�pf�߻	�1a5f2�|�kSL8L���>d�P�L��	�2
�b΍��M��r�_>:o����P�bu�����/��ڙ!�e�L>���{��m`�G�����=כ�
�z.�X6i��ӓ�)��ʫQ�Fk/�?����|U�*T�mo��L朚��`�9ט���UաМ{���:{.       �|1��M?���&W�Pzw̽as�����`{w!�  �����DGG����WHH��1�1&8&'P�F�� �'>�      \�T9_�9��*���\״�F���VP�ۃ�v;���L���׿���ܤ�����������k4Wq(� ?3H�"�A�@IbB�Zd�3�xV�9�mq�-Ǝ�;���'v+:!Z)�)6TÄ �P�Z��ԸZc�dB�2k�,=<�a:�x��E�E��߭;c��k>�&�v�Z�翨�~>��*VҰ��l)��;������ݯ�b�[Vb�'�߯&ݠLg����2f�u����6욫��5�ѴH��mMX�pWFN���Tês�u��ɖ�x��l،'�����5���j�9�7���w��������+(fƦe&�p��o�a0& ./!�!�b�-eBI���zℂ3p����E���?���>6�       ���ܓ}����9���ץ~[̄6_��J���_ �/���R\\�-QQQ��M�Lxxx��<((H �m�      �`��GyGy�U���1��H�g�TV���W6��X�9��p��6[S�MQif���>Q
;�9�	�AId�Z}>�
~���l�WLǜ�v�qg���zqދ�9G�OV~���|J�.��7�K�]�U�W���?��ӆ�&�\~���0n��Tf����x��YzV��|1D�]�6��x��w����~xL�v,��$��|��bad��������+?�'�s��IC���Okl����v�zk�[
���r�ޗ��&'�%�aY����_���|����q����.%�'	        #�?�N���S�i��^ŀ���OtS��O�f���I�����@��k (ݒ��lq"|:8�$cdr�+WN PT��     p�ԩS�Z��_��%l�mD[��h���Uڙ���_��y���!�l�2�ݫ���6�8p�y��*���qf;�dfЮ)& ���wk`ˁn;DJf�f�1K��H�w/�OZV�^]������eLF�O��َ���e�-:�pH�t{�#7�M���P�zX��Ly�)��ګ����|�������1'c�}Bw�9C�/�]���~��O��^\�ݦ�޻L?��Q�k�.r{'RN莯�Џ�(o0���濤_#�;���e.��E���g�?<�.M\3Qc��v�-������(�LX�u_^�g{=��z=�@[�6l�0m=�U8?L8�#���?f
       �3}p�����.��}�����c�
ӯw��K�]����^�o��a�=^  J���T[���s�9�����c�cre���U�|�M P�     �B~?{j ֹ%(Ƹ��]z��T����\�*T;/ۯTYߎ�V=�'Uژ]̠Âj�T?��Y
����|Y�k�-�3̀�ԳqOuo����y<RK��hѮE��ϟ����}��=u�S6 ͕~���s��Z�oe��ϸ�~x̆��q�j\�q�ߓ$��̇�~��o�^���^�����_��]���S��b���z�gl JqHHKP�O��.��~/��s��`�;H��#�������~^��x��JWP&`h��i��O��E޶��Zu����B�p����m�H�v3y�d-ۻ,��(8�Y�WP��+?���|�8�E}��;�g�ԧi�B���/�����?�pfg{��'l8�	��������=má6n����       ���۴��g�޲�<�-�'k��f{,$�L/�}Q���:a
 �	� ���t*..Ζ�����L_�ʕ+��1A2g>
*x�- �A1      .�e��k�
T��h^��G]2J��Stb�J���>dj�O.��#&k�C�}*[���6Cպv��g:\X�B�8�C�T�r�B����*�4ILK��Sm1*T�� ��6Rx�p�<�`��P���ǵ'v�v��,�!W��_�!G9�7�7�\l��\���6R/��v����|�7k�,���']��z�������IG5w�\}��K�*�e<5�)����2mo��h��^V��*6��z��b~f.Բ��zB3}�t��7�}������n�n�x������:�3�t�3�6��HK�,����y��n���:�yzV�=6�Y����~�6��9�aUL`�����Cn��}�3miV����k�_c��
.g�����&��O|/k�u{ܬ;�N��<�t�]_�&jX��ۺ���PZ|��3-��:�+>-^�&�D��}i����5Y�Yn���`B@��ϣڐ�V�Z���w�ϾF��s=smh���l�FS�M�ǘ�Ŝ�9ￗc��
��9O�b΍�+VW׆]���\����^1�u��k�y�\�m9�E        �ӱnG���n���~���5�-���[����z��r �Wذ�x��o˞={r���1�J�*��d�c4�� (     ��)'�\�*�T�D�)��A�As�=<�a�FW4�B�x]�`H�!z���򥁈EU9�������@o���_�u�ғ�H�43�N7Eo����oo�W�Rx�3۩�f�b�l_�_d8�bfK�HQ\j� 0�w��ps�����i&(���ڒÜ�L�)5+մ�G��++�?оw�d޿	�1�&�W$�'�Y�L	S�:�l�I�J5b�1��q����Vpc�����Rf0���^�%"4�ș�Z�j�XI��L�=�>�[[�lՖ#[ι��/���U[���բf�`��{���1��2!5A������)�x�"�Ez%,� �� �9�ڢ�TR��ҿ����q��*-�gsIr �@�ڗ��iIz��`B����-&t�e����_5����6�t��dB�r>����d��%��b�nr��r���a�y�^X=U(_A�A���2�S^N`������o�S�ګ���       ��Ż���w=���\f������������6��3 �+VTbb��▚�jKtt�c����
�1��Ǧ@��Q     ���fЏ���A�fPQ�Z��܎�i�֒��7v�J�&՛�ۑߪ���|Ř+����z�7��)�׮yMu*�)����u֤���M�6(�:�w e���l�2[J
���:[J230~ѮE��TщѶ̉���ĄE�!S��L���V�����C���K�i��	�ۘ�Q�7
        o�դ���M@��m�=��'�k߰_�Ä؛>fb���t��i��{]���̋���L"��� J�ڵk�������[\	>cʙ�2�q~�� |A1      .D'D+?̌еBjٙ���cݎ	A1����>P�O���ӏw�������{���גӧi�"�ӹ~gy������ w   ��{�ܣ@�@�u&�g���         �ӏ��.vY7�Y�>���\��:u����}��;=7�9m;��e}ŀ����-z��+���;fb��W~,g�S ���ׯ���H%Ijj�-�ѹ�N��1��Ǖ+W&D�Q�      �����|/� ��W�b<�ѷY_�|���j�W*�̍�w�U���U&,���Ы_UIԤzM�eZ���ߺvk{��d�Iy�i�q��^� �9   �G�#@�_v��zf        @Yզv;a�+�m��c���~�ai��1����<�3��>Z�~���~��:\���rf���M�j��� _תU+͛7O�N�P����ȑ#�����Phh����N�ȘǦT�VM���'��}�      �p4���ӓU)��9�m_��V�[���ɠ���h�����W%UNHLǺ���l(&Lh����tf��
լ;f�9�K~����S�N�m�o�K�]b�QP�   ���퇫N�:.��S�5y�d         eѥ�.u�z\j���f�Ж���s����9Cb�d&���i?-p���̕am��D0�]t�"##�vN�Sqqq�DEE媯T����$��Ք�+
��     ��Iy�zt���g�R�����}�����<S�B5ͼ}�.������Q��f�9�D��丧�=j�D7L�A�)��u&$�����5�{���^��\^����*   ��G�=�n��%��0         �'�I�\Y��c����8R~���֯ڿJ/����O>�ۦ�f�bʕ+��~@�r�9��v
 |]�^��k�.��e��ɶ8p W����BBBN��T�R�t�L�5l=���     pc����
����e^{��5R���o�mD[}1��8�Fe��VIѪV+�8�G5��@%͕��Ԛ����i������W��i��sԩn'��۷i_��?N�P�cp��u  ���f��έ��-��         |��O���k=�����Y�ܯ�:�ež�z�׺��M��V��5[h��- _��]�j����ZVV����l���:����O���6@&'H&�)����7�b      ��o����Z+���$��{�׬���x�D�9��1��Y|}��

UIe��%�/ѫ_��^��,.�Ҹzc}��j]�����\����K��h�A�A����^/6%V{��
   ��d�3����6L���         �U�6t��ڃ�	�1}���n�~á��c^��1~�x�A1F�z�	�Pb���S111ںu� Lvv����mq�bŊ�Ccr�dr�� �      ��$jI���uQ/MY7�����A1�moS�#@#��TVv�|�y/�}QO�|B~��T�9��G�����h?�!����៫rPe������M{k���m�O�>�
2?�S�N	   �_��m(dDh��z���          ��*�(��U꺬[p�G�a&�2��ܙ�aj���b�
�ۧ�a�sյ��B PR�+WNC���˖- �9y�-�U�p8lXLN�L�*UN��T�^]��b      ���S����^�z�\vX�a�	.�+_!o3�sT�XM7u�bN�ȗ���RSFLQ��vi/1-��jb~��ߩ��x�zRz��jMBCl�Z��Wo��K���pA�B���b����/֌M3����no~��{�o���|��i�M����xP̰v�
�ނ�  ��a�;��t����S��z�ި��N̫������;         PVլT��m��Lg���<�m�{wy��qF��a&���c����\uM�7 �$��C�^�t�j�6ԂI�r:�����%**�:sL��� �5'D�<PZ     ���;�k�%�ι\�z�Jpŧ�{l�=/�
�+�8����6i����|�XI�\�������N�3���%QK�1z����B�g�������uQ/]}��
p-u܄j9H��M֛����c�U��b�a���_�V�Z�l�o���+��S�iτ)]���B�;o�<  �x4��\��)��Wtb�����         �����s%.5�c�]�wq[�+f��x�6Gov��	����aÆ���;�������� ���[rgdd�w�k��c�sfp̙�2&`�ۓ��DP     @f�13_A1&�Ą}|��K�m�_�~*NT�@��_��{]//xY'3N����[:ܢW����ЈB�a���8j������|�ؔX��?2���z[�^���V��!��h��#tŅW���f��ۥ��ڏ��OW}�9�s�l/��;:ݡ�]G��j�8ըTC�u��݋=Ҟ�ه�x�?�����  �o3���7۹         (�*Tt����{��w[�t�Ry�G�p���� %YHH�Z�l�.++�ɘ����X������5S�sOp-55Ֆ���\u�Æ��Ș ��P��ի+ �h���FP     @�Ĵ�|݀4��
�q�9t]��T��;�뙫��moӘ�c4u��b�����GꉞO�I�&�j#Ù�i����oj��-*&��՟�Һvk=��Q�h?�����n�L9�rB36ΰaE��./RpOp�`]��
���v�����;���Ʒ��   |����?�_��"         ��s�������h�g�����.O9�|���� (����O�N4j�(W��A2���JLL��1&TƼ������l���i�5S���r��>�M1A2&P&�qa'�
��     �<�g�۠br.=.�Nu;í5E���]�:���|1۞2b������[��&�����d�o�E����5�Q�R�Pmd������Ϲ�ԡ�C:_L8ͨ���/��>/����V�
�t�e�ْ��e�+s�}�����S;��A5iYi��1A?a�a�Q��Z�j��m�.���7+�� _0��P��9����9F��&/36�   |������6�         ���E�X�#�w��c��m�����\!(@Yvf��+&�"%%�t��)&H�<7%&&F�����DGG�3�oHH�=~Mx�	��Q�����U�re��~L�A1      ���O�c<��I�<��ۼ����j4ӄ�&h\�q�n�w���l��1W'3N�=?u����h|���V蠏K�,�#3��C��+��u�7wi��	zk�[�ya�"�i~n]�w��s����p;k�/1nhs�>_�y����/�z+����#[   �s0�>[�����}K>&          �_|j���CC<Ҿ�$ϝg��8�<%)=���f24�W�L� 8���A�DDD�\ƄX� ���d%&&� ��PSL= ����:}�EEE�Ug����гBdrB��U����@�AP     �9�0�mG��y���\���שQ�F�:�ªZ���(_R%����N[ҳҵ��jm9�E�o�?���8{#:9=�._9�����T;��.
�HM�7Q�ڭuY��<2�Ijf����	}���:uJ�hc�F]�ᕺ�˽z��7�Mlo)i3��q�E
����U�դW���x�� �(V�_��f?�ń5�����n����D
���z��#          �%�%�|��7,�(�Lgf���\���:31��7�)�r��;��r�r
 P8�����c�,���l�Ell��1�s^3�}�_6PR9�N�!2�9fs�cL1A2&P&�q�r��BP     @>�����9�s�9�J�Wt�������dCV|U���5�f������<�fP���͒~�@�v-ҔS���ԵAW�����.*���C�j�Ǔ�k��� �(LP�) �/:1Z�-zM          
�L���OլF3;�[a���m#ں�_h�<�B��Iגғ(  /���?FѨQ�\�&�"11�Z$''��&<Ƅʘ����- ����jKttt�:s̆���cքǘ���c8<<\�˗�.�b      �a��z���T�R�s.;��0}��s����oǯ����~���6�[�ݪ��T�$ۏm���/ק7|�[:ܢ��$���b��O^�u�����P�.{���;             ����Lg��;r6!/E	��\���qgٞe����._7�# ��q8�C(�1�&4&��@���$�8&&F�YYY������\����gǘ�*��3�     ȇ�������7._˿5�--ܹP΂����6׫E�Bn�.|U���L��1$=+]#��=�{�l�gmXJY6��P�AaS��|�Ӹzc��+3�̄�             %�3۩�w�e����4�)���-�Y�x�byR�*u]���FP �:LaJDD����  ��������A&P� �a�7S���s՝"cJ�*Ul�L��>��4 (      ��/�G�=��J��\�Y�f6���9��}?���!�Gg=������΄ܘ}�X�1�;��2�V��C��]��U�Z�b@E}���X�P�3AOq�q            ��h��ͮ�bZP���xe��l9�m���vr4Oj�������	 P��ɸ���e�bLpLll��1�<6��`��:�(�K�
�q8
��1&<����T�^]��#(      ��l/��|��?z�C+�����~����]v���l.��韟.!1g2�C���z��7T�]��J��d�&��x�e?����ݺP�9�tT�^�o            @I�8j�njS���$\w{X�,|��m�>\M�7q[�p�ByZ���._�<) @����:��Q�F��N�mx���c�dL��y���) �g�3sl���ބ=���� (�����     ��pŇ�ut�7Fs���ӔS��펊:���6�K}_�6n�8���U�Fo.~S!�!�{�J��o��}?����V�[�mG��]Ƅ.����_c�URz�             ���9���*W�\����zZ��Mҡ�Cj��W�=���f��:������Ƕ P�9�<�(�y��$$$ؐ�Մǘ�9�	��&55Ֆ���\uAAAjР��7o�6mڸ�.E� (     � 2��������_�|Xp�f�>SW}t��'w�L�����+��
�3k�,=7�9�f/�{A�j���m�WI�}*[��,ӂ��t�R�8�CG��*+;��PӠjum�U�[V��}��؄�̹k����]{c���g�)Lǵ5�tէ            ��lO��>�Z�ֻ4W��5�����~%�%䫽�/�Y�/���X�1N�Iu*�Q��.�"�G
 ����ȡ���ԭ[��2'O�t ���` (���4m߾ݖ�˗k�������A1      4'r�����[:ܒ��[�n����M�>�É�Ϫ3!1_������"��	�m�m6��43����P��բf�&f���v����w��Ɍ��zd�-�����m�k�r����V�����Ճ�?�o6#g�S?����1W�)�{5�5ws�m             J�W|�2(�h�V��_�۾�M��7��Έ�#�ٰ��\f����'�I�\1�m>�Y  UŊmq^����+<�̯��ɥ�;�	ǎ����C��iӦB�"(     ���1{�2�Rx��7! �����kîzw�j_���?��0�|�jR�%�'��w����(_u$�^^�>]��R3��ofz��`;��\����V����2Mo'�mhWo���"��7����             ����S��>���s�b�b�<�F�o�^36Ͱ�����W�O�Ck�~�wt�C=.��v2��zg�;���+&$&>5^  x[@@����mq��t*%%EIII�����������L��	��׌����ot�m��nݺB�!(     ��'ם3�Ԭ;f�\�r�Z�I�&��}q�lPF��ZBn�.|������?5n�8{�ט�s����/)1-�Hm}��+���5M͐����C�5v�X            @ia�s��=FSo��v���ݍ�������nyR��uԣ�뀚Ż  _�p8bKDDD��S�N)99نǘИ����P�dP�deeٰ�|�1�x     PH?������}=p�Z�~X}��mG���/�,29C�U��m�+�\���F� O1�4�am��[Nf�Ԉ)#���.             (M��������-z����$;������V9�.�D-  %��d6'H�nݺ.�IMM=+<Ƅ�$&&��9y����ߋ/��W_-�b      ��ɟ���/W��vŲ=�2o�<ܱ��eeg)%3E5+�T�*uբfui�E�j���_����#�)����L=:�Q-�w��~+rf;��q����i����7�J���|��"�G
             J�S�Ni��QZ��
5���������:�pУm�A�#;�tY�}*�� @�lK�Z�\�gee)))Ɇ�$''��������0���l%ɪU�ԵkW����J�h!      ��������W�F�^ن	��r�����؀�����\��z�k֯D��,߻\sw�UY�p�B-ڵHW4�⼽��IG5���x��D��ʏ�x��=����޵�             �V'RN���}��E�V�c��W_o�Z�vM�kԼfs�u��`�� PV���+,,�W�N��1�1&@&���9ń� ���[�l�%�\"x��     �q���i�C���*�(�Ѷ��n�h"�Gh���8�a��/�=]��=��Qx�p���s�
�s�>�e.;/�^�o�ݗ�����w�����>��cf��z�χ�             ����G]���n�N]�w)R[�N�ҿ��K/�{A����ϻ��vӷ  ��p8T�J[��w������8%''+11�ɘ�9���m׮]��b      <`鞥��n�F]2�cm�٩��w����Ej�`�A>�ڢ�4���z���Z��|��C�m����(&���7���s��w(-+�X�w ��~��G]��:�����(+�t|             e�����>��������U	�R�6v���?>�Y[g��7�Nu;��35�o�^  �`���mq'--͆�$$$��z��I�v��{}W�\9���     �������t�4��!1gJNO�+_�+>п��K�_v�~���V}&�ϧ�>-֠�q���9��?����屠���1��C             P��ɵ^��u����N����]D;���s���h�<NY?E��N��]�_��ۺ��W���  �g�V�Z���t:������8%''��&@&66־fe���Djj�RRRT�bE��1���b      <džk��e�jc�FyC|j����&�����~�K�]��)53US7L�gƦz{��
	��vL0̘�cl'��a���JLKThPh��Z�oe��             ���K��[K޲�Z�jj_��Wo��A�U1��bSb���h��*%3���)�?P������  ����PXX�-���SL�LRR�}���UZ�b���	�     (��nCX�W)R;&8��/��L���/�SW>eg�(�(��������'9=Y?l�A7_|�׶aBUF��	�'�|1��,ڽH�Z*r[ff             �t"���o��d�����   
'88ؖ����'O�T||�r}5�͠�)EB~�a�      xH��l�ڿJ}��)R;S7L-�����,�4�%���͸u�Uk��67r����s���v��o����u���1�#A1+��                ��*V�hK�:u\�gee)))Iqqq���Urr�-�ÿ́ʘ�OA1      �bߊ"�|���uש��5�I�b@�n��B\3:���ʕ�h�&h䴑��a�|��]��܆	�Ys`�                 矿�����li�(���N�S���6<�|�	�1A2&`�<������     ����^���%;o�q�q��@���=��Y���u"J{b��I:��G��U�Vk����j����|��cە���J��
���Û���$                ��s8��d�IMM�29ńʘ��ĉJOOP     �AK��)�b����>����ԩSz~���}b�>��c8���-G���q���<��}*$�0�����ְ[���y��                �����DDD��7A29�1�������!2�)�#�6�      xPzV��휧!��j�u��|��K�?��w�TH`�׶���6��?��鱶���W|(_�9zs��bfo�-                @ّ$�F����ʲ�1&<�ɘPS�c�A2(��     ���.tP̦�M�w-��]�_��Ea�a^���c��<3a��k޿�v��]�u�'ת��                @�����*Hf���v�����'O�`$c�&$$(##C��!(     ��fo���S��+�W�u�NDɗ� �+>�B��J�o�P�!��É���ƌM3��̇�ˊ�����g{�                �_���P�V-5l�P*TP����W��i�dLxLLL����l�LZZ���FP     ��I:�uשS�NZϤPG'F��l�ޤ�����*,8̣m'g$�%�%i����֩��|�ʾ�}�^�3                �	��������7Vpp�U�jU5j�H��???egg�����d�Ή'l�LRR�}nƊ �DP     ���cf��b����._�1z��~�W�РP�����$���Z����t����̐�;�r�P�e�iN�                PL�KVV�-9ʕ+���[�֭k�� ��	�9r�v�ޭ��%$$��>P�      x����K}_��˯��4����Wk����]�*���6S2R�R2��1�C7L�A1'cTĦ�j���VbZ�              (I���T�Y�@�TtT  (�&�ؒ#55ՆƘ�h�"egg��b      � �D�VX�K�]��uҝ��u�v-Ҩ�4���
�q�b 7-�R)�R��{j�SZ��J��'���(p �	d            ���[�n�b�����tf�h�QM>j�Mn9�Em����Bޚ�4U��zZ'44T  ����Z�j�����      /�z��
��+秒��_�~X}��7��m�q�2/���,ݳT�.{W%��0P�����$��6[         ���;����?���� E�}�ZQQ����.W��^�.�k���^[�����jk{���*j�D�wqd	$�$�,��NO������L��p���w��y�O{f&�  �3��%6�id����c�?���a&]�  2�P   �Z2z���;WFvVv��w�����~�n�k��᫵OQ~Q��J
JZ5�zYu�:��hlj�L���Ԫ��M�/j��         �����1���o�o�~+~��c��1���  �eB1    k������G�ƾ�m���y]#S$o֞zש�Sߝ�_i�UާoI���-m����'.M_�%�6n���         h߶�`����w�+����>%����   V�P   �Z4�͑-����GIAIT�VD&(�.���~<}�ӑJ�Vi����*�j[�޲�s�@���}d���K-�^ONy2         ����=�8��8c�q�k7  �j�b    ֢{޺'�t�"/;�E������9��I<��3q��7��=����-�ky�3jMH���uu��
s[��g�=��aY         �9
r
�cnJV��O�:  ���   X��,�'>x"��շ[4�oI�xg�;�I.x����oÒ[�v�>�_��ߟq�����=�����U�GM         d�K�]5q���  �:B1    k��7G�8�E�-���LRQ[>ra�v�m�^ۧ�Ol��V������_i��kP�����_F&�ѥG��Ϊ��~�l         t&sω�'��A��.�%�K�?��q��#+�ժ=�>��x�7��� @gWPPK�,	h	�   ���w��e��7EWf����Lt�;�?����ӆ;�z큃�Y�7?�E��N�O>2�&=6i�ܻ&��M�        ЙL�5)�w���=J>��z[ƶl: ������k�dge����[��*�K �άw��1}���   X˪�V���&�^��ҹ۬�Md�$�q����S�?���6x���:h�Z4��'.�L׿G��}a�        @���^������[ґ�C�>4~���b����uw�8�������� @g֥��/L̈́b    ��;��ӢP̎��9���~id�q���sӟ����ݪuC���֏9���Խ�{��!+��������L�i�M[<w���        @���nI�|sd��8:���q��.����=��q�sפ/� �Y��P   @xg�;-�W�S;��9^��bd��>��������d��I��W<}E�O'�|B����\����l�g�ͫYV�L         ڿƦƸꙫ⽹��}'߷�XLIAI��N�׿t}  tVYYY-%   �&Ϟ��{��;cC1���hL�lB��N�Zw��ƈ�#���)����n��tά�Yq�[�D�K�R�Sߖ�{y��w���!         ����H�s�9�����O���  h!�   �6����xW<}Ed��^�.�����j����q�GƘ��Dgw���}�_�[^�%�5,�L���vo�ܷ�         d��_�>��������c{n�g���3T/  ��	�    ���3�g�&=6Y�ܽ��%%QQ[�hԛ���\����ZwɁ��}��Ʀ��R�T\:��ͽ��ۢ#H��o�W>y%         �<MMMq铗���c��XvVv: s���  ���b    ��S����8m��r�s�-��GG&�^V��q{����[�n����cw86���ߣ�:l��b׍v]鼗>~)>��At�lyH��>9��          3��6.fUΊ>�}���N}w� ��   h#I�%���w��nƆbwL��ա�Ĉo����{8*j+����5���U-�;��Q��e�Ű͇�h����1m��          3555�����;��Ƕ�`�   VN(   ��$W�hhl������Vߎ��ca���D��|-��ߣ��mX�a���ŏ��(:�K�]���t��7�������l�(.(n��$�        @f{z��+�lT�Q   +'   �Fʫ��O߈���ҹ9��׿t}d�$frפ��}/h���{��G���Y��q���h��&�'�>����]On��'�<         d�)��xr�9  `�b    �И�cZ�I���)�I<��C��I�R1򄑱��w�Y�����խW�>qtdge�h���>A�.=�m�j�ܪ�U���         �mA��/.(  `�b    �Н����EQ�$(���{����(y��QRP������tO��k���*'+'F�0:���k񚧧=�I���9�-����X         �m���b��#+��M�  |5�   �6�Y�g1v������?g�s26S�X㦍�#�9b����q��7�F� �����I�Rq���ƾ�m�e5��'�D�+�)�s�yn������        @櫭�]���3u�E��b  ���    ���^��š���=*����O}�蹏�[�PL�]N���8�3;\,f�!#�G{��Uk�h�����钿wߒ�-�;�|F<��3        @��ѥ�
�746Ĳ�e  |=�   �6v���Gyu�W���E�ٹ�����9=2ѫ����{$Q��
"�=x^���\:���ɐ��z�k3_�LW�_�wa�����-���
1         �W}v�zYu   +'   �ƒ73����.n��Sv;%F�-�(2͛��������z/C���s�oI�8i�IQ��&2U�}��a�3��J��g������^�z�h%���         t���^��Us  X9�   �u��箍���-��J��f��EC/�SF��&��|���ؼ�櫽���oG�rD�_2?2Miai����c�������Y#���>�������Ƽ�y        @ǰ��{�����>  `�b    ց��������9�E�O��=qt<���i>��fB1�o��FL8wB�4�xz�ӑ)��d����;�����GCcCL�?-2U׼�q��n��TV���5��U�
         :�!�Y���t  ��	�    �#W?su���Q�[�ҹI\��co���!�,��dM�y�Q�F1v�ظꙫ�G/JEګ��ܸ������.�����kV嬨o��L��G�wl�s�Ͽ��[��
W�        �(�v����������   VN(   `I�W��2���j����֋�'������Ɔ���sMK�9�9?������?��'���ЁC��C��m7�v����#S�h��	;������.�_>��         ��8}��#/;o���:��   VN(   `�ݸ��ɻ��nԢ�C6?�����'����b��=�l@�u�]���Oƅ�\o|�F�k�m�]��[��om��5��ܪ���v�h�����o՚��^�+g         ��E���]����U͋�g�  ��	�    �C�˪��4F�0��k.9�2oJ��8:2���Ek�: =�MW��2��hjj��4t���ɐ�ā��T*���_R�$2M�.=�!������:j���?         Cnvn�s�%%+|��w�Ʀ�   VN(   `=it���i��}[4?���r�-��O�/D{זo��7`��HB:#��&���羿��7�l`��1q܎��V�mkSu]ud����x������Z���G�5�         ��[~�����=�l6�+����  ��P   �:�����uJL��(.(nњ�������^�+�Ο�Y^v^��sP�A����fM���>�|�L<?��(�._�}���|��7⛛~3�;m�S��L�ZJvVv��/�7ܪuɛ����X         ���⠸��k�e�*/}�R���+  ��P   @;0�|F��s��cnn񚲮e1�G�b���׮c1���������>=~�Ϗӱ�|S�M�)��G>��UuUQ��*��-��y]�K^�(�/�^]{�f=7�e�����$��.$�'S\w�uq�և�jM�s9���        ��շ�o��1q�NǷ�bl?{�g  ��P   @;q�k��w��N��-^���:����X��>��hÒ���Je�c/������$���ޥR����1|��Z������t�        �/��΍ny����H_<.� [򙶒����j��b�������:�Zo��g�Z��o�g?z6  ���   hG������l��ܬ�k��I�b�^?4ޙ�N�7�t�$X}�)��"�Y���#���qZ�����_ċ3^         Vl���c��Xt��O���?;  �hhhh)�   �v���<���x���(�����/Z?^<��8�������d��	Vߖ�m���JcSc�7ɕjn;�8v�c[�v��Q1b��         �s��d~�C���2  ����	h)�   �v��9o�I#O�1'��T*��u������>�Ӹ����=�ѥG��g�`�u�����,�Ο�I�.=cԉ�b����^��goƩ�O����         ��^>=�s�wbʼ) �?UWW��P   @;t���Ņ�\�;�w�Z���W}�إ�.qƽgĢ�E�.0��Jek��[S�o?��7�1�=��ؤ�&�^;s��8��âz��        :���}(N��Ԙ[57  �_s���G��P   @;u��WD�.��}/h���v<.�'�:9���t�+���9�osx\�������I������^;�j^p��X         ����qѣ����{  �euuu-%   Ў]�ȅQZP��l}p�_i�;|l��ſ�ŏ_���іv�p��ِ`��g�}b�����缽ΞC��>�@̡[�J�+k+����}         t\/�x!n|�Ƹs��aY   �O(   �kjj�3�=#R�T���i�^��ʊ3���xl\���q���GCcC�m9Y9�ף��~ެ9���a��Q����N~���zJ\��+���t��XX�0��x��7        ��#���G��?�����)O�G>
  `��   h����1�Geme�d�OVi��]z�uG^��}N�xzD����Q�PkKٹ����w�6Gı;�&�j�s0���!���6�i���|��1��bҬI        @�3�~��h/���U.�����]9;>Y�IT-�
Zfi�Ҩ�k��+'ׯ     ��+m������fa\v�e�J�Vi�A�ō߻1.vI\��u�`̧���癗���Ĝ�����#���t�M1s��xa�k�\C6���:p�j�3�|z�aXL�?5         h��~7�|C�1�����h�
7�S��  ��P   @����c��iq�7G��.��φ%��ߺ<.;��7m\��8:���d|���Uگ{a�8n�����46�q�w�˪c^ռ�Mj��Dm}���_%%��ʊ��z�G~N~�k���1���q��+�7O�f�^��[~�8~����gŶl���=7��8�֣��o            V�P   @��k�]�Q�Gq�����/�#	�84=S�M��?�gO��f����Y<'��-Y�&	��-��{��7�=��x�����"��Es��ƄO'��>H�=��'�>Y�hI�.=b����c���6�o�m�]z���+�JNVN�l����=�ǟ_�s���m�ߪ�٥g|k�oő��6�Ѭ	{�oqƘ3���.            X=B1    ����ǎ��1n=��8x���ؾ�zJ���fYM,kX���-�Y��|5�����&Ifm(�.O�w?�K�%�m7�6o28����m��";+;֦���C��s�������x{��1oɼt'��%!�$ԧ�Ol�}�ش禱�;���v��{m�Tj�=�$,t�}g�-��           �?566Fuuu��Ԥ�&#9-%   ��� �!;$��缸���!���0�0=ړ$���{���>/~�b446��s�I�'�<�z�WQZX��/t@:�q������Zo��X�&͚��ql�?��           �� �xkVVV�k}}}��եc0�/�y���g�}�<������b    2X����㯌G�4�������v�����1�8>Ƽ5&y���Q>#ڻE5������G�b��M�	;���t|�EGR�P�?uyz,kX           ������I�$�D`�.]����dɒX�pa̟??�Ν����6	�    t ��y'�ip�5���Ձ������(>��,nx�����[��G�J�>�O>=~��O��]N���J�E�{��g���ώɳ'           d�����ڵk��0I�%	�TWW�{��/Na-Z��� X��b    :��Ɔ��k��	wƥ�.������΍L����c��#b���Q�PIeme\���q�����=��/�e���#2ʹ����G.�{޺'           �=�������t��{���Leee̞=;},��	�    t0�̏3�=#F��wa����-�[d���f�ŏ_��~[465FG��~i:sפ��/G�%������}?�x����;���>           `]KB0.L�� L���ҥK2�P   @5�|F�gx���y���?���1x���^555�/��?t~,^ڹ*�sω#o=2.zQ\r�%�J���I~&c�wL�#�M��y          @[hhh������,Z�(�����***���.���   �ખV�-�ݒg�uF\u�UQ�S�I�����;�-���謒�ʯ��u����%�.�������1w-�(           `M���_���������!��X�ill��b    :�?���x��c�c@ـh�������~�j�뱿��������^�O%�����>��XZ�4           `U|1��_�Lr��Xr?�;���b    :�	�M����s�x�q��G��'�:I$���G<=b��b�,�SF���}_           �ש��I_������2~I�'�9�>�   �N���2�w���ψ��:�s����x��������j]�s��{Ǳ1�|z           й%DMB/��K�5	�|1S__��'   Љ���?����O����ox����r�s��y��y�������.           �����:�I�/�H0����c��e˖|�.]�DG�J���   ��&|6!v���q�a��ɻ�ܦ�2oJ�e;�١��9�rv����#�=           t�����/����ͣ��"�I.<
����0:��hǄb    ��������?��G\���w��mr�n�݂/;~����|wM�+�sF,�^           d�$��^�Lyyy: ��N�%#�/��TZZ��R��hǄb    X����g������#�9b���[[|+^����,Gowt��+	Ü}��1�͑          @��dɒt�%��������R�~���!   ���[57����8r�#�G�1��Yk����ꙫ���"����ٹk�<wN�3�}�ܘW5/           Xwjjjb��GUUU,^�8}{���QWWОm��VA��   `��|o<5����+�=N�T*���ѻ[��������"N���8|����9f�ψ���x���          �����!***bѢE��H0�ǒ L22UQQQ4(hB1    |��ڊ8}��q���5�_�n��?Ǚ{���x<��Cљm�k���\k��,�����*~7�w��nI           �����ӱ�$�R^^UUU��N�%1������j�}������m�    �R/}�R�q���]��|ylP���;�J�m��{^�g|0��ʺ��C�>%%ke��'��?t~|���           ��jjj���"=��/����ɨ���6�`��y睃�#   @�465�-��c��{A���9�-��ٻ{a�xb�1����ӊO�3)�/�Ny �X�{'���=��x��g          �/KB0I ���jy &�����򨭭��
�裏N_@��#   @�,^�8.z좸��k���3�:#
sW{�~�����O���ib1Ih�>{n���w�g���.���{8           :�����񗊊�����OF}}} �STT�w\���#h[B1    ��yU��'�$�~��p���N�.�]Vk�-zoϝ�\�~h|�����zv������L�51.{Y�;���           Yyi�|1�|;��466��4(���oGqqq���b    X-�*g����=zQ����q���cÒWy�Mzl/�����۾�|�LtD�{�G���ؼ��kd�f�W��"z�!�          �è��KG_.\�<���(LUU��P�Z�a�w�m�Ql��ѷo�`��   `�����k��&���8q���o��n��*�Uֵ,�����1��-���ЁC������խ�j�S��:FO���1y��           �4555����ŋ���<I�0��d$��``����^��ѣG����o'���,����C(   �5���6���_�c�~�ǩ����pl��j��������c�M����;+��-�L�J�����<.9����^�}&|6!������	w��<           �U�I�/�h�4�O�0����}�����/�Hb0I��v�;d�    ֚W>y%=��ǹq��ĕ߹2�vo�'�zr�����ߏ�f�����q�17Ő͆����@\��%�P          @{��L2-Z���$c���QWW@�XQf��֋^�zEAAA�1�    ��-�[7�zS�5��x�'����U��E�t�Kq�s��=�_Q��:2AV*+��9<�8�(�/Z�}F�92Nyb446          @[hhh���ʨ��Jm�����oWTTDccc m#'''�����=z�C0�Q�$���t|B1    ���g��p`<q����dgeǏ��q��q���=o�MMM�^��o����]6�e��5q�H          �������ŋ�ї$��D`���ǒ���3��.��$#��$Q��۩T*�܄b    hS��|-������>������{�N�+^��B�������/E{2�l@\|��q�N'���7�rc�>�t�          ��jjj���*~i�$�d$ǒǄ`�meggGqqq:��`��Ks�gϞ����u�b    hso~�f�}����i���/�b�&��ų_���>�?uy��6.֥�e����<N�����Z��ݮx������          �P�i�4a��'a���� �^NNN-�����+=��%%%������b    X'�Ο��48�?��ح�n�����O��g�7�|C��8*/]m!+��6g>+�����U�X������^�.          �Ω��!����%��hѢ��d̟??���X7
���QZZ���4�N�Rk�P    �����1�/C��cn�cv8f���e�]���C���ߺ;�|_��:6j��Ě��X��F��w��n��ѱq����ދj�1�OLy"          ��+	�TVV�0UUU��I���<}���"X7������8~I0I��9
SVVyyy�P    �Tr9���b�g�7�&r�V�%�n����� =��U��)c�ُ��W?y5�������Je�������{�77�f�;`��[�7ִ�f�G�vtL�7%          ��V__�/NG_��K�I�7K�755��.��$#��$Q���Ʌf���   `�K����xi�K1򄑱aɆkd�.�]�ЭM�D}c}L/��,�$>Y�I̭�u�u��n�?��u�����^�=zu���ŀ��ck�M��g�wV:�          d�����>}z̜93����HG`jkkX���KIII:���/�`�QPP�i�b    h7���\ls�6q�!W�i{������ʉ�eӣ=�W5/~t�b�[c          ���/��ҥKX7���_��In'����쀎D(   �veQ͢~��7m\\s�5�^�z����=q�g�ܪ�          d�����뮻b����}ݺu[a&]�v�L�b    h�FO��x\2�8s�3#;�cT�?\�a�������H           ����!F��q kFvvv/����.��E^^^ �$   @���fQ�s�9q�+7Ư�U���J�"-�^�}�q��Em}m           ���G��UPPP���4`��0�ג����]hkB1    �{�gO��n=*��}:s�ևe̋�kƟ��S\�����          ��f͚o��F +VXX�/!������ �O(   ��1i֤8�#b�w��� �����ɏ�hʼ)q��7��⥋          �lcǎ������*'''|I�/��b&��<�]�+    ��ٛq��FIAI��aq��'����T*�N�WEmE<��q���SӞ�&          t.��ӧtt�����K���1�u��}��b    �XI�%��$c����c�?&����o����k���iŧ1n�x��G�o�#j�k          �X&O��B�tYYYQRR�<�D`�C0�������   �Cx����WO�*=��u�o��F�;`����ؼ��ѫ[��>G]C]|�ࣘ8kb��p|:3u��           :��3gd����(**Z�)--]��ݻw�q 3��   �gIݒx���ӣY���1���X606�i:&���%��u���Xְ,��VŢ�EQ]W��g��9���ySc�����          @�2k֬���!��L��]��1	�    �),�Y�~�jz           �TSSS��������(..^�)--]�)++���� :�               �
uuu�����.��$1�� L�5�ĤR� �"�               �
"1��/�`����իW@k�                �����t�%��$�$��Ib0������                |������d$1�$
�|;�J@[�               :����())I�_� Li��$�

�=�               :����(**�R�w��ѳg�t,���               2^aaa:��<�L�i��J� �	�                �^vvv��/I &��4Ga���"/// :2�               �](,,\IF�I�0ͷS�T tVB1               @���1�޽{GYYY:SPP ��P               |�����urss�ї�Lr���t����� ���b               �+����&��*,,\�IFs��v*�
 �,�               �]�v�����L�8N|�b�9����� �m	�               ���h���wމ�&'''�����޽{GYY��LIIIdee �P               |����gd(&�J-�$��L�����  s�               ���n��b�رQ[[�Mvvv/�����.�����E^^^ �1�               ��Hb+{�G�?~���K�.��/I拷���"�J �P               ���{�|�A̞={�������������FAAA �P               �Dvvv�p�	q��ǜ9sZ�>'''����% ���ݻw�q �:��               Z�k׮q�)��s�=���j,]��_OB0I &	�4�`�o'k`u�               @���������o̙3'#???���� X[�b               ������O�> mE(                ���                h�b                 �9�                �vN(                ���                h�b                 �9�             ����݆Jv���3�qf�I�E��Z��(V�|�����Kɦ.jC[(�鋢/��R�j�m��aq�!�I��c6�4�<h�n��&1���n��y�Ng.�U�Iv����|��̙��������  '                �8�                ��	�                 $N(                 qB1                 ��                H�P                @�b                 '                �8�                ��	�                 $N(                 qB1                 ��                H�P                @�b                 '                �8�                ��<�~����U*��fB1                @)�������3��2�z=��P                P
�f3:�Nt�ݟ\˲,VVVvb1�L(                �6�Y����/V*��ꪫ�ӧO/���׆�)��߿���ػ܄�~3&                L�޻���/��                �M妛n���q��T���j�����{�ޓY���Ї>�dL�                `������O]�����#��N�V�0<��Z�~�^��:�~���~$F(                �9��`4�^��×���q�R�7�x��z��sssy�С�F�b                 ~���g����8���7�x����ڿ����ַnM�{	�                 <��`?��|tcc��o����]s�52�`�P                �elooׇ��'O�<t��я>|���r}�              (�,ˢV�E�� 0M���n��� R��t�/\��w7�t�\}��o>p���^�+              %2
�,..���\  L�Q,fcc#��~�f�Y]]}��;>v���߾�뾵�k
�              @IT*�h4��y  L�Z��f3���v�1)���j�z��;��믿���\K(              J ˲X^^� J��=�ŋ���G�z�^����w=z��>|�n�#              %����J%  �f�YZZډŤ���W�����[^~�����XC(              ��h����\  �U�Z݉����HU��i\�x�߆�oߍ��b              `ʍ6M�b1  eV�ՒŌ�������㯻����B1              0�F� ����<R7bss���o��B1              0劢  Ұ���;��rK�����q�+              S��� @�M�=O��˷���hx���W(              ��h��`0�<� �����O·�=[����Xů�z�������P�������              ~���f,-- @moo��~J��n��K/�9��߿���s�t:������t��_��B1              P����z=j�Z  �I�ߏ�����̑#GF�ύƱc�^1�'��J��K�E�3~�(>�|�G�R�槯]�~�8��9#�{�śo���~���cL�b              �$���byyY, (�Qxeuu�Yc.����lxx��������U�^��N'�<����q�+              %1�@=�H]��c~~>�Uۉ��4
�loo����K��������xx�K��F�`?��?�y              (�N��3�,�J��s ����`0�c��xOL�����O(              ��]���=̖z�~㇣�U��3�.��'.<�����CO= �������Ȋq�{���`0����
�E�+�O(              ��[�[�5�-�v|�?���iT��]�i�����=(�[/���q$���Lj�,���s>�                �����EQ\��/|a��|��8��                J���?\�T&���������8��                J��}���o��3<�Ob��(�b                 �O�e�m��������
׌k"�                ���ĄB1Y��b\s	�                 �Uř,�&��Ҹ��                J+˲��Z;���q�%                ���I-\�Ҹ��                J+˲��(&��P                ��E�>���b                 .g�ɲl"k��                ��<��s0�ᄖ�Ѹ&�                J������S1�b                 '                �8�                ��	�                 $N(                 qB1                 ��                H�P                @�b                 '                �8�                ��	�                 $N(               1�۫����W `D(               1�A7y�xU�U 0"              ���|�3���D  ��               $��7��o�!^}ի @(               A�A/����/}�K�\h 0ۄb               uv�l���;����xY�e �.�              ��=r�����g���x�k�Y� 0{�b               ��ߊC�z(^������q�+����zt����  �O(              `J<p�8�/#˲X�.�Fw��l�ڈ��RL�(t \�              �)Sŋ�Č��Vw 0��b                 '                �8�                ��	�                 $N(   �	sO�E  �H�NU7�         �l�   J��F4��  �\ν�\���          �B1   @��?6��Db            ��&   �V�b5Zw�"�             �jB1   @)�<�w�#�f            0�b   ��)"Z_mEuͣ            ��   J�y_3��            ���   Je��B,�Z            �2�   J�v�+��            @��    ��o���r;�^             e#   L��Ȣ}W;*�             (#�   `���ھ���            @Y	�    Sm��K���b             ��P   0��O֣���             (;�   `*U�+�>юl�            @�	�    S'�g;��|+            �Y    L��{V�v�             �B(   �*�'�c��            0K�b   ��1wf.�6            `��    S��Z��]��"             f�P   ����E��v��<             f�P   ��"���VT��            �]vX   Ik<؈��            �,�   �5��|4N6            `�	�    I�=U��ݭ             @(   HP�ɣug+�^             �    �D�N����            �%v\   I�w���{b.             �B1   @2��K��            ��%   $�v�+��             �$   L\��G��vd�,             x&�   `��"��W�Q٨             �N(   ��}����z             �܄b   ��Y:���Y             ��P   0�s�h��             .O(   �s��J�O�#d            ��	�    {*�g;��|;             ^�   `O�ܽ��             ���   �L�d#Y             ^�   `O̝��ƃ�             ���   v]�b5Zw�"�             �%�   vU�͢}�y7             ^�   `�������G             W�.-   `�4l����            ���   v����|r9             �rB1   ��՞�E��V             0B1   �X��y��lG��            ���   �&+�h�hEe�             ��P   06ͯ7c��\             0^B1   �X,~o1���             ��P   p��?�Ǿ��             ��   ��T�*�:ъl�             �C(   xɲ~�;ZQ٬             �G(   x��}m_���            ��%   �$˧�c�            ���   ^���sѼ�             ��b��Y��۠�fw3  �r��W�����?             �#B1Dc�y��[o�� ���zY��hG���H            ��$   �`+w�D��Z             ���b   ����F,<�             �=�v�������J����;q��  �|���	�             0B1����?o�շ\�3��?��   ʥz�+w�D            ���    �)��Ѿ�y7             &G(   xvED뫭��y|             0ivz   Ϫy3��             &O(   x�������              B1   �Ϩ]��ʽ+            @:�b�sk�b��p��E?ή�  `z�[y��܎��             ��!���0;�O  �Tʊ,�w���Q	             �"   �h�ی��z             ��    �^���,             i�  �W�ͯ7            �t	�   ���W�}��              �%   3*�gѾ��V             �M(   f��=+Q�Q-             H�P   ̠��Y���/             �A(   f��ٹh>�             ��P   ̐�j5Z'ZE             0E�b   `Fd�,�w�#��            �t�  �Ѻ�է=
             �Fv�  �h<؈�G�            ��$   %7
�4j             �K(   J�z��{Z            �t�  ���;y��hG��            ��&   %���KQ]�?            @�-   e5             JB(                 qB1                 ��                H�P                @�b                 '                �8�                ��	�                 $N(                 qB1                 ��          `O->���� ��Yg�w6   ��	�           ���AY/ `����   0-�b                 '                �8�                ��	�                 $N(                 qB1                 ��                H�P                @�b                 '                �8�                ��	�                 $N(                 qB1                 ��                H�P                @�b                 '                �8�                ��	�                 $N(        ��c�nB��������ή%K��H��đ�(k�"BsU�Cq��=de�=$��D/S��Ň
���KC_�\�^JEӀc� e�4���tf��M��2�������`��{����
       HN(                 9�                ��b                 ��                HN(                 9�                ��b                 ��                HN(                 9�                ��b                 ��                HN(                 9�                ��b                 ��                HN(                 9�                ��b                 ��                HN(                 9�                ��b                 ��                HN(                 9�                ��b                 ��                HN(                 9�                ��b                 ��                HN(                 9�                ��b                 ��                HN(                 9�                ��b                 ��                HN(                 9�                ��b                 ��                HN(                 9�                ��b                 ��                HN(                 9�                ��b                 ��                HN(                 9�                ��b                 ��                HN(                 9�                ��b                 ��                HN(                 9�                ��b                 ��                HN(                 9�                ��b                 ��                HN(                 9�                ��b                 ��                HN(                 9�                ��b                 ��                HN(                 9�                ��b                 ��a�������Z���<�������7�                ��P{n߽?i�$�Amw����                `��b                 ��                HN(                 9�                ��b                 ��                HN(                 9�                ��b                 ��                HN(                 9�                ��b                 ��                HN(                 9�                ��b                 ��                HN(                 9�                ��b                 ��                HN(                 9�                ��b                 ��                HN(                 9�                ��b                 ��                HN(                 9�                ��b                 ��                HN(                 9�                ��b                 ��                HN(                 9�                ��b                 ��                HN(                 9�                ��b                 ��                HN(                 9�                ��b                 ��                HN(                 9�                ��b                 ��                HN(                 9�                ��b                 ��                HN(                 9�                ��b�Wt�ƍ��؈y����V�w ��c               0W�b�W��K/�͛7���b�                sG(                 9�                ��b                 ��                HN(                 9�                ��b                 ��                Hn�C1�$��fp�х��=Z{4���1�~��A��               `��:���_�����<����{��sq��.�4�¿|!ֻ�               �_s�                �B1                 �	�                 $7ס�����(6�{vvv�}O76�����                �0�:��v�����z�������?�eY               ��1ס                �i                 ��P              ����X,c����ȮSvb�� ���              �O՟��4?���cii)���c|{����_ ��	�               $�TY�k���#�G"� �!�              ��N�N����(zE  �K(               ����qu�j}� �wB1               	U�j�-�E1� �b               R�P���  #B1               	]�] ���b               �9T��� p�P              @2ã  �	�                 $'                ��P                @rB1                 �	�                 $'                ��P                @rB1                 �	�                 $'                ��P                @rB1                 ��u(������NpO��Ȯ��zn              �}{뭷��T*�LbvY�߻r��gǱ�\�b�׷������S�Nd����nM�s;               �!)��ceY>1���k���                 ��(�VY��=��=���b                ��U�ek���b                 ~��(ZeYNj�P�8|���X�S�˸2< ���7{7c���v                �`0x�(������Zs��տ��~����v���               ��(��㓚]����֚�P                0�>:��EQ��ZB1                �,;1��eY~\k	�                 3�wީw:�G'5�(
�                ��O�����bR�+���k-�                `&�ߜ��λ���q-&                ̪���_ׯ_�k1�              H��c��S/�Տbx�"�Z5v��4�T�S��_ f�����?��w/_�����CeY�����8�             ��j��h�����(�V�E�R�;�B �+�hY�1���G���y���Rr��o�\L(�*E%Z��G�����             ��(����z=  f�(s����v���nܸ�k��bB����q�'�S�P�R})��Vgk��             �t�V�����J%  f��w�v��w���o�}�,˿^6�y/��`��1:G�#�^o�z���?���F����l�              �EQ��  3��l�YF�_�7��d����������G���r?��A�0���0�U�V�'N܈1�             �0�8- ̺����t:?��������W��v���Y__����<l��ѥK�vc��b              `�E�z=  f����v����k����{�0T���a�k
�              ���V�{�� �A�V��w��^o!���믎{M�~�V�              �g� ��J%2k4뫫��4�u�b�s��/�W~�+             ��)�2  �E�w�F��W��P̜���+�^�/�ޗ�ZQ�             �F�~?  �E�w�Z�����O��A�=ס��}�s�x���J��F+����N�����#��ŧ�:��|L����ע�o             ��h��`0��3 0��nd�l6��g�9���P��G����g�����z��`��̙x�'���0MN-��g�>�l��             �ص��h�Z 0�F��N�---}cmm�/j����oeY���N̺�G����J,//              �cww7�V� ����ގ�Z��?^�z��/�������j5�|��8s�LE              ̞����&�` �,)�2677���E&������߭��=w�ڵ�5ס�^��~?fݱc�����/U��S�ܖ�             �h�(3
�4�8th�� 3`��t:�n���u2�k��������e^̱;�w���N̪j�+++q�ܹ��̂�?�w�L�s�Lw�            ��F��G�h�i�R�� �J�H���hii�G�z�����>��s��eǏ��/Ƒ#G             ��T�e���t �qi4�V���7o�|�����b#3c��j���Ĺs�               `��������F�O����$�A(f�?~<.^�G�	                ���j�~���^����^xᯋ�('y?B13�Z����s�Qr����?�3���&�$K���Tp��A*��b�Z�U+R����ފ�zzN�p@���{�-�
�E�mk�c-�F�X�AE
Jи���������|=��Ͳ	I�a^�9�3�������a~	�컻;���b�*                ��K͎���ʾ�ɾ��b��١���]}��Si��o~�bD��害�3zzz���#                ��r������XX?��o
�T���&j��ľ��|>�Ծk�---��v��o\~��b	�Y��}Ѣ��;����"                4�\.7��w���h B1�Pggg���DGGG                 +�P�2��磻�;���R�(                �A����p�\����]�v'&&���:::&�>����z�\.��e�}8�(��e���3zzzb�/                ����r�k�}qjj*�P(Ě5k�k���1<<�֭{����7B1�|>�����Օ�C                �-a���g]����, �\-�O� :;;���':::                �_�\�wM(�C*��GwwwtuuE.�                ��j��Z[�b��c�9&�?�����                �D(f�������]]]���                �N(f	��쌞�����                �g�YD�|>������+r�\                 �E(f�tvvFOOOttt                �|�b��|>�������\.                 ��P����===���                 %s���������r                p �b������鉎��                 8B1�I>��������\.                 K(�0��쌞�����                ��K(�*
�m۶8��3#��                �� s�tvvFOOOttt                ���С����=��y�G�P�W��Uq��gG.����ݻ��}��j               p@:S)Wb�<~Я?������}lܸ1�#�\.����߷K�P               p�:s������/�W�����                 ��P�ڲeK��/�rlܸ1                 ����<5�T�s��m.4��^����DSSS �cd�����U�=                DC�b�y���ΉO^��8�� ׽�{���               �H:�\Z����?�=���o�                �b�ُ�O8;n��8��                 XLB1s��rq��F��                 XlB1s��j�w�i��7�"~�����㘵�                �b�����h���o�u\}����all�                 G�P���ǲ`�����wo��                 8��b�De"               `ll,}�ј���|>�~��X�n]�r� �CM(               htt4n��������Zm�z=s�QGe�4�~���9 �`�               �Ƨ>����j�{���f.�bq& ���Q�t��� �"               ϡ\.?g$f!J�R6}}}��ZZZ���O
ɤ�L>� �P               <��o��yGb�K���ڵ+�g��r�nݺg�c��)���&               ��;v,�g��j188�ͣ�>:k=�b����蘉ɤ��`y�              �y�HL�R���T*e���7k-��g���I�z@�>�����'               �����Z��޽{��K�X|F8&Ee�1�t�����'               ���닕�T*e3�����2���c�������!               �Q�Tbbb"U�\�]�ve3�b���xLggglذ!�ʴ�� ��P               �G#Gb�T*e���7k��Iј4Oʴ��G.� ��C1m��hijY��5�5,�b��-˻885�Z-              X��^���/"���XL=$���1�ٰaC��,� �(:s�����N_��M�6����rE\��Xή��U145              ,}�\.8���jd���;k�X,΄cҤ�L
�ԏ�wQC�b               `>�$��T*e���7k�P(�ڵk�hL�ǤpL=(��ٙ��D�v               ��J������Z/�Y4f�ƍ��#2)*��� ˕P               �b�J�l���f��#2�����2��\. KUC�bF�Gb4?���,����]�}�Uk�              `yYY�����hooϢ1)��1��̆���% SC�b&�)��,�J���M�Z-              ���Z����@6����֋��L8&M
ɤ�L�XT8�:               ����T*e���7k�P(�ڵk�hL�ǤpL=(��ٙ�<_�&               x*�Jd���;k=Ed6n�8+"��[[[`!�b               `?��|��522��\�իW�d�s= ��S`&��@"               ���Ғ�b��j��0>>��Ν;g���^{{�L<&�d�q�6d�O�q�               �<���bxx8�HK�����lz{{�����b�ڵ3��\�ȤI�[`e�              �y{�B1,9�Z-�^��Y(��L���c2��Lggg�,/�Z               ��	'�?�p�rR�Tb`` ����g�555e�4)"S�ԏW�Z��#               �8�3���o�Z��LOOG6ώ�$�bq&���A�t���8�b               `���q�)���?�J�R6}}}��
��L@��y��u��pw              �s�袋�G�j���*�J�޽;����g�c:::f�2�8��pp�b               �9lܸ1�;Ｘ��;ؿR��M__߬����g�c��i֭[MMM�P               ,@OOO�ٳ'~��p�&&&��'������|���cRD��I�����b               `r�\��o�"w�uW �N�Z����l�R,g"2i���q�?a��              �J1��.�(^���׿��x��ǣV�px�J�l���f�
�,��1i��I��&              �:����+����������3344�M�Z �_�R�ݻwg�l)�v��g�d�q��X,,B1               p�����E/zќk)^122������٤�t-Eej�Z �O�ǆ���y���g�
���Lggglذa&&�nݺhjj
X*�b               �0H��H�u��Y��j5�W�xLz��cRH&f����T �O
:�{/Moo�3���|���g�p��ttt���G}t�Z�*�H�              �E�"�����J���E��I�t�w�ޘ����H1��Ed�b�8s�I!����r��CI(               ���H�y��9�SH��������,j��Ӥ�Z�����4}}}��R���=�ƤxL
�ԃ26l�����%               �T=$�q��غu��J��cR<&�dRT&M:Nׄd��V��=����w�z�o��4)$��2�s��P               �P�Ba&<1WH&�,���gb2�xL
ɤkCCCQ.�8�J�R6}}}���}�v������"PO�Ȭ[�.�����$               *��gA�4�7o�sO�Y�#2���ψʤ����D �N�R���~��g��{���=�ƤxL���cPG}t�Z�*X��b               ��*���/$���xL
�f��Z�t^��x����LD���w�z�W��4)$��2��\.,_B1               �A+
3Q��[��ZzHftt4����xL�ʤkCCC1==��W*����뛵��յk�f�j�ǤpL��ݸqc477K[C�bR%ijjj���?>��:��              X\O��%�����LL&M
ɤ�4{��r����{���w�z�X��WӤ�L
��w�rd5t(ft`4��b�R	X\�8W�lY3             ��|>�}�4�7o��^��btt4�]��I�������d �O�T�f���ߴiS�~��q�YgEKKK�8:               ,m�\n&$s�q�͹'�-�
�ԟ���8xO>�d6��ַ�~��/|ap�	�                �Z�X�fӦMs�W*�92������j�ott4>��ĥ�^�����%               �h�B!6lؐ���J�����fϞ=Q.��,���/})֬Y��zjp�4t(��o�ڦ��?T�_�� σ�c���X�&�=              ���X,f�y��9�GGG�x����̤����	�GL�H�����w�������y��hDu���T�����~"��z"               ��5k�ds�q�͹�B1�x�ӟ��)4+I�T��۷ǥ�^�               8Z[[�9�c�\�V�1<<�c����@����ώSPfzz:`9ٱcG\p����~B1                �Y>�����g3�Z��dR0&�c��)&S�J���� �w���8��s��O(               `��r�X�n]6���{J�R��B2)��ӌ��dG�#�<"s��                ,�b1��)��Y<�>CCC3��S`�V�J;w�̾W)v����9��!               ����Dggg6s�V�1<<�c����@������xjj*�@�@���x����
��%L(               ����X�~}6�S*���L}RT&Ed��޽{crr2��VJ(�V�5�&               @�X,f�y��9����bhh(���q�<�fh<�r9V�                �����l���T*122������٤�t-ej�Z N(               �C�P(����ٺu��j����31�z<&�dҵ���(���&               ����c�ڵ�l޼y�=�Ri&"3::���L
�LLL4"�                ��b���|!�z@&�c��L:O��k�Z�J#               ��Q�lܸ1�n�:k�R�d���IA����,��2����PLOO,7B1                ��B!֯_��\���lOSSS�)�JYXfll,���ٳ'��r�R#               @�H!���Y�&6l�g�qF���D{{{�j�,$SȤ�����#M(               ��W�¤I��ڢX,ƪU����#�?����r��磩�)�_.�cll,ɤI�ݻw���`���P                ,@��T*����Y�fM6�7o���B2���D�ٳ'{�,$�"4),355p��b                �I1�j��777Ǳ���ӥ`���x|��_���逅h�P�%�^[�[���Mg���=��x�֗�rv�c����d               И��b6�\.`�:s�Qg���N_��M�7��Ni?%~~���rv�On�               HC�b              �Hj�j���z͚��   �              8BN�{j?|�����=  ��C1ӵ阞�^��Z���J��ܷKQ-�]               ���������_�fM �k||<��~�.E��j                ���                 ,B1                ���b���,�P                ,��7
Ű`B1                �V�^�PB1                ���b�B	�                �"��r%                ��	�                 ,qB1                 K�P -ߔ��� N<��lֵ���ͫc�Q���?1��RLLM���P���c��c���S�O               �0B1 ,H[K[��/��oyy6��u�IG����z���x詇������|;{~���2]	               ���b د�Go��N�(.{�e���B��[�{�n^/{�˲y���Ȯ�x̿��_�~1��_��C;               ��YN�<-��į��W�P̑��1����lj�Zܷ�����-�y2               �Q	� Ŏ,����+�E,�\.�mٖ͇/�p������������(W�               �D(���t�I��s��<��Y,f�*4�/zm6�Fv�_��W��>{��               4���m˶���k�ug�.�M�XN�Y{L|�>��yo|��?7~��x���               ��L(�������揳@L.�;��"  ��IDATd����S��ȓ129��R���c�2���Y�&���Ѿ�=֮Z[:�dמ������s+�>�������ߟe�               V"��p�Q'���旽9�M��z�������ߏ��}/���w��]�����ӡ��De�ޫ��=�[w\����8��3�%Ǿ$��:Oˢ2�%��s���U��*�򮿌����               ��D(`+6����k_}m�Z�c屸����w�����1]�>$�kxb8�x0��|����\/4�ksW\t�Eq�)�y'�����������g�3>t����w}��}^               XlB1 +��_��cq�Q'.�5;�v��������}|��oFe�GR����y_67l�!V7���O�8^����/�u���=�Z}T�s��g�������w               �;���ӿ��xK�[�w�4��������{~|O�j�X*Ƨ���|>��|K\x����f�U�U���Ύ{�����/�7>���               ,gB1 +ж-۞s�};�9>���Xy,��r�_}��t;�]o�w���q�g��5��|��/               X�b He����s�����=�X�K�Y�&�E'_��?�O�0               `��h �j9���?���XI������柍��������Z��               +�P�
V����|�o�ۯ�'����������o��������\���               ����C1��R�O�/x����X\����߿��vI��?�����{��O|?�O>��ͥq�	�č��               �4t(�<Q�����/�J,����Y�}�$�P��n}]<��C���~������sqʆS               ���� �T�����j���               �;�                �%��C1C��X�[���c�������XΪ�               P���s��C1�T�����%�}`�|������7               �����j�P                ,�R��PB1 +X���Ľ?�7ƧT�               ��]�v,�P�
�+]������Ͻ=���;              ��cjj*`��b V���:)�����o}"~�~/Ƨ�               X^�b @.��w���������^w=zW                ˇP@���&��k{|�Ώ������L               ��	� 4�BS!���ڸ�E���>���o�}               ,mB1 ��M��=�{O|�Ώ���E�Z               `i�h`��B\{����b����}�             ��Da"FZF�5��|  �P�
vףw�U��*Z���{ɱ/�{~�����>��#Q��             �����@[<6~c� X���j������X���gS*�bzz:`��b V��v���������Wm}ռ{WV���\�;�uq�g����z(               ؿ\.�|>��������T�����x�'b�Ν�ux��b V�����q��� �>������<V7��w�Yǟ;޳#>���G��HT��              �HR����9Z[[�P(dA�J����1<<�E`���CCC122���j���I(�Lצ��{n���+n��x��wk�5�����������^?���               XIR&�`��ڢ��%�������TٱcGDLLL,6�������q����u_�
����	����?�����Ưߘg               ��R��E_ҬY�&�����O��سgO��倥N(��T�+q���~1n}ӭ��-/�w���_r}\��K��{{<��               X*��jg���b0�����ߟ�ki,wB1 ��]ƹ?7�9������bUaռ��;鼸���������D�j�               8�*�J���dїIA�4�L����g�P@�LW��7ė��Kq��ƶ-������7��x�������ձshg               <�R)��L����K
���4B0�_:���"��ܾ��V�}X���? ?x�q��ωkο&����XUX5���O�8x���_������              `R&�_�ԃ0�������5t(�_��;}��7m���zۉo��ν,����}UM�RS����o�/�Ǘ�+n�m[�ͻ]뺸�7��_��3���              h<O���b0i����r9�篡C1 �����9?'�9����k>-��y���E����q헯���9              ���R����P�??�xxx8j�Z��r�\�K��,�,��Jܰ�����_�[�tktm�wG�#nz�Mq��������9쟱\-�Xy,              ���B0###100���Y�%�ׯ�s!���իc���%L(���������mq���ć^�hɷ̻��]o��H��w>o�۷              �cccY�ehh(���g�/�<M�T
x>r�܊	���Y���5t(flb,ƛ��rr2��U.�c||���R4][��Y*ӕ�a�񕇾����x�^��ٻ��{���$!aH�L��xEq�Zg�׹(2*��[�Z��[](�hۧ�>�`U@E�Z��@���TGpDEP�B2<�y+<���$�|N���s����Y�`��w              ���KI���ˣ��t��E�i%��u��1���9����� @�ŬX�"V��b�)Y�f�PL#��������|I�9fL䥚�_�              ��*++cٲe�t��())I?�l׌d4��ݻ�E�b ��5�kb�������c�>��T               ���"JKKcɒ%�|��Q�ŋ��K����2�{�4� ��]��[O�U$            �dG�tDL�35 ��Z�re:�RRR�~��v�\VVДu��!z��4� �0�0�?���d             ��ާĻ_�o/x;2Mn*7�=���a�F�_� h����cɒ%�|��X�lY: ����~hΎ8����
�P tT������o            @ӰK�]⮳�Q�����12E���1q��8�ǁQ��,  SUWWGii���K�)))I��-UϞ=c�]w�P �jת]���_�y��W������q��������            `��s��o��v8(ν��(YYҨ��=N����� 4����t�e�����$��_/^��$��``݊���SN	�P 딜��}��ѳc�:Ϳ�����Ϗ�e            �,��yZ��u�8a`�6�?~��Vq���Ņ] �PV�^%%%��K2j�k��@Luuu �өS�8묳�u��A���[
rb�Q�㧇�4���78I����ńY            �\�:���/|>F=2*n|��=�!�b�n{ lN����	�|���+�|R�T���';�����P k��q�w�O��ţ�<��w^�[6/            �̗��7�xC|���9��I�HzK�gH�|��ѶU� ��*--]~��L2V�^��ӦM�h߾}l��V��v�E�^����(h<B1 �O�\q�q��/�Tvj��KV��������            ��9y��c�m��3�<#^��;~AnA��_Ņ] P����X�d�ڑ�_�8L2.\(�]�vѩS�t���8��������E(��ۿ��q�w�.�w���'�{"ν�����             ����o3Ο������]TWWo�u{w��O�]�������� �Seee,[�,�/_�~�	�,^�8�]RRUUUlY999�LM��1�Ν;���t���B�r㗇�2.;�He�68��e�ӿ�4���6�	            `˙����wX��ԫ�9y������О�ƈI#b�śt̑�G��+�-X＊�����+��i� MSEEE�����/I�%��$�k�K^�&FAA���K2�L������
���hϮ{Ƹ3���������s��9�Ή�K�            �4�5���{C߸��[�}�Z��w?1^��8��3�ُ����ڵj8�q�>gnp�g%�Š;��= d����X�|y:�R�I0�H�K�	�@�H�RQXX��$�$�R��رc���-�P@���?��Ob�1cҥ�Y�fE�yrL\���QU]            @�R��4�=8���d�|���&�M�s�+�.�:���f�51fʘ:_S��6�Ƥ!��gǞ������{�Ǣ��ƕ�`j�/5A���If�ʕ4����t��s����$�Daj�����b Z�=��#Ɲ9.}ҥ.����8���c��9            4m�g���?}9&�����u^r���G���v8(��_:�ֹ���ta�=nl��i���WTU�;@�ƫ���+V|+��t����d,\�0V�^@�*((H�_j�7c0ɀ�h�3?��O�ʣ���ɖD�����+����w�            ��w���n���q�J^�����.y-�LSfO������������:}���d�'q�g��< lk#0˗/�e˖�C0�/N�WRRUU����J����0}I0I�&ӱc�����B1 �خ]v��g���������D�������            @��h���^3?�7�rs�mնֹ]�u���},��zu\5�����L�߯{��g�=��V;l�xy�/qΤsbI�� ���I�/I&y]�^򺺺:��WPP�6���$�Daj�������f�?�G�"1++V�O\����'k            ��k¬	��ܗbҐI�W��j���N��F���rp�8$N�����#7�����k�F=2*n|�� ��������˗ǲe����u2j�0@�Ib0�:u�Ν;��/5Q�$����X�b Z�7�x#�M��{-            ��㽯ދn: n<��8o���;�О�Ƈ��a��6��_�'L_��RՄ`jF�I�/���E�bժU4����h׮����7c0I&����3Z�Օ���WǵӮ����hJ�v�]����L            `㕯)�������}<���?GqAq�s���0kB�����|�� h	�����s��MG`JJJbٲeQYY@�j۶��LM&�NF�6m�"�����oư����_��"9�t��Gǐ>C���'Ǥ�&	�            �f��?L_ot��{b������Ip�?'�g��?@KPQQӧO�_|1�4�T*�����K��7�sss������"~3�71��ѱ�bU4�u�-������v            `��x�������]�x��#++�N�{{��1p����Z���Ҙ8qb̛7/�-+???ڷo��$�5#y]TTT��@s!�B$'[ξ��x�ӗ#����A:3�ǀ             Fr���oN�a}�EQ~��/Z�(���1�t~ �"1��|+S\\��0��	� 4sU�Uq닷�œ/�kVD���ʎ�z��Ü���:�u             '���ˏ�<.;��v]th�!^���8��3㹏�����z���Y}�f �f$����kh��|5'�����'Xzv�g�=;��7,�-�6            ��׹m�sНqd�#������c��3⚩�Ę)c�7�h�>����?��w|+�R\\�6
�lgee��Zv(����UW�}z=�[F�;�[����!2Q~N~���	1���8����a            ���OGb�n��F������v��J@s3e�׹�b%���/��f&���ly-:S��$�.�[��I�
h\K�,��s����H-8��g�>�8̙���Z�            ��$q����*~~��7x3�E+Ōf�)�OY�#v:"f���t�x�����X�`A|��g�YNNN�k�.~���Ԅ`:w��4.�B ��n��bH�!1���ع�Λ�^�겘����[            �8�mO��v8h�s_��R�q������
�|��ѶU���=�G���W�US��ʪ� h��|�̀�m۶k�/I&5��}@f�`��K���;�>�s�'En*w��KN�0��?s|L|ub��*            `����q�wD���;���:nz�����KcM��{fM����L����]�gS٩}��8�_��w�y��@S�駟4�T*
׆`���׆`:t��Z�
���`�٭�n1�������ܶ�&������q�q3�����            l��윸����#/�����]X�0�N����w���jv�b��c�.\�:��<4^��z��x�������/2E~~���KM&yNFQQQdee�<��P�/D�׏�ZQ�"�~� ���QRQM٪��IQ~Q�{`:3�ǀM^���Ǥ�'ş_�s�Y8'            �M׽�{L<1�q����`F�u�Y�y���YY�2.��E���Oş�9���un�����s����).}��XS�& �����X��y]J�+((X�IFM�f[Z���]9�^�Tu	�q}Z�i|Z�iи�ZprBhH�!1���h��z�֛�l^����q���ų?���            l'�~b�6�ت�V띗\�Sߘ�_��K���+���P��b��0�w�g�yF|��� h*V�\�����|+S���~��O �l�;�������튷�,k���Mq�CGeUe             �O��Vq���ŏ�8jY���C&�'�{����d�'q��98.;Ⲹ����7��M�����K^�s�=7}�i�� 	i��(((�V����xm&����� �L(����ɏv?!F���<|���s~�|�            �.��Eq�Anp޴9�⬻ϊ�6�XUqœW�+����=�j�U�s����!��O���+W 4Uߌ�t��)=��$��� ��P �t`�c�~��{� 
�7i��K�F�T��ҮK             #'{���&7��rʕq��k���j���}~�O�=���c@��Z_|�ű��c��> [NNN�k�nm�����[a���� h(B1 ��u��c��cD��g�=7i��5���fM�G�}4�8�	�            �_.�2�=8�̞���Nn<}�͇�eG\�yydge�:w�n{ 4������d$1�$
S��� 2�P@��Nš;#�����8)rS_-L����|��9>&�:1JW�            �Y�͙����/��ŎQQUW<yE<���q�;�7��ƒJ����0~I0I��&
ӡC�hժU 4B1 -Ԯ]v�a}�����G綝7i���z/�y��?k||���             2Oo�f�51fʘ�M�B���7{ńA�^G l)999Ѯ]��1�N�:�G򺨨(������hA��b��chߡ1�ǀMZki��x��c���1��iQ]]            @f���8��3㙏�i�c���8�O����Y\��D*; �1


�ᗚQ\\����lgee@s&��egeǁ=�!}���>��un�^���2�0=&̚��~�X�"            ��6u��|��XP��ѾCr�����s_��Ϻ;�v��j��[GѪ�z}�C���R�(,,L�_� L���t��1����%�h�����{���^�}��y��Wc��q1�Չ�z/            ���T��+��2�LU�U�	f|0#���^1�qq��FK�ey�辬~�|�)�梠�`m�%I&���lgee �&Ќ}�_��ё�/�}��q_�{y\���+            4-7<}C:�i�-��o;>~v�����" 2]vvvPwI襨�(~�	�Ԍ�u~~~ �q�b XkUŪ�2{J��5>���_3�$            P7�|}Puuu��>6��?- 2]AAA:~���������ڵ[)..^��ԩS��� ��P 1�Y1aք�땻�5^            ��0�ә�鲳��u��QVV-I�6m����7��H O(��Jj�����ƭ/��/|?              X��ݻ�;��I*�����h߾�� L���:D�V���"�B�r���
�����c��Ӣ��:              ���={6�PL{���$1�dԼ.**���� ���h���cH�!���W��=���g��}              �?�{���S�Fyyyd������d��$�YYY@� @�Νv��G��ˏ�<����?s|L|ub��*             ��,///���4����t�%	�$��LM&�@��O| �%;+;��7�tc<���1aքx��Ǣ��"              Z�$3{��;w�f_���`m�& S3
#+++ �E�b���{�u��u��o�}h\{����M�C��UU��X������^��}���/������uzz�[6/��������y�             @K��Zw�uW|����lQQ����?�`�P lH�����ؽh�:�ߺSݣ2���O�}��'DS��',S��$����c�.�ư��b�~ãs���^�[a������o�������o�/�              -A~~~�}����K/ŋ/�K�.]�/''�[�d��uqqq�R� �MѢC1 -�;މQ���_>��8t�Ccd��q�'En*��k��e���q��k�������t�f�cu��              hΒ���˖-����t$�]�v [�P@SYUS�LM���m�#���=��Y�R٩8b�#�ci�Ҹ��{c¬	����Fuuu             �ka��١gtl�1rR9��bu|��˘���X�bQ�|�����K��;ﯪXC&	�����0 ��� �`�K�ǍOߘ}��#���3�93ڵ�����8��d���1�I1n��h�G            l9YYYq莇Ɛ>C��^G�6E��:w��91e���s֝��'�7�wܮx�8}�ӿ�~�겈�  �A��,\�0�YX���[��q����u��f�����D�>�?���q�C��i{�#�������I��ڥ�.1���q���������Y� �             ��눝���Ǐ�}�ٷN�w�Sz���1�әq�ԫ⡷
   ��PL�� �-)���9.=�J�}ſ���c��^+;+;����             6��T^���w��m�͢}����O�)���^s�	   s��P ����Oc���q�S��a=��}�Ʃ{��s[            �8�䵉�G<��<t��wd�#㕋_��rA��9>  ��$�UUW��9S����Ǡ}ň~#b�n{o���:U1�Չ�0            P��Tn<x���-S�m��1�qqx�����嫖  �Y�b ��E+�M�ܔ�o�{�3$F�7":��Q���a�{�ظ��k��O���^�/�~���j�W            |ۯ��U��-��оC������;N���  @��`��5���Ȩ����ɥ$sr�#'���dgeǀ��7'�&�0=&̚��@��.            h��������qzu�3Ο��阘�٬   2�P �lUŪx��ӣ[a�t0���ύ�{n�z��T���q˩��#o?���<��cQQU            ��$7j���"++k�󪪫��O����z(}���DUUUl]�u�;qܮ�������:�t�i�>-������G�  ���b ج�-�c��M�>�����GƠ}E�Vm7j�ֹ����NO�E+�o<���<��Q]]            ���穱��{�w�s?�9�?��O_����#}�Ѹz�ձ[��b�a�b���)�/���{<N��xr��  4.� ��Y�͊��ø��Kc��c�~���n�zZwH�g�q�s����            �����w��_�s�Z�ʪ������c�ġq�K��N�C��ԫֹm���C#�3�<#���_  h<B1 lq��J��oM��;�g�sf�7<�w��5�            Z���o�8����f����;/�����S<{�f�}�����?����u�k��*�z_�4<�ug   �C(���W��O^c����z#����81�Ry            |ױ�[k����^P�HL��+���"^���wƸh۪�:��d����kx�  4<� EUuUL�35=�����:=~t��b�n{            ��%7l�ͨGGE��M>ƃ�x0�_�~L>9zl�c�s����SnI�4��gn
  �a	� �薔/�?�����}��cH�!q���F��            Z��n���W������f;�_��~�/�r�_b@�뜓��7�xc�r�3~  @�� ��5���Ȩ�������-����˿F*;            ��$A���/��7���QU]�Y������?��O��w:|�s�X�oN�M���W�U   C(����bU���}�mѶq־g���#k=�            �Q��������}3>��E�Y��,���������]��u޵�^��Ō�2&  �-O(���Y�g1v�ظ�����Ɛ>C            Z�$S��_��b�]Y�2N���8xb����Z�]y���&�M����  �e	� �dTUW�3=��U�           �9).(�uߢ�E[�ث+W�&� nx�zo���C��T\��  l9B1 4II4            ��6ymjݷ�b�?~eUe�4<�|�~g�:�'��I�d���]���  l~B1 d���!�j��w�_�bq|���            ��l٪e���ئc�]:w��$3��Q��4~|Џk�w��.��܂��?r�h  ��b �hWsU���Y�y��W��w            hΖ�XR�Nm;5H(&Q]]M�(*�*��/�u���##������� ��L(              C-)�=ӹm�hHI,撇.�U�b�a�j�wN�s"';'ι�����  `��             �P�W,N��Zo��}������}����/�E��)�+����9����Tn�8,*�*  �tB1              ��y�ǡ=����pP\7��hc���kV���__�A���T^�kP   �N(              ��6�ZC1�Y�QU]���O�:}�_�����Z���<-
r���	  `��              d�$�.��G﮽��y�Gc���FEeE�p���b�����w�}  �4B1              lڜiQ]]�����6j(&�g~�k�����>����9�ka�   6M�Ŭ\�2��YZ��:t�q����ҥu��f��             ���K>�7�����ξ�}���_�U�ј��⟢���N�C��  `Ӵ�P̪����G]���и�PLII��I(            ����{|���m����z���X4�[_�5V�^����T   �W��              4I槇�t����wNF�bw�zw:s����bj�E�/�,��^��ئc  �P             @���������ئh���;i��b�λĻ_��`¬	��bU�u�]���R��e�/ӣ>�
�� �yj���^S�&*�+�<�*�*��U�U�Yu��f��             �QU]_��r�w���Sq����Yw������M�Ϻ;rS�  l����zb�����8���x�^����ʿ          MWY���   �玙w�3�����z���΂w"S����Q��<�@��i  ��iѡ             ����o�_�{v��;�R٩����c�]�"�<��#q�'ǃg?�9�  l<�             �&�����T�:�U��D���Xv�aѻk��쫨�  �n�b              ����e�<���?y>=  ��'                ��b                 2�P                @��                �pB1                 N(                 �	�                 d8�                �'                ��b                 2�P@3�K�]bۢm�)�Z�5               ���h�~|Џ���               �i�                �pB1                 N(                 õ�P̨]F�n���y�6]�	�q�nP��h�.x��(]S                uբC1�S��MN�:��O�и�Ry���f��                �ѢC1                 M�P@36��c㶗n��h��               -E�ŬX�"����<���4�5k���w������Xs��M               �ikѡ���(�.����+Wи�`SYY����!C1               @�ТC1                 M�P                @��                �pB1                 N(                 �	�                 d8�                �'@Z��n���ѻk��ѾG�o�>��I�+]U��ǋ?���/~�b,Z�(               ��!Ђ%!�����}�F�m�FVVV�>WYUO�t���1�Չ��ru                [�P@�a��wn\{ܵѡu�z>���Cv<$=�3&.y�x��               �2�b Z�����0hB���	�e���������m/�<xA��X               ��%Ђ$��'G>�����k��7"�-�6N��D�               �̄b Z�Tv*&��E"15��uT�6�tנ             ���m;ǀb����V�������ͧK�K�E�+���/|?  ��K(����ῌ�w>z���}Ό'�{"��            @�P\P��;'F��u�m���.�w�rW���ߧ� �M'���a����h��]��1��ɱ�|i             '?'?v�ctl�1r�sc٪e��|>Z�Q��\S������.�����h�צΟ�^�=~q�/⒃/��~�����/��5�  l<�� ��$'x6��E���=����ļ�y�hŢHe��C��}���О���;[��z��tj�)�?���_��W             [�6E�Ĉ~#��v���g�}�����+���_��oN�q3�����\7����a��!;��߭UN������rl���k�Z�n�ݢ�����L��  �b ���Zo����9I���.�{^�'���j��� J�3��?/F5:}��6� �N�U�            l~�q�1W���t�e}������s̘�n�uq��k��u�ҮKL9%zw�Y��]v����8��c�W��%�T�)�/�^��V  � 4s��>u�'yf|0#Nwj,Z��N�%'~nz�x�G���n]v[�n��ҥ�is�            �y�تG�m��b��w��g�Ryq���1;G���X�b��'�#=v�c�-S#��<~�������9&  �aB1 ��q�W�7���zl�X����~���8���ū�]��sNr�H(            6�m����/x:��)�n�7��d����b����>���g�}bK�a����!Nz  ���{������˵�Isk�
��B��r�# �P��eDgG8�Ł3�=��3�KE��((

3xA��P�S(��M���ٹ�$��~Wz�씴�ms�|��+����<OX������2B1 cXaAa;�؜��ޞ8��s�*3`m����_�]��S��9?�]�            �?�E�q�'���H̀Cv?$�;庸��Wg_��e^|�}_����ύS�95~���  �P���=�6U�sv۳��������{�w���'�șG���Q\X��L             ��ړ���]���]�~�۱�uu����{�X�9�-y(�\�d�k_�]�QV\��'ǾS���>1�������Ӿ"  [H(`K~�2��?����'�V�P̄�	1kҬxm�k            l�ݪw�+��2��-)*�O�����?��:?�9+�W���>n^x�;�b���8<���/��sN�$vs̬c�7	  `x�b ư�����ؽ1�Z�T����k9�V9M(            ���#.�TIj��m[�,�'}��X׾.:3�1�bJ̝67Θ{F6㰜_wּ�bEӊl4�o=���8��ψ�tӰ��'W<�������+�}%


r�w��  ��ê˪s�/\�0zz{�v�7[ތ����^5}��            0|Il�C.r�������7������y���>N�sr�t�M���z���]���?�k^Y�J�������zK}��_͆g�?�����������  �;��jR59�W�����V�����{             �神G��HB+���'㖅���u�{��8���C�=s��ٴ_TX��9e�u?q�'�*3 �ל���1���fS&N�y�̋V�  �;ס����x���a�_^^�����o�9��vD��q��.�ι��є�{5v4n��             �IsNr��'~8�H̀�F�g�'���l f(��v<������L|����mݖs~�G
�  �0��PL_���c����ع�簷w��툴C1�'��O���~��������T             �f�n�s�o�����-��ӫ��[��5.9��!���?�|��Ż���zR��A��v�/  ��ס             ���������_g#,[�gO�l����_�?�+����H�5�A��&�  ���              �`�*c��=r�������>�����{cT�V��l^6n�|yf�39C15��   �g\�b��<+
V����� v�e�ˢ��7F����             ��Tm�=�����n�/��.��f6h�ʺW"���^uYu   �3�C1��n���T�V�s-�[K2K            `��,�̹�����/ަk���圡��ts��P׫N	�  �p��P             �HW5�*�~{W{���lӵ�;s\Z�Z#�Z:[r�W�	�  �p	�              �`'L̹��ն��n��}�Ξ�ȧtO:�~q��� �p��3             �VXP�s�+ӵ�����}���~   #�P                �'03�����z����s����ǔ�S"ߞ]�l���m               �P�8t،òkG8a��+�n}�V�               ��                �N(                `��                �b                 F8�                �N(`��tS�E�7               �B1 c����.               `t�             �f�̈%W/٦kԖ��ܿ�K��}O�|)-.  `��              �B%E%1{���r���  F�               �B����aÆ����O�4)R�T ��"               ����O>�d<��c�����YYYY6S[[�i�������� ��5�C1Vu�u�>����`�ګb��c�1�=��H���              �KWWW���?��˗�wvvF}}}v�����������۠LIII ���P̹������]v�%���S�g�}f�fi�K���              �G���2�Nz{{���!�r�����I^WTT ��P               ��?˖-�n�okkˮ+V����f�1ɪ��y�q�
��O(             `[ټ2~��c,��t�h��d�G�i����5k�d��J"1���Q[[�)��.++ ��             �l��E�;> �</��b����������)��.]:h^QQ�)�րL򹲲2 =�u(���!{�}~�@`�������?�#Q�/              ����z�V7n̮7�|sЬ��8������l��L�2%JJJ��c\�b�2Z�����?��+y��ed)+.�y�̋�����Q^R}�}�a�Xָ,^]�jt�t             �H�+�2d2�hjjʮ�K��mVPP��՛�1IH��eee��5�C1 l�T��zI�2�8jϣ"U������xj�Sq�swĭ�����             ������M477g�o�1h�J�6�c�USS�)&�'� �K(���:�;�����ˣ��tX_��w��Gg�WN�J|���ė��r�u���y             F��������.�NgW}}��Yqq���1�z�q2`���'�8�[�n1�xB�YSGS4���z�#�8"n����Y;s��Q^RWU��������O�x2              v4��-��dbÆٕK*���I�[�2�qAAA 0�P�W\X/\�BԦjsΏ���xh�Cy��I{�����̆^�a֤Y����1ι������            �h��zU���l���U��X�N�����~Ь��8*++�ј�S�F]]ݦ�Luuu�x%0ƽw�{��ļ���xx��y��>S��_]�EbT�V�]�+N��	���'            `�ڐڐ][�+� �E&������Z�t��fEEEQUU���$񘚚��q�&O�&L��L(`�;}��C�n|�������}jR5q��ݓ��=�JRq�E�Ł���h�l              Ɨ���!#2�T*�)��$$�e�

`4��Θ{F��������[�v��O�>���;����3��o�����              ��J���U__?hV\\����hL�I�1A��S�f� #�S�a�V��M�/���go�tO:/�I1���a�ۜn�^{ �[�\4ll����V9-��6?N���(-*���_z��G���5              `82�L455e�ҥK�S�TL�2%�ykD&�ʔ���H 0���C��|�μ��+�}%J�J6{N�����M��]����Ԧj��]WՐ�K�2�9���3            �X��{��-��q1m⴨��������?��7[ތ��ǂeb��E �E:��+Vd��J"2�d%!�$ 3p\PP ;�P�v����߰qC�i��r�i���C|h��,oZ���i��ڗ7{^S�)���ڸ������C6���/�+�2ں�            ����uL|������yL�0qX_�F��~�]��h�h ���L����͊�����*�I�1I8f (SWW����/B1 cؑ{�s��E�D�/��{\x���
�P�=�8��������Z�ra|�G��?s�JR����N�{z����            l?�U�7�sS��ߙ[���&͊�O�>�x�q����1��� ƒ���hjjʮ�K���R�M�d%!�$(3eʔ����-!0��{��s�?���y�����f���{m����-��c���xC�A�$?X�           `<9|����圭jY�y�7y��������cw�����t�������k���iq�-�EKgK �&���[+�NgW}}���@D&	�|�TUUEAAA ��P�U���_�'�-|sa^��=�]r��p�{������C߈K��4v��}�콳�            0�|崯�I{��s��w�c^�u��c��KⲼ]��9'ǃ�=��t�X0����fc1}}}����LQQQ6�րLr������K`���fM��s���-�[��{$?�ٜ�.�ntf:���=q�S7�5']3h6�vf�R�K�i[            0�U�U�~��������^�{��䎼Fb��m~��_�i�~Z����hPPP�T*6n������FSSSv-]�t�| "3�8NVEEE c�P�5{�����?}��)Vn.����x��|�۞�-g(&1w�\�            ƅ���E�9gI$&���Cr����Ɣ�Sb{I�Y�x���� �Ŵi�r�:`gimmͮ�˗�Gee妈LMMML�:5�L����QXX��$0F�Z�k��5���l.��ʧbY�m�ǋk^�խ�cת��<s�̉_0            `�;}��s�'���;�~'o�����]����S��_<�Xټ2 F�3f�0jd2�hjjʮ��s[TT���$�$$3�^���0r	� �Q�*s�7t4���uu�w��C�\��������:qj            �xp��cr�/|sa��ᵼܣ&U����9�s_�x�����`ق�/���tf����>g�vT�U��e�e�{}�W���`�����~8`���������%�J�- SSS�)"���� �Q�9����y��!����#K�|yi�Kq�>�گ�P            0�M*�{M�+�����}�p�br��͞��}]��/�.~��׃fk����_��x�?b��)q�Y7�G�t�k]t�Eq�o���/�؞�M�ӧO������,�NgW�?륥��2�e���ؾ�b ƨ�	�C1I�7�q�f�O,"�%��Q.�*            ƺ��8<


rΒ(K>����f�y���8�{�Œ�%�x�����[/�W׿_:�K9�I���/�o?�� N:餸�[ƫ���X�vmv�J��ј)S�d�[�2eeel;��1���?���҉y�����Yָ,��֮֜�UeU            c�{�s��/�����r���u\̬�9�<ӗ��z��"1ou���^w�͇��P0j̞=;�͛/��R ����쪯�4+//[8�Ǖ��CF���Z:[r�WN�����qؐ��W=���՞s?_�,            0�͝:7��c���=.>������c��[u�+�2>8�1�|Ҡ�{g�7�>���� �:�hhh�5k�0|ٵjժA��������������������� �B1 cTK:w(fת]���3jf�nջ9f�3�OE�E9��2]            c��ɳs�/\�0o�8y��CΒ��|���n��:�k~-�v��͊���=�^{  F�$Xq�����+V�`����FSSSv-]��m��������d�1����T*0�� �Q͝�9����m���3����/o�%򩢴"�~kWk            �X7kҬ���zϻ&�k��X��E�ě-on�=n}�����_��A�Cv?D(U***�c�X,X� {����`��������Z�l٠yYY٠���quuu64c�P���}}����3�6UM馭�����r����-{,�i�ĩ9�[;�b            ۪ʪ���.���5/����>f��_<�m�Ǫ�U����|o�>S�	�Ѧ��(�=��8�#b�ҥ�|��hjj�����J��lI����>��V����l
��mP��Xr��g\����ꎍ�.%7�������n�s;������I���yg�-o��k`���=���h�l�|�Q3#�P            c����9�7vo�tO~"��:�����ro^�����s�bfO� �Մ	b�ܹ��V�L&��ڲ����hooϮ�8�knn���� �����hhhȮ\R�ԦpL����@L&9Nޗ#͸Ť�ұ�mðϟ<yr ;W����܎H};�6��Es�9jR5�fy�G�:3����=��?���ȷ���˚�            �e�9�;�v�#�8b��S+���������/�ܯM��XS\\�)>1{�� V�hmm;w6�<�IB2I`&9���	`�I���U__?h�<Õ���g8��$��x�ԩ��Daaa��0�C1 cY__<��#q�~g����ǡ3��+n�u/;���x�ȧ�8p�s��[            0��iJ7����N�w��#K�|Y�>����˪`�)**��J�H2�J�2I@f�u����`��d2����K��m�Db���Ed^���l/B1 c��^�]�PL_��Yߊ�w\d�2þތ�q��9O*���z_�Ӽ]���	sΆ��            �C�b
����w�E�ECΟ\�d�Ks�9�~eYe 0X*�ʮ�ӧ�'!���L�inn�F-���J^����_}}}CFd�s;�IV�I2���{�P�v��wƷ��v����{?8��_}jX�O�27�sS���yί��Ut�vG>���	9�:b��            cYg�3�~���U����Ο^�t�K[W[���	U���L�2%fϞ=h��d���$f��d��L���dOH��$┬���A���⨬��Fc�xL��$�rIII���P�/{~%�HN�=5.����<��h<��_�vg���ǎ��}]���q�A����OƤ�Iqٝ�Ś�5C^���:���3枱�����E������f�3            c]KgK��ʲ��b�qؐ�Ǝ�X޴<�;�{�J�J��,;ӗ	 �'	R(r�dz{{���cSLf ��Nֆ���;��IN��ҥK͓���s���S�F]]]6*SVV0�C1�}��|W�/�����]�]��}���Ǉ���(,(�9?{��ㄽN�;_�3�~��XҰ$ֶ������=iv�����#>uu��ςe��7���>�rZ�4礜���<            0�5��s�O.���%�I�e[�g�{����ͿD>���~ssg�S$`'(**�����>}z�s�����E{{�ۢ2�����9����,y�U__?h������l@fภ� ��u(`<xf�3q���}b�s�(L2��9����]�v���%�\�b            �
�$��e����?m��w��%f��r��P��҉9��:���)	S$k��L&���I�1�����{����� ���"2I����*�I�1I8f (SWW����� 0\yϕq��'Ō�����y�7�В��~݋�8�~�'O�|2            `��ؽ1��MQ��4;|�÷)sҜ�6;xi~����ܑ�֮� `t*..���={���[C2�����ښ��$Q�d���%����6����g*YK�.4O�O�j���L�x��!04v4�G~������GyIy^���eU|��OF���1��9g�-{,�2]            �������=��ށ��7��V_����r���Ă7D>�Q�G����O �Mo�%�No
\$+	�$q�dmذ!����6�s�����A��9����>�S�N����M����(,,F��q����y��w\rG�JRy�f�'�Ьk_�v�qW9��Ż            Ƌ�V>�3s،�bߩ��+�^��kVN����=m��3������ȧ�w�?��k^ ƯT*�]ӧO�9ooo��cZZZ6����^ggg [/��l
5-]��m��������Fc��sϘ;wnL�<9�y�b Ƒ߾��8���㗗�2���#�����q֏����)��L���ќ�������#            `�x�����|a�~AAA�p�q�����k~���gc1C���{#��~P���� e�ĉٵ���'���x�[?������`<��퍆���z������:(N>��(//v<��q��+�~����i_�O��(-*ݢ�OB-�={[\��bU˪��=^s�5QTX�s���ǣ��>            `�����cc�ƨ(�4;k�Yq�����1��U�U�U�_��s~���#����g��䜽�� ��UVV�]ӦM�9�d2o�$!��5�Ib�;���g�y&�-[\pAL�2%ر�b ơ�Ζ����!����㓇2�9�������,iX��z_|g�w�5/m��mﺽゃ/r~��w            �'I$����0����4��M��k�㵊��sn�ݫw�+�=�2��Q���9�`{*..�ɓ'g�P��t455mZ���ـLr���]]]�?ɳq�-�ĥ�^UUU��#0��l^�����\>9��u��5iV���g�b���x��X޴|�|OI���o9�����            �77>r㐡��������o��������͙2'�}����}N��~��'�og�;+�~[W[,Z�( `gJ�R�5}����7Fsss���FKKK�8	e$��JB30�$1��n�-�)((v� �:��%g�δ�}]v            ��S+��߼��8c�9��/���+���q߫��3�����k���*��1����gŅ�k�-oƏ����~���/:����o,�L_& `$���Ȯ�v�-�<��d�I<���1��۳+9N���L�XS__.��;,�1�b              F�+��8q����l�s&O������������ȧ$R��=s�^�s�5 �Cqqq���f��ٳ�{{{���%��h��~nmm͞��C=|p۟P             �(�x���+�;��v��S+��?��_��C/r���
 뒀ƤI��k(�t:�������=���6�nll������ _6n��/����/���b              F��.�n����|&��m�h������ۓ��V�UŹ��s֜n��i ��T*�]ӧO�9OB2�����Ғ�sGGG�βh�"��D(             `��]����~|�=����ںڲ��e��"�>���GuYu��=���{� ƪ��̮��s��d���-������=Z[[������^�����V�X�B1              �Ho_o\v�e�\�s�3��[}�$s��=3^\�b�[UYU�ӱ�4�����  ?������6�r���͆d�xL��Ǽu%��I����3���b����/�L(             `���ߏ߽����/����ams�9���oƷ�V�v�n�������T>)笭�-��� �EEEQSS�]CI��ـL���۳a��׍���e�ƍB1;�P             �(��iy|��O�U��*>��ǉ{���~H̨������խ��%�����^��l,f{I����}"��M9�w�xwtf�� F�T*�]ӧO�9OB2---���ܜ]���$��5�BB�1�	�              �r����w|7�e�eQUV�������;��I��c�� `����.9�L&��ڢ��)��ۣ��5�ill��%1���� �޸�|�]��9Us�}������u�ng�������?bcF            �~:3����  ;Jqqq���f�P��t63����@\fÆ������u(fZٴ�=���ϯ+�`�)�٢�v$*.���              ƩT*�]ӧO�9�$����hnn��I�2ɂ�L� `��������ڻ�c]��               Ɔ���P2�L6��c�!���L��������b ư�O�>.?���n}�ָ��              0>Gmmmv͞={м��7Z[[���=�y �De��Lr���0Z��PLWOWtww���,�\�s�%��H���               �WQQѦ��P��t�����Օ=NV�I�2�}��u(�uck$�USS�Ε�G5)��fB1               ;G*��+V�m���2�M����QRR���===و̆�!�丽�=;��a\�b                ߒ LKKKv��^{�uuu1{��(**ʮ���������l4&��$_�~��lL���YH��F(                ���_2�Lv(((�����>}z��~ِLqqq���Fwww���l@�7ވU�Ve�4�-�b                `�mL&	ɔ���̙3�+���7n̮������_|1��0B1              ����:c�����:�  F�	&dפI�6�-Z�(z{{�C(`�џ-y(ƢM+            ƃ��c�n�c$��tEGOG�������cm���������0�����k  @(`{z���            �^��84����2}�Xټ2��.��6x�xb��}   ��b              �*Ņ�1kҬ�:{���S���ts���m�����˛	   ?�b              ț�TM|�=�ͮ߾�۸�w�ĳ��  �m�b              �.N�{z���)q�o���_���'  ��#             �vS\Xמtm��Qq���Ds�9  �-'             �vw�^'ă�=�}�h�l	  "������7`8�b              �!�~P�������L  �wS�N��+W�P             ��p��8�'�HP[^�Q^Ruu1w�ܘ7m^�3u�(-*�5�������k�?\  ��ĉ�K(             `k�h��_�?F����8�]��G�4>����&U���9隸�����/ �xV^^0\B1              l��ޞ�������;/�ˏ�<�t򗢪�*��Ņ���ӿg���  �
�K(             ����tƿ>��q�w�ݟ�;�����}p�Ɯ)s����  �΄b �ٓgg(�G��{��1�jzL(�5��(,(����H>�:��+��ZWŪ�U��iE<���x��             Ƈ��D��t|,�����}�

�3G~&���   ޙP CJj����8e�)q،òA�mєn��V>�_������+^��z             cWcGc�s�9����Ң�A�s<G(  �I(���8ab\t�Eq�Q�����kצj�љd��3�O<W�\|��ŭO��7            0�,Z�(���w������ڙ1o�y�Қ�  �<� �&O�<������T��继�;~p��3n��>�ո����;            ���[�|+�p����p�쨙G	�  �0� ��u|��y�����r��Tm|�_�O���W��CK
            `�Xټ2��.��6�,�  0�P�8VPP����g~#�w����+���������r߿D__             c�_�c�(�>S�	  ����*  ;EQaQ���?����I���K�|)�Ý�~qd�2            �~���h\�+��^�{   �L(`*((���q�!�Hu�A�G\�󋢯�/            ��mu����*�  �΄b ơkN�f�"1K��ӫ��V�˚�Ś�5���m]m���d�)),��&Ɣ�Sb��i1kҬ�������o����h��������s             �[�^�\�K�  xg�:���6d}2��'�s�������nG���{�S�ןz���l�c�ӿ�4~����F��t�$s�>��E�\G�y���暓��'V<�}��            �^s�bJ�J���x�/�  rס��޾�����������-y����܎H;1��ux����p����������w}��楼�?	�|���g�~���>���w����'�����ܯύ���             F�$3����   6o\�b ƛ�O�:f����9K���~�X�l�v�^�]�����柾7���g�>C��{��q͉��տ�:            ��ir���]�.�  ��q���.���/n��{_�7���y���;ʟW�9�׃��o���?{�������1ִ�	            `�����s��{ǽ�	  F�q�y��h.h��e�e�\k���b��1������^~��Q^R>�����#�ӻ㿿���8��s���q\|��9ϙP<!��迏k�6            ��g��Y9��[�  xg�:�x��[t~o�7���ޗ�-SZT�;�sC�����q��H̀޾���/?�{�%g]|�73{�lvs�$�%\BJ�R.���@Т�
U+ڣ�ZK{<mEO߾�}{U(��K�*o+r{=h[���P�\� �����wf�}�ξ`f�&l��3�Ϝ������>τ���r�|w��e�C�V�O�����[����            �.'/?����=�  ���:P/N;��X2wIŽ�сR$��+#��8������>�v�_4gQ��u���            ��rʊS*��ݴ6  �W'P���'�����Y<����z7���~q��9�Pq�G}@(            f�c�;&�/Z^q��  ��b j\:���W�]qoKߖ�l�eQm��������Q�����z�Yєi���H             �ß��O*��Ÿ뙻  xuB1 5�}���sVܻ�Ǘ���@T�$��;�_zϗv؛�<7�����{��            T�3^F����W�{d�#�|��  �:��w��*�'��k�6���y���_��Wјi�a��U(            f�7t�!�q�7&�����-  ����qo:�M��{�xf�3Q�^̽w<sG������r�[�o�o            @�z���U��,�.��?<6_��  L�P@�[չ������~T�۟��b(��            P�������;>�un�R�I���+K�p  ����N�ce�ʊ{w>sgT�;������Eˣ)�#��             fVkSk�~�����N���I����������
 �zW(�J(��-��,��ي{k7��j�<�b��C5�!�+���7?            P�^xp�{Թ3�4J��z^v^�5��ܦ��p��R &y~�ޮ��M��s/ @�
�*������+�o��z7E�������لb            ��.>4����;jŕ�\�x� @���@�T	� ԰��Ί����l1Y(fi��             f���)~��	  ~a۶mS%PÖ�]Rq}S輦-&{�K�
�            �lrُ.������B>  ���������a��,���R�K1[l�m������            �./�^�߹�w�Go  `�	� ԰����냣�1[L�\'��            աw�7.����;�.��  xm�b jXSCS����p��c��ksCs             �e4??Z�����k�3���  �B1 5�)S9�/�c�-�V\oih	            `f�s�5���<�u?��p<��X����{l�c��?ۥ���v�o��  �oB1 5�1�Xq�X,�l7ٟ            j�mO���0�A�H��G�ݗO�#����h  @]�bj=(��v�x`f�ӲOt���짽?�|q�~�            ��h~4��  �ou���bռUS>���3��uz��z���.����	               �O�X����(�a��:                �%�N����|���D___lݺ5�l�2���r1��                ؉$ ��dJ��I�/I&��ݱiӦ����a��               �n�R�hii����hnn.�`��Klٲ%�n�Z
���00S�:ӝ뎞��T���0���g��j�/�              ��/���ҥK#�����XEwwwlܸ1�o�^zժ�C1�c�1:::��80�
��.�n�QR�              `z%񗁁���닮���H"0��d���K1220[�u(�^���q�!'�l�O�>              ��`z{{K�\.W�'!��۷��zzz�P(�*��:��mii               T�������+E_��K�I�ג��b1�^	�                ��F.�+�_�!�$ ��r��P                �Y�)�_�A���m۶���p �O(               ������Kwww�����/�}2�k�1��#               P����J!�$ ��墷���پ}�D�P(T���5�����                Ը��`��K�I�ג��b1`w̙3'jA*��G��a��P|�oE-�wý              �B)����[�/��������l���D-�`�\u�U�              �nI襫��4r�\���M<޶m[̄8 	�{�P               �����Kww����陸OFrT��+W{�P               �466V
�tuuE.�����Rf���$S(f����8�#��C(               �5*�^��K2������Ԣ�;.�����C(               `'��K|��흈���0�}��z���'�|r���                umpp0���&F.������|۶m1<<���N��}�{_477{�P               P���|���Fwww��������H��&�Ĝ}�ٱ|��`��               f������Ꚉ���0�����b1�׮��-�����!��}B1               @����$������9�L&���8����㏏���`f�                3fpp0���"��Eooo) �<NF___i {VCCC���łb��x���Hϛ7/��t0�b               �=��)�$��_���m�bxx8�=/�͖�/�1��R�<O�RAu�               vK>�������K2���c���d>::����d����~I0I�����舦��`v�               *����r�������0�b1��#��N�_���`�(Ly�J���%P�>����5�]{7F=;zߣ��e�Ǖ�\              ���!�$���_���5!���1�ŋ�F9
�aZZZ��%P�>t���S/��_�����E��D=Y6Y|�����~�cq��
�              ukpp�|��r���[
�$��#������hkk���̟?"�dɒ�>T�o@���8'���A|��/ƕw_�Q��m�7>���ƅo�0��             �֕C0�a���J�^z)FFF�����D�%I&��T*`W�u(ftd4RS�&0��oDj;v2��]_~ϗ��~>.���q�Kc����%-<(.:���~;���              ��|����r�%��ݱ}���Z2`��d2���^
�$�$�R��tttDSSS�t��P�@�@l�MU��fVR0ܺu�۪T���v�vğ��OKA�����+?�J<�환��t����o�t�{Թ�Ig             `6���$��������0�b1�����P
�,Y��t��`��Dy�J����� ԣ������>x��mO�W�}E����1��������ѿ���8zߣ             �Z�<��_��K2O֒!3/�͖�/���L2��� Ԡ�}�sq�{/�e�MzL:��SW�Z��6���^7<zC���]�/䣚�i�g���x���իV�O�}����uI              �)�\.�{�R ����IF2
`f544��/I����d>o޼�>���Ԡ��)������}!.:�h�4���ζ���[>U/�^�������w�g���	���?޾�����q��gN9��6��˹Ɜ�P,             �t[�n]�z뭥H0�Z[['�/�L�q[[[@���P̷G�M�SuZ������9��kc6(����������K�{I���wN���]�x�'J#��<�����S?����I<��xz���_inh�UKWő�'|b�|��qȢCv�<c�����������             �n�b1�����ޑN�c޼y����"���P�:�]�ޣ��/W�E�����/�<N���8e�)��g�y�p�	S��t*��wLi������n�il��{7�=/��ͱ}`{)"�=�]�O��!�m�mєi��sƾ���~���e���G���+�!��oI�T�?z}|�?�Ol}"              ��[n�%x�� �Wss�+�/�(?N"1I,�]]�b ��mO�o��q��S�W�u��ѻu�9�s��eǗF5��� ��;<�*             `Ϻ��{Eb`7�R�hkk{E�<OFkkk ;'Pg��ʱ_:6NYqJ|����Y���M�X������[�w��;              �������~��2�L���O�`�ϟ?���舦�� v�P@JB+I0&�-;.��?����h�4F5��+�2�~��ǆ�             ���v�m122P���D&�L2okk�T*��!P����8����wo����Q���x�Ao�j�Dmn{���_��!�G�             `o��{,�^�c0�dɒ���(�`ZZZ�B1 �tv�w_Q�:W���`����_��W�z�o$?k�]���w�����ػ1              fJ��MMM��$����O�g2� ��P ;x|������|it�uƻ^��8����W��j��X1��+��c�����I����>uk�s             P֭[0�d��W�`�!��<�J0�� �S��6�5�]S��q��������C:�X�? ��wz���Xߵ>�m_��œ[�����?��p�             @5z��M&�)_�!�r�<����-B1 쒮���ޓ�+�_���--1/;/���͏���p�����@i             0��r������mmm�dɒX�xq)S�̛7/��t �C(�i�?�_��             @-�����=!�J�B0I���I���l6 eB1   P�F�����   �UŦb        �����^�L&�����������舦�� �
�   �QC��            {V6����$#��$Q��<�J�k%               �*���b��ť L)Ga��---��	�                u�����)�_^�Y�dIi`&�W               ��lv"���$�Da��T* �J(               �	�L&���K�$ ��_�Q����hjj
��J(               �5���D�%I&��T* j�P               PU&��,^�8�����u(�#~$V�]1��W,�������zK�f��?���`              @�jhh(_�L�IB0�(L�ill ^��C1��=$�w���������v���5���b              f�T*����R��y�<�� �k�:               ;���\������2�L���ǂ&0�<�-*��`��               �$�H̜9s���?�QKKK) ��`��d��$�N�����C1�c�1666����| 3+y���C-             `6��쌧�~:jU6����$��a�d��r �yu���uGw�{��'53`fEw��_��(_�             �M>��Y�ihhxE��)�d���_k               ؉��:*n������Q����+�/��ϟ�$�T* �nB1               �mmmq�G��?<c�!�NG{{{)�R�$#�'!���� ��	�               ��8���㩧��\.�Ǯ���P�Ҽ< S�,Y���@��.                �"���?����7�����}�$�`�L9S���� LF(               �`����.� n��X�~}�c2�L)��`��� L2/���� ��!               S�x����G?�7o�6���h̙3g"3o޼H�R �M(               vQgggi ��"                P�b                 ��P                @��                �rB1                 UN(                ��	�                 T9�                �*'                P�b                 ��P                @��                �rB1                 UN(                ��	�                 T9���{o��X�juԢ�������"               �� ԰Ö��<5jі�-               �B(                ���u(&ד�-�-S>���=�����[�L�u[��               �K�:�����Д�	`f�������_�UI(               �Eu�                ��b                 �\]�b67E!U����o����m��fc㷽������=���               �zQס��|����?�3�������\����                f���                 �B1                @MH�RQ,+���̈́b                ���������c6�                jB{{{G�P�a��av�Vf��                ��p*���_^lll�d�lْllhh(,Z�h���}��NX(���	�                 ���Yg���QG�b                 ��P                0�
��/}�K�]��T*U�/444������L&������;���n��'>1UH(                �y�b�|�i�&c��X>>�1>~?�����񥆆��������yST	�                �q�|>5>�Oߕ���u�e��477��3gΟ������s�`�H��q�>G�qˎ�%s�Ģ9�bn��͏�������gc����E��               �i���M�㔁��{���u��������ߙx.B1 �Q��8%~�����<5:Z;^��ޡ޸�����{��5Ϯ	               �i�B!��������zfΜ9g�w�y���� �q�����s.���]�������q.��?����M��'�>             �t:]�T*  f�$ʒ�������[>00���k���o��o��޺�P@x�o��Ms+�=����нaZ��D^��D�1���sڡ�Ń�`\xÅ�/��K             05�������L&  f�$3<<CCC�8K���󩮮����ꪓ����|����k
� Ը9�s��o������7�#���i�ޅo�0.��˧�.�<�k~��X�]_���            ���v͝;7 `6K�ӑ�f���)r�\f�j���w��������j��?���{�ZB1 5�+�Q1������͏M۵N;������N[$�,9�ߝ�w�B��G�             T& ԚL&mmm����b1����P���}��_=��h����P@�;��gN�w�]�N�u�/Z���7�!�g�Z�X�U�*��po��Z             �RKK�H P���t���F.��j544�p���rO]��C1��G6�ݥす��qA�e�b6{n�(�ީ�%q�3��yv��q��n��k�ՙ�bOjoi��~�X�ϫ            �WJB1  ������)
Q����V\}�՗|�c�̞8]�b>��ӱjު)�����z�~�տ2�#!�wA���k-_�<���Ž}�_#_�O�u�z�[�}G�oJ��d�O�;?�N<���ֿ-2�L�ӾO����>+;vG;��J�[��             �J� �e���1<<լ���S7�x��<�s�M���:P�N8��I�n\{�]�����-?�o�0�x�����z�[q�_\
�\�k�Eg��q��N�H(            �eDb �z��d�����tWW�WƧ��s� ԰��Y�}]<��r�C'|�N����YW�]�]�z��!�z殸�w��V�W�]
�l��               PM���W��Ը�t�W(���p@�P�͏��o*�r����s�t?����s��){1�b����~��Xڶt���tC)s��W             �B!  j�l��gxx���k�}�����<o]�bzr=ћ������̬����������v�UKWU\_��i9��б��1���3��o�.�{C���ܿ.�>���g��L�            ��666V��;���  ������|����l6��P(�7��1~��*244��!3}F�Fbddd��'� 3+�����%?h�K�.���s+������r�7t�!��_6���Mk��G����_s�5q�I�����|ЛK��bo��            �v�/k�f� P��HL�(K�R����'�I��b1u�W��N�?><<|����1�FFF���s�u(��-_�������Xߵ~Z�q��'�t��_�ba�ϟ|m������^GkG��xv��            �/B1MMM��d �����t?�J����#����}|�{����J
;~�=9g2~��c4�ו�{���������.8���b�� Ԩ�\q��M�N�5NZ~Ҥ{��Ѹ���_�5�{����:yc�a�%�	�             �����}}}���& Ԍ��8/����|�#W}�������ȵ��{A�<��866V��v2���7��B1 5j��%׷�o��k�,s�3wƶ�m���u?W��,_�|���V             �_�P�����f����\�x �Ile``��=ή:�3����555�c����Ò�J#��ښ�-��k� Ԩ��s+�o������}���t��g��v�ڊ��E��            �W*��T�>��N�c �Y#�^&	Ì����Ź�;x��7?0>}G̀���t�O(�F�6�V\�잖����;ݿ�;c��t�O�=�޳�z{s{             Ժ��P�yqMP_2�L�츝F~�����'f�����6�- �=o�x���t��]v��T*������H(f��+��|B1 5j�PL�����'?\N&_������e������-B1            @��銿��_�eava<v�c;=fӦM�q�Ƙ~����Ԫ����Q����^���<�P@���>�i��e�O����'��?�K�p_����               �ɤ�駊��L]~�뮻���s��i P�z�z*������J*��c�?v���^x(��dљ����              �6���=��df������e��OO�Ʉb j�d��������%���sN�����tj�4W\�,                ��n���)�O�3�
� v�{����:���}�'�t�C1s��T\��               ��������o�y��t�L\?�N8]���Q�z7U\�l������<���>e�)���Ž��O�>�{�z               ^E��	�
���\B1 5��-�O�w��ĥk.ݭ�fҙx���=��=��)�b���+��uv               �L*��T,���k�O׹�b jԦ�M��wc�۾�{�s�n�b�v�ۢ��c��;��3���K������               v�P(lJ�R3u���u"���ç���y;��p�	q����ۏ{�����|j���{�{1��2M��sUŽ����               �W�=�מ3]'��a��������߮�۸�;�{p��g��wL�>|�����Ǐ��(��qˎ+�b~Y�X�'�>               �3�t�?���i��	� ԰o?����bn���Vt��o_��8���cpt�U����W��ՑIg&=�_�ט�7�SV�Rq}c����               ؙb��?���������?����{o����'|b<xу���>?Z��I�s�>G��>��8zߣ'=&	�|����t;��*���ܽ            ��c�ރ���D�  �*D\jAQD�hA�^�`��n���[w�;���ә�gw��O�Ut��p��#��h�(JѕZQ��E֘r!�<�sH�ےh~O~��o~�����.O2��� �'�d2���-@����M�dƒ�[Է��	b�_�����M<���QY]��vEYIY�:.�~fn�w�y�+��c�����iצn}���3�����3o=               �	2�̝G���v׍�b z���[㟞�������c�M=vj�y(��lܰ��nW�vu�s�z�W               ���K/}�����	� ��?>��q�c���������iצn�g&��ŧ.nw�vomlܱ1                -�b R`_v_,\�0����b��Q�z�ׯ�>�۹�΍1Cƴ;��[OE.�               H���x��8�����%���A����־�/�<�Z���}{�;�{�Շ               �D( E6��g�rfܳ�8w���u�u[����̏��ދ�6k̬������5�4���V               ��P@��س#�.�v������:�K׿_�~|����mkn����O�[߫#On~2v7�               H�T�b��l�߿���[ZZ8���oi_>���_�;��_�ta,8yA�3���1Սձ����7~�m�/��?�w��'3���p~�++               �&ա�����Q�������8�v��;vt~�&R.�%����X��j@�3xL���G&��?������5.s$lؾ!�|gH��{��               �M�C1 ��=M{╝��whjij;              ���                 $�P                @¥:�D�����Y�fύk�ѳ!�!�ny;
����                �T�b�˾ץ�s8����Q��               �4Iu(               ��Z�"��G&�	 �VB1               	Ӹ�1�ox?*�* ��P              @���}�_ @+� ��~C�؁�Fi��X:0z���|>r�\�6�F���رgGT7V             �u��xk,>yq�?8  �b �X�!��Ǟ�GO�ӎ;-�������E};u}����Z�5^��j���X�m}��\�-�             t�~_}\��5��G���4 ��� 8HI�������K')�?���_����կ�_L���v�޳U}s}��ݪX��X�ʊؗ�             ��^��R|���O��$�� �^B1 ��!��ķ>��Xr撨(��ԞSVR�,h;w]�+�|����3?���5             ���﬎y��Ž��� @:	� }z��o�������m��I�ˇ�w��N\7뺸a����K�%�             �G6�l�?�_������b��� ��P@ʍ8*X�@�=���C���.�-��zE\yϕ�}��              >���㮍w��c�����F�޺(�]ک����G���q4T5U px�b R�1g�#_}$�����=vv���^��~zY�ݲ6             ��m�� @�� �Ԭ1��_���1�t@$MEYE<q�q�ݗ��7W               ��P@
M1)�mɿEyI�!]_�\[k��κ�Q�X�M������2�L*C���#��A�GYIY��ѿ�<���b�m�b㎍               i&�2K�C�P�"1�Օ����/��elؾ������$�����FM�Ϗ�|\��℡'t���X̊?]�8=j��               ��P@��z٭q�?q]K�%��p������r�!?�5(��o����`�ج1�bəKbѴEQԻ�c�7t\ܾ����+               �J( Ef���O]���{�����]�����{<�并�����ޅߋS|���L�J���]����               i$��L&n�얶�ٻo\��u��zD��ͪ7cᲅ�hڢX�pi���u����7�)7��|.                m�b R���BL=vj��{k㒻/�g+��#������/��_bXٰv�L19.�xq<�ڣ               i��P�e�.�1��tz��c'pt}���i�9-
��o�M��#���Ϲ�ù������,8*�����/���B<��D������s�V(              �TJu(fڠi1i�N�1pD G�	e'���ΎBv����x(f��q����p���|3V��:���������=��iw~���1q��شkS               @��:���ry�s�����/�����{�˧|9.�tI��s�}�               i"��,lw<��Ƿ�V��$�~���œ��{�>h�5z#              @ڤ:��e#��uz}�B
�F���+�6��qd����8uԩ��=��ظcc$���q���c�i���8|b�4:ޭ}7                -R���S���N�/++��jll������$j�TI��ΎL&��ܝ��Iu׺��Ŵ�5fV<�               �"ա�48{��펿_�~<�'"���|6�To�1C�47���B1               ��P@7mԴvǟx�hɵDR���x�w��_�����:�L               �S	� �p���l�����H���|��P�I'               ��P@6�t@�,��܋�I��;�;(F������               H���!'D&�9h|v����t[j�D}s}���47���B1               ��P@6�|x���Լ���"���|l���FM;h���               =�P@6�|D��;��B�s���C1eB1               ��P@6�lX���ս�bg��v�+�*               �B(�+/)ow���.
EG���g              ��H(�+�]��xsKs���M펗�)	               H����P̾�(EmJ�J               �B(�+�S��x.��B�?p���               �DB1 =X&����W�W               @Z�                 $�P                @�	�                 $�P                @�	�                 $�P                @�	� �Љ�N��O�<
���               �N( �.�xQ�	               ��.سgOlܸ���KJJbȐ!1t���ݻw                 
��.����u��}�L&�w\L�<9F�                 �K(�������1�                ��"s�&L��N:)JJJ                ���:�X�U{��ڱc��ԩS�"1�L&�#���!��m�&F>                �$ա����������KJJbʔ)q�YgEEEE G^sss[,��	�                ]��PLWd2����c���P(nXuC�����'�o�               H��N������ǖ-[��K/���� H�����               (l��T8J3�]����E������+�F�Њ ���LCTe
;|�=p                tE�C1?o���]X�����X�pi\9�� ���[��盞               �4Iu(�p�5�Ţ{�3o??��Qڧ4                 >B1��_���Y~��4bR                 t7��n�iצ�y�̸c��hڢ                 �NB1ݤ��.����X��Uq��ۣ_Q�                 �B1�l��e��������1iĤ                 8\B1��M�6ř��w,�#�:��                 8B1�����X|��x������Dߢ�                p(�b>e���c��u����1�bB                 t�P����W���O���q�iW                @W�!���q���ē��l��/�                 �!s�-[�,^��B,�zy�<��                 �$B1G����z̸eF�<��X2cI                 |���d���q���6�T����ѿ�                 �G(�([�~Y����X~��8y��                �Ǆb���x=f�2#�����7��f                 �wB1	�w����G�&^��R��EYIY                 ��I�e�źw���k�ǔ�S                 ա��^�ѧW��k���͍�Ǎ�Y��#%�J��OQ��lC���                ��UR��o���4pR$֮�����ԩS�O�T���\y��q�G!�ڋ_���w               @g��$�֭[���&�8�8p`                 �#S ����駟�ɓ'Ǹq�                H����fc�ƍQ]]ӦM�>}��                 -R]�k�����QH~�������cΜ91x����inn����ڷ,��               @W�:Ӵ�)����д��C=3f̈ɓ'�IKKKA���.��               @W�:SȲ�l�]�6v��s�̉���                 z&��WYY���1o޼:th                 =�PL�{��x�Gbƌ1y��                 z��"���ڵkc�Ν1gΜ(..                �g��a*++���*�Ν                >�����.V�\3gΌ�'                P؄bz�l6k֬�m۶�9����                &��n˖-���Ƽy󢢢"                ��#�����r�ʘ1cFL�<9                ��"��l6֮];v�9s�DIII                 �A(��ZC*555��UUU��͛c���1jԨ                 �O(��r�\444D�~ΥK�Ƽy�b��ّ�d                H.����f��jժضm[,\�0���                H&���{��"��Ǽy�b���                $�PQ__+W��.� F�                @���&��Eee�P                $�P                @�	�                 $�P                @�	�                 $�P��e2�(..                �����>}��ȑ#                 i�b                 N(                 �R���r��f�������o              �4Ju(���.�Uo>4r�Ȁ�����m�
|��               �KR�                (B1                 	'                �p�ŬiY2���Jc��������A��(d�               ��Hu(�����GNϞ�t�s�c{��                H�T�b                 
�P                @�	�                 $�P                @�	�                 $�P                @�	�                 $�P                @�	�                 $�P                @�	�                 $�P                @�	�                 $�P                @�	�                 $�P                @�	�                 $\�C1s+�ƨ����:3 ���db�����h�5               @g�:3g؜�4pR�1��$�䁓��QG!{tǣB1               @��:                P�b                 .ա����H�               �T�b�j��jU�c�9& ������m6�       ���+N�(�p<��Sq���"       ��Iu(        ����cXٰ��1��        �I(                 �b                 N(                 �b                 N(                 �b                 N(                 �b                 N(                 �b                 N(                 �b                 N(                 �b                 N(                 �b                 N(                 �b�0�x㍱{��H�g+��6<�c��㢡u�sƏ                i#�骫�
"z��W<���PL��~q��s               ��#                �pB1                 	'                �pB1                 	'                �p����5�j�566t�\DM�=v�|                tI�C1���Ş�=������S>��={챃�                ]��P                @!�                H�T�b��ث1�оt�l&�{��                ]��P̊}+��4�o�/8��|�� ~���                ��:                P�b                 N(                 �b                 N(                 �b                 N(                 �b                 N(                 �b                 N(            �����o����߹�>�9�/q(�H�D�Vh*�Ũ��a5�Q��J(h6�:,�/�RUQeӑʂJH��ĂQ;�tjK��R4�����v��>�3�}3�$��㜘�������^?'�mE��5    ��                H�P                @�b                 '                �8�                ��	�                 $N(                 qB1                 ��                H�P                @�b                 '                �8�                ��	�                 $N(                 qB1                 ��                H�P                @�b                 '                �8�                ��	�                 $N(                 qB1                 ��a͛�o����tp����bk���]�˙_                ��Pk�8�F>ܢ���8��;��               @b�bȍ�Gb�4@�?�ؚv�gd��z��ڼ                �P��?������
�_bG�t;Q�'�V                M�                 qB1                 ��                H�P                @�b                 '                �8�                ��	�                 $N(                 qB1                 ��                H�P                @�b                 '                �8�                ��	�                 $N(                 qB1                 ��                H�P                @�b                 '                �8�                ��	�                 $N(                 qB1                 ��                H�P                @�b                 '                �8�                ��	�                 $N(                 qB1                 ��                H�P                @�b                 '                �8�                ��	�                 $N(                 qB1                 ��                H�P                @�b                 '                �8�                ��	�                 $N(                 qB1                 ��                H�P                @�b                 '                �8�                ��	�                 $N(                 qB1                 ��                H�P                @�b                 '                �8�                ��	�                 $N(                 qB1                 ��                H�P                @�b                 '                �8�                ��	�                 $N(                 qB1                 ��                H�P                @�b                 '                �8�                ��	�                 $N(                 qB1                 ��                H�P                @�b                 '                �8�                ��	�                 $N(                 qB1                 ��                H�P                @�b                 '                �8�                ��	�                 $N(                 qB1                 ��       �M��X���r��lD�݌+�+       �LB1        �	���oƫ�?��lďN�(���       ؙ�b                 '                �8�                ��	�                 $N(                 qB1                l��阪L������:����b����                6�w��n<��#�����n��l6��j�0��F#߳�ެ��l����r�r,�c����y���G��uR'               ��+
144�O�Z����"1YH&�z���Y@&��~��ɑ�b�����4�^;��\h]��q�}q�v�׻���                ��,(322������e�V����fee%�B����_.�czh:�c��>��Rg)�\l�@�\�\,4b���Y�b                ؒ�����p>�y��`����y8&�W�w��u�Q+��9X9���P�Bs!��y@&�ݜ�K�Ky�I(               �m�X,F�Z�grrr��,���bV2�,//G�ټ�3F��q�r8��tW�l�l�����\>�?�(�                6���(Ky��Bq��/
���t:7�c��L�w�ݛ>�Z�����|���]�����\�Z8����1ߜ�F��Y�b                �4O���|2��ɘ��;F�=�=���7�T������[�w�sS�2�R)j�Z>�k47�c�^��VkCg�G����|V���b�b�Y���6f�R�R���b                �\|X�0�w����)���/ľ]�b����Wۗ����v��r���Ǒ��|��n���1����F�k���|�=���Jw%��1S��'��,4�;�P                �jw�1�4�ϯ����犅b�Q�#��S�'��'�������;��o�r��Z-����n����xL6�fs�gT��8\9�Ϫz�gg�h�l}6��6�F���?�                ��,�rv�l>�9���*��C����C����/����^�x���x>�:�N�����c��L�^���b%�T��vF��[�c�>��c�=�V�l/B1                l;�n+����|��Eb��7�̣1G&��ǿw���{(�JQ���Y�n��h���R��ng�m��B)��+���W~F�s���i�ğW��5ދ��B����K(               ���i�;����z��Z�92y$ߏN�C㇢Z���r��w��gU�^_��d���Jt�ݍ�Q(ǽ�{����׮�ѭ�lcv-3S��K�K��!               ����Z��^�m>���b����<�O�Ǧ��Tej�gW*�|��ٓ���W����1Y4&��v�����J��g�rg9�s�~���k�řƙ�o�G���#       ����P(Ķ�����.��W��Y�ta)�{� ���Q,��+�W�P������_g       ��n��Wf������=���7Ƭ�c���N���gī��u:��pL�^��1�t����hi4�T��s���b��gb�1���Xh.���ϏP        ��D剘�M�vs�̙x���o�9/f�_".^���W�X�/��O?;M�Ўg��      @J.�\�s�s�X{�v�c2�R)j�Z>�[��\�z5�d��D]����ڗ�YU��c�9�d�"2��`��                �-��x�������<"sh���ϮV��LMM���HL�^h<�R�����|V-w��Z��k�d���>��t�x��'���P                �����N�S��=�����xp���5�k��
���c:�N�YZZ�'���vo���h�=�Mvf�\��'O�ۿ��c����_;q��!             �⾱����|�
�Bz�  �AZj.�O�秛v�ʕ�8}�t��9��/�q`�@<0�@�>���]Ã�d����R���J�&k���������`>�]>�ng��.����=|��?��ɦX,��s�=w��l�z���{���	r�N���K/���5B1        ���*M�v�����������4�+   �s�������w  ؞�������,7�j��^[[ɹ8w�3^r�?�穉����N���oś�F(       �u��Vblx,����р��������,�n=        �                ��	�                �c�J�����L�v����               `Ǫ�j���l�F�Qx��go��                ��	�                 $N(                 qB1                 ��                H�P                @�b                 'C�{�}/~���܊n�                �P����                H�P                @�b                 '                �8�                ��	�                 $N(                 qB1                 ��!�Jz�W�O-                �EB1D�����;�P               �-�                H�P                @�b                 '       ���K�(�J���ŀ�
�m���YJ���o      �O"       ��M�O�de2������ԍ���������,�n#        �                ��	�                 $N(                 qB1D�o`�|^      l;'�x2Fˣ��\�����]�]<�gb�iw�       Ő�       �uy룷b[�( y���W�*       ��I(                 qB1                 ��                H�P                @�b                 '                �8�                ��	�                 $N(                 qB1                 ��                H�P                @�b                 '                �8�                ��	�                 $N(        `��N       �s	�        �n��F�.�����������=v������ ~���b'i�Zq�y*       `��       `ݎ���Do"��������x���}8N�:�f3v�v��B(       �b         ���z(���/��B�;w.    ���Ft:�   �Ai��7}�P        ��w��8q�D���+���    ��Rs)�F   �������F(       �u+��1�_�M�&��}��Gc������/G�� �_��L��\���}�(U@����أ"(F��u��$�S<����x4&�$�ģ�E%�1���B�PD@@iK�]�|�|����.�����\�{��<�����      sy�        ��z���)�Sd�u��4V��Ot��-&M�˖-�LSZU1'       `�'        ���	'����J���       d�        �������;�s�=���       d�        �ҽ{�hݺu<��S���Gc�����       �K(         �������'���^z)��m�F���       �_B1         (777�=���޽{<��CQZZ       @�%        ��z���:u���?>��        '�        �WTT�{n<�����/       ���         lrsscذa��.���?�ׯ       ���        ؎���;:u��ƍ����       �8�         lg�����΋��~:^xᅨ��       �a�        �egg�����k׮��C����       h��b         �c�z���.�(����?~        �P        �v�U�Vq�y�ų�>�'O����        �         ";;;�8��޽{<��QZZ��K~~~        _%        ��H�bF��&M�ŋ       �0�         �͚5��;.fΜ3f̈���        �-�         j��Ύ~��E�bʔ)�nݺ        ��         ��ܹs�x�1iҤX�xq        ۆP         լY�6lX̘1#y���       `��        �keeeE�~��cǎ1y��X�n]        [�P         �֩S�8餓bʔ)�`��        ��         6I�&MbȐ!1cƌ䭺�:       ��%        �&��ʊ~��Eǎc��ɱnݺ        �P         ��S�Nq��''c1,       �~�         �E
c�С��o��/�UUU       �-�        j�U�VѪ�Ud�f͚������ڵK�b֯__'kT               �&��ˏ����4���Fu%�<xpL�6-�,Y���U�T                @+((�A����o��vTWW       �e�b         �sYYY��{D۶m��^����       ���b        ��wKލ��>�L3�� ��;��~hLxaB|���M�YUY        B1        l����ia ��ia�8���⦩7�'�06Tn       `��         Pﲲ���.��#�-�(       ���        `��e@̼lf����1���       ԎP         [U��V���⦩7ŏ&�(�+�       �8�         ���������c����ȱ#c��y       �'        �6��̾lv������       HM(        �m�ea�w����߈?��(�,       ૄb         �沲�⒃/���#�s��       �	�         �`�۩_����8��1nָ        ��         �gĆ�       �/�         �����x`�q����럾       �W	�         ��,*Y��|{���M�lݲ        R�        `�+�,���k��?��bM������       HM(        ��.?'?��G�&��nY�2       ��b                 8�                �N(                ���                h��b        ����m#/+/2Myvy,���v�g7�9j�����UK       �wB1        �ڈ�QT]�擜O��/>�m�ov��;��񊬊����       ��P                @'                ��	�                 4pB1        �ZQ��h��>2�ڵkض�5k��׼��U�E|       ���       �����0�02M~~~ �Vnnn���T       B1                 �P                @'         �Ԧi��ܪst-�Zt���(jRY_|TUWŪ�UQQU�W/��+���Uc��       [J(         RHD`uG�~d�۩_��y��ز�&�����\83�/�O��T�2�����       �B1         �O�qH����ql�c�M�6[�^�V����z?=���lݲx������o���       ԆP         ۽���oT\~��ѳ]�zݫmӶqv�����������o�}QU]       ��P         ۵������]�����{��a�{��d��G/�g>x&        �         �K�
[�u�]�p��~(�Wǽ�������>|a�.[       �τb         ���n�;&��=����dT�Q���㸿|�A       ���b         خ��Q��YF��V�������/ǉw���|       @�P         ۍ#v="�h�n�}+�*��eƻKߍOK>�ū���cu���,/'/��7���M�C�ѱe��ٮg�h�#r�s6i�6M�����{�mpL�75       @(        ������o��u$���:^���x��'bʜ)1}��(�(��}����?����sh��ZݯY~�x����[�Y�f       �7�         2��v��g���Ϳ�����-So������x��[�wiEi��ы��5O_=���s�?7�s�w��I�F�۪�U<t�C��w�b���      ��K(        ��7�1ѥ��F�)�(��\�={]�)[So���e��"~=��q�7����,�r�Ҟ���1�~�� ��m�G��mR��Z�V2"��z��M��8^]]3�      2�P         mdߑ1�琍�3{��8��S���ޏ����$��������z0z������'�9!&�9!���ڡ�&�?���=6�z3nԸ�ӡO����QpyA      �لb         �X����ύ�3���q�}gǺ�b[xk�[1��3��z������x�'c���      ��G(        ��u����N�vJ;�o�}q�}gEEUElKk���Iw��F�������m�G����[�̗�Z_y�=�G��(~��       �B1         d��윸蠋��_���(W��#1_*�,��ƞ�_�|�2 �9?8�����U�Af���F��=6z�^       ��         2�q����m�������)cN����hHJ+Jc��#����՘'�!����A��ӡO����k�;r�#�kQט�r~       �O(        ��t�>���]��U�`Ղh�>Z�Q����o��M��){�"��F]�󲳲��g�5O_      @��         ��İ��R��,�?���h�����C.��-�ט��񑗓*7�'?'?����Z�_<�8~��/���:      ��&        @��S�hY�2��o����h�J+J��7�5�\Sc֦i��۩o���kA���ر���>�{��qh�C�ٹ�      �لb         �8�|`�����q����1�g�=���?������(�����&ߧx@�P�v�ꧮNƢ�UUuU      ���b         �8�w�������Gc���b֢Y�o�}k�vd��-;�1=�I9[�ny4�o�5f'�sr\4�()-	2����      �/�        j-?/?���#�����m��䤼�TUVm�z��k��/|�B4&/|�B�P�.mw	2���ώ���o�g�=ѹU������yM��}N����       2�P        �֪E�hY�22MӦMض


�e˚ח����Z�[�n)�O[0-�W翚�x�6݃̓Ť3f����2u(&�x@�P      d8�         2Jana��l����}�I��ۮy�(�-���� 3|c�oD�v=S��Y�NL�dZ�ʞKV/��-��8g�΃�W�^�s     ��$        @Fi��,�l���ј|���ǳ�����PL�(X�v6f���U1n������S�wN�s���/       3	�         �Q6�Y�~U4&%e%igM���/>h���S�95嬪�*�N�?�뵻҆bF�?y�'ɠu�EA���ʎU�����5�,l9Y9��|Ml��      �/�        j�o�"�s�#Ӕ�/`�zj�Sq��j�����
rR����Ҋ�hL֕�K>��¼� 3���)�I*��L���ϟg,�o.~3�t�S�܎-;�1=����~�^g�摗��r���$�6u��I*+֯��Х�K���8r�#����mvNFb��lݲxk�[ɯ��o?�}��V�l��$a�f;Đ�C������m{D���rN��:o��x����?���k����      uG(       �Z[\�82R��F@FZU�*毝_'k�U��?%b+��C]�,�S���$��<i|�����6�Ʊ����y��<�����ypԃ�M*��KV/���^���ث�^5�WTUDޏSk6W"
��c~��>>r�sҞ׶i�8��!�ۥ_�������q��[�J�j������W�G��#Y[�]����,��������s^�[=��Lގ�����}��r{��ҭQRZ      l�         2����ig��Ū�U�X4/h�v�~C�ϓ�c�v����r��lM<���5��3����_����h׼],]�4�z�9���!������b�٩�Nqð�.���F��yS#$b/:�Oq�.�n�:=���_�U�����"n{��F�     hh�b         �(+֭�ʪʔч�M[7�PL��mRO|~+ׯ��ő���r�����5�Z�i<���qL�cj��r���Έ��1ظ�M��c�~,�v���������L��</�L�ٿ�o�o�.
r�l��MZ�O�c����1r���|��     ���         �TTU��5K�cˎ5f���%�-��ŮmwMy|����ϓ�-3:��Yi���5����D|F(f�vl�c<��g�w��u�f~N~�9�Ψ���{g��M"X����|i����ݾ�\�J|���lT�b     ��B(        �����R�b��q�����h,v�q���篜4~G�~T��j������ٹϦ�����[�*]�
[՘��q��e@���kAMM�ģŏ�*SU]s�͍OK>�E%��y~��ܪs�h�#�s����1⎘�lN46�{]�#1����d᪅QZQ훷O>/EM������nʿM��o98�Z      ԞP         ��O_�A;�q��nĭ/��E��!a���A�7z�贳���&#%�߰>��@���y)����bҸ���ׂ��d�'q�s7Ľ3���|Vc�����8$.>��8��	_��ĝ#��>{/�s�?<�_{���<���N�3%��W����3�=#�3�;Ѧi�����f�x���[����      �v�b         �83�Ly��]��$�He֢YA�ֶi�8~�����L�k$�I���ȸ��ˢ��4�_C{��`���2����c?�u֥=���2KI܎��ȸ����C��3OSv�q�hv�a��u��Z�p������|7�%�ĕ��2n|���É���==���k�\?���      �v�b         �8��}6��E]c���Ō�3��KD:��r�������Έ�܂���?~9��콯]c꼩1w��إ�.5f�����:1�y_�����Ǎ�߸�s�z���k6i�g>x&�q�7b���~%���8ަ{��[�I^���9�ω�o98�^\�5��[g�sF,\�0~t؏Ҟw����c�ƽ      ����(         ���~�_9?��W��wz�Ō�;2��E%��ݥ��[��ⴳ1���j����3mL\=����G����s����������ɑ�/}��������w��-����nߌ�v?*��ӒO��ێޤH�?����c�f;D�ԯ�DL�C~�|�      �zB1         d��^(���k?g�9��'k��FC�4�i��7*��7	�};�};�M9+�(�q���z����?;�g���UcvĮGD�������.;+;���K|�A\2�-�c�q�߯��N�)��8�?6:?��s��m������/�����Jyΐ�C�'�      '        @F���)�m�����q�ԛ��:w�sc�f;��=0���q=pt��co?��-��Z������8��,G9��Yq�����.����i�=zY�W�o�>��?�y�{w�;���윌	�3������Om�>*7�E.�g.x&�9�kޅ_      l�P         ������E�c�N�Ԙ]~���_��W�-_M���Ǘ����/~�b�x������v>f��M^�iw��$$�H�x�Q]]۳S�95�,q�Hz�BeUe�������GCw�~gDVVV�Y��r�㩯C�c�����#��yL��Ⱦ#�	�DEUE      4V����z��X�n]�]�6��į_�֬Y���ӟ7��xB1         d�?������q|�V;��q�?�����#��N-;���<�横�
���m��I9�l�g�ĻOl��_7�xS4�kZcֽM�8l��bʜ)�=�sH���c�t��oM��떧�:7C{M;{�����e��~�8W�PL��u`�4�      ��6lؐ�|z�2��ϡ�T��+WFUU�~?W(        ��uό{⪣��n��՘��ƃ�?�͎��o��q�����-]�4Z�q+P�vv߬�bC�M^���$&�9!N����{nϡ�D,g�6;��UVUƃ�����+���7�s�?7�-�a�t�N��xN£o=+ׯ��&E)�G�v�P     P'6'�R^^��-_�<2�         2VYEY\���qǈ;j�
r��3���6��m�0�0Ɯ6&��R�vҵ��lM�xu)ꒌa�3fژ�^����J�9i��{�|/�����?��%o��Ջ�|�g>x�A�b��w�f���>Q�{�V���9�c�^�S���i�      ����^�<?q�L%        @F3}L|w�wS�"z��>��q��gEuuul+YYY�S�{u�+����ދ?�������gENvN��[�ߊ��o�ړ�L���F�V�k̚�5��}G�m/�ۣ=��v6{��zٳ�֭+}:�I;[�zI,*YT/��\83m(&�     2���^JJJ���"�I(        ��VYU�~��1���#7������wf�Y6'�~���V~z�O���H9Kl���w���,h�1�s���v�m������ď�q��9��nC1���%�l֢Y�����6�KFz�mz���X8���M�b��Z�5RJ��    ��csc/�V���J�޿�	�         ��^���h{U����I9���c[����߿�����c[�~eи���u�]Sξ��l���ݕ6s`��W�^�Βwb{ӡe�����}T/{&���ϋ��{GCԱeǴ�����۾��~�Y"Ӿy�XT�(     ���.�RVV�?�t���+WFUUU�p�        Pk'�����4K���_| �N�ܾ1�`t��������:٣��$*!��W<�8�lҜI�p��-���%oǴO�E�.��>�?�:$��vl�c�YIY�]V�����mӶig�y����d�f;�  ۅ�8?����ǧ-��M�.   �_���|yKzIKܗ�!       @���jE�E�i!
`�j��G�/>�UEVE@c׼�y���Ii�c������L�6sV���'O�$6Tn_���$�I�Y}FQV����j[='_�)�+ ���~���S�9������    3m,�R^^������\�2����b          ��Ⱦ#���T1�G�x����o�}q���#?��`ھE�8f�cb��c{��������o}W������ܔU�EyeyگIa�P     ��b/�[��KIIITT���         �z4z�贳-b��/V�ow����ʴ��Ed�TC��TT�3za^�=�����K;�P�!     �����~%���˸˺u�|���Kb�~����@(       �Z��Ϗ&�M"��m���F�&5�/�������;�t= �a��E�b��ű�(ݐ�"Ҳ�e��۪I�h��*���Z��s�X;+++��    ��S^^S�NM��͛K�.h�b        ��VmZE��v�iJJJض�5k��ռ��V�F�
h��=��clm�ٹq�~��o��m4t9�9u���ҕig�����ʖZ�>���^���Y���?�    �媪��'��{�'֬YSo���.1r���s�=�y���������ˋ�����_�bE4m�4��������:�����?N���H<Ɯ������I|߸>�JD�JK�>X�nݺؚ��:g}����?.����c/���>2t�й��#         PQ�Q�FECS<��Q�bZ7i]'�|Z�i�Y���th�!�OW�N:��Xo�vj�i��E%�     ��ʕ+��k��w�}����ҥK\y��P��~`@nnn�y"��X#�IHcnH?� ��V(���J<��Y�E����������M�����������8q�3_�~�o}��>_(         ��9�^���O�>1���xu���t��ʲ���yM���iڦN��d�'ig{w�;�C�퓷�jc�I�N}�m߾�ӯ����c���     �k�ҥq�UWŢE�&?�������j��kGfggO�8q����/
�         �Ѿ=�۱ێ����)[���˨�����Т�E��a��߈���G�fm�I^��KV/�9��$�/|�B�1��GCU<�x�C1%�%ig��x]JDV
r�d����v�O�}�>�׺u��%o����n�,�Y�-_[����yߴ��}�     ��lذ!~��_�k$�.�SN9%�����D���>�h��?�'_         ��T�[7~�ƴ��L�M�Fb���/~z�OcH�!����o�[�a}<��#qó7Č�3�ƫ]�vq\����=��1�������5<���)g#�����,����U����Z7muiP�Au��럾�v�����Gyeyԥ������?'9�9���c��u��A;�v6kѬ     ��u���ܹs�m��;,N>�d���/^wWL�8qްa�n�         c�cp�H̚�5q�s7�˾���m'ߖ�qlʛE��5���==N�{Z��16.�pI�X�"h|��wf��䥜UVU�M/��J��'Z&,\�0.?��d��_5)����μ��땔����j�+���\ԕ��ue���lu�kA����ķ'F]�ψh��Zs>���k��i��V硘�:����J;���     6��駟���sss�?�adgglC��0a�?�b         �X'�}R�٭/��������R�%�h���w��H�eF���rh��c���o�K�ⴳ)s��{$&a���1iΤ8z��S΋oR(f��yig{w�;�JAnA2TRW*�*�ٹ�ư��R�{�e(&�w�{FC���O��$���{�{QVQVg���?*�,�5�2gJ     ��x�������ֿ���I�&�X������b         �H�9�q��ǧ��-_�?w}��٢�E<u�Sѳ]�:Y�kQ�x����?��
��]F�}���Q�8˖J�.sĮGD������j�g���cp2pT]][��}O��-;F]�����������6��:���C.������w}'�u��q�����So���ڷh��x�S�=+֯     �T�@̫��Z�{z��B1         d����
[����5.>[�Y����S�Rg��/5)�'�{"���/�,
��1J+J��7�j��7�?n�c4ɫ�S.�������O]]�����(�,OF��U��=��n�K�^ڢǛ��l�Ϣ�MxsB�.[��9���s��~��=m���e@��7*��?|>�-�;��9�����<�u|���-���C��z�p�;     6�;�k׮���;u�-[�h ��         ���%�O��{��u�߈�#��}N��СE�������?���AÕ����;2�����U�����))-��oOL��<���q���DUu�׮����Z8+v�r�ӣ�o�E�7[�Z�5�Z�y���;⒃/I9�ψ��;������=
s��$<�A�k~�s7�M'ޔr����|��q�=�m�ugH�!��Y:s�͍G�x$     `s,]��^�?���#+++���         #�㐔�篜��|��W��V�&��V̋%��$�שU�d���G�zD��ߙ�������(jR�v~ό{bkK�.ӽM�8l��b�ɵZk҆b����8�ߙ1v��M~�9�9qˉ���G}IDQ�;�h�״�,���z0���1}��M^;���;��e@4&}��q���N�vJ9O��^�����Z�΃b���7��D����"     `s�\��^��ܹs@C"        @�)�-���r��fTUW��~����=v�c��,]�4��tm�?��d$�u)�y\~��c�Ӯ��!�L�C冠a=pt�ي�+�w������#��[m��I9/P\�P��c�Q������;N�#J7��������%"%>��1��ШO���$����ꨫR�[������~��:oj��mݤu�v�mqB���Y�a}\2�x��Ҟs���$�V�=zY�W��z��5-�uM��ҋ�c��	     �\���wכ�y���P         g@�Q�[�rv����|��q�F�͊!��ū��'7<wC2��_#�+��ul��A�}G���c��g�6;���v����U��֖�{<8�����R·�=<����bU骯]+�ZMĊq�T�F=�f���=��x��Ү�g�=�~g�E]M�|e���W�Ua��ٮgԥD�)tٻ��)�횷�g��l�<�����ߤ�;�������?��ѩe����mXo/~;�w���o<�μ7N�����$�q������b���"����_��s�1%�%1z�訮�     h�����         2N�}R_�zI����:�+��S���D��;��hp�K���,��9<��cq��G�<g��B1�9��I�Cҹwƽ��$B �B1M�&D��|[����?IF@��7K9O�azdߑ�������5��Yk��F�fm�C�ɀJע�)�b��8m�i��E]K�zN���x�{/E�)���΍K�4�;�1eΔx�㗓��OW-ZFǖ�1�c�8&oJ�'�I��m�F�I8�����t��ĵ���L~-'ϙ|�A򺶺lu2��S�N1h�A�o�}��M�U�q��g��      ԞP         g�v{�<��TWW��^g�w�F翜��dd���+��{ψ���hUت����D����D ���g��'^��|l+/|�B�_9?m��x@q�C1���	��_N��מ����'o�UZQߺ�[��򏢾����8��Sc�艑������������mS�7������{�m�0ЦJD|���Q1�;S�w��=�]�v��檪�����	oN  �*�Ϡ�����,��i�|	�ٻ8;�o��3{&�e��&��"�5)!�j�P"�S����E���M��.��Ւ�U���Q$��Z��ElY%Dd_g�Y��y��Й��d�̼���{9�}��u͙��q]��  ꆠ         ��AU��������N��*kɋ�~���j���-����7�O��i�ZzZz���x`�A�1����ծW��dxH2 ��$��{����?��~H�CR!o}�V�ֻ뵻bP�A��#�_k��e��;el*Ԧ�=��Sq�'��	S#73���}�'�Ϋ�@���j˪8������L���¦m���Ί��z,  ���A�ƺ����lʬ)1�O   ��b         hrvXi��sku;�:��5����Gc}���Z;0s�W�O�Q��}�ח�42�t����q_4��>T�t�s����������Ćm�c���D�.���5c��1{ŧ�e'  ��IDAT�/O��D��}D���ѿC�]Z+s�?�K�$J�Jbw�f�8��G��'?����ȩ���_�|����+�[�^      �s�         ��tiݥ��Ek��vF��D����o>��k'f�~��8�K�W���y���hۢm���)U��\�f�Y1'ڼ���܏���.�+��}��qœWDqiq��K���0�xn�sqǩw�~]���>ĝ/��<uM�y}{�����: ���ÿ���5^㭏�J�<��3�$�n�s�����8��������J��s���3      �<A1         4)�陑��S�?P���ku[_��*k�e���{O����L�4(���A�|��s�9U���݀�]q���F�}��'�R6�n�њ/-})���Ձ_��<+�xL��m_���򲘱|F<2{�ݱz��J�}���G�m*��v��֢�q�߮�[��5�=��8m�i1���HOK�rΚ�k��w��?���ۻ�t�n{�xx�Õ��h�G;������*}M��im[�vq|��o��O\c�M}��h��f���2����pz<0��xu٫b      j��         ���٭+��V�-�jӡ=�����oņ�������U��.�]�x�ܼ2�Ι���?|=�j[2$��l�D"���]Zu�-;DǼ��1������O��ز}����AK5��`m�칟�Z2e�=����zG��V�z2P&�Ϊwbنe_~�����Zm���$)�s�?�L��DZ�j�+�����:E^v^jLIYI�+X���.Z�(6m�      �>A1         4)�s*�),.���d�eľ]�����Wwy�@���f�FVzV�46� ��k���j㶍u���++/��k�      �OP         MJ2Ƞ2�i鵺����+Zd���^A1k�VYkӢM�޲:       h�         Фl޾������H$Q^^^+��m��3����m�Gaqa��4��[�  hB�����<sr���<?   ��#(        �&���������̍�E[ke;C�W�w����
�)*-
   ��k�O��i    TEP         MJqiql+�99j=�{���]+��{D���+f��cW%�h�Ӻ�ږ�[      ��CP         M���ӪbP��.�k%(�m���_�����\>3jC��֑�V��~[��       ͇�        ��}���.�]45�[��a�h�"ڵ�����l�N��|��أ����<0���U�����DZ�������]n培�J�EQiQ       �|�       �����R��I$4�����>_>��٩��YC�Z����O�˟�<v���������6�n׻��e�       ͋�         ���͍38�B�^{��u�/欘��k��m�}�*�ɐ��6}����Vڿx��       �y        @�����TY��+bܔq;�����~�d�TY�ǢDm�*(fɺ%      @�"(       �j{a����M��u+hX��,�gV>S�{���Z��e�FAqA�f�V��<6��sG<����ۧ}�����p����2l�a��/\�0       h^�        Pm,����FeE l��Y��ſ���
�������>�B-�H��g�����.���99��)���lò��¿Gm�q`*��23��      �nĚ5kvjnfff���UY_�vm�l�2u��S����re��M�V�"==�^�������m۶Tk
�         �$�a�*�I�ҺK<��g�?��-{���вC��ܿ�A=��)3�DYyYԆ1��T�_RV�>�      @�J�������ܴ��(..���\7Y�lPL��n���S�>$�uv����u��g������         �$=:���p�ѭM�J�}���^����+��I3'�k�_�pr`��=��C����4�[��p{��Uk�_UP̛+ߌ�E[      ��EP         MRqiq�0�����;����va��޲:�mX����V٭�k뮩0����s?O�Ԇ���ƐnC*����+      @�#(        �&����>.<��ط˾_8�c^�T�m�(n~��-zA�����       ��        @�U\Zg���x�ۯDNFN�m��?�[�o���r3s���ί���d{L[0-       h~�         Ф�Y1'&�iB�����H������o�s������zv��mWi�م��֢�      @�#(        �&oꜩ������'2�3ke������+��/�:jӡ=�Y̪�v��       ͓�         ��?���X�vqL>cr���o��Z�eu������[�Em�x��       �'(        �f���_��?va|���E��]k4C���+����~S�9       �A1         4+�Ņ�_�������~G�1��/��r���?�����u�bنe�ܢ�b������gck��       ��&(        �f���4�~��T�Tˬ����i��X�um���   Ԧ����q��W�/.+   �         ���E[S   �JAqA�   Ԕ�                �FNP                @#'(            �j�ݮw��mW�m��X�ni    uCP            @=9e�S���W���b��ɱ;����Ψ�?e֔��	   �A1             �䘁���^P������rP�y�i/��`Z,^�8   �ݛ�        �m���"�GS�%}K,��4��i�「*��~�[27   �/�˓-�ZV�?}��b   �	       @���m��FS�<m��h`���ű��V�/I��      �               �n(;;�N�߾}{@c"(               ��N~~~���z���DP         MNFZF��u�h�毜�J�      4g]�v����y�8���A1        T[�N�Kf�hj�o�@�jݺut�޽B���mKj�^~n~̼df4U�~:(�]�n      @s֯_���Ϗ������o��F���EZZZ@c (       �jK�����M����%�J?_�M�3      �����vX<���u�~yyy,_�<z����               �ni�ر1mڴؾ}{����_�"n��ր����v��                vK�ڵ�1c��}��W'�Z�*f͚x`@CI$�w�q               �n���O�w�}7�R~��ǭ���:u
h �dgg��|"(               ��VZZZ\z�q�7�ܹs�d�����n�=��3��QZZz��ѣ7&� (               ��Znnn\{�����6�z�(//���KJJ��.��.�(9�HOO�C�?i����]9r��m�v
�        ���X�1F�ft4U�7,      ��222�[��Vy�1y��?~���q�q�}��\����H$�d�'�O޷�>����{QP         MNQiQL[0-      ��gРAq�7�ʕ+��W_���?>���زe˿ZII�N��~���馛R�۶m����.]���j>���{�g�k,[�,���S!3YYY����ڧ�EcѪU���̬�u�>���g%_˺�VAAAlݺ��g���Q�>�f���{t��'?i+�����p'�                ��t��9N:�Jk��ũ��͛7�BD>"�lɾ�jɾ��Omذ!f̘�3z��EP                �Jfff���ZM�V�Ԕ�                ����)**J�/
�Y�n]м	�         ����=Z������{cŖ     �jWBf�*��l�*df���Q^^���          �B��Nq�~GF��'��)()�[߸5     ���l�L2`��1�(���֒�

���0h�         �����
�v�I}N����M�8    ��S2`�m۶��3�A3�(�����3���7FiiiP;�    �f�/_{�ݳ��[��gN�����1�w����O�5%毜�Sk���'���E%E��hk����-�j˪�x�Ǳz��X�~ٿjm��qT���5�����ݯ���{��q����=��'�����o�uN��+��?8��x���   �ҳRA ;�UV�8�ױ��     ��d�L~~~���Ά�����#(     ���<;�qp������z�i��>.yY��W�u��b&��w�?�ʲ�R�+o�|3^\�b�%�d�����w�~V2�fꜩ�y���|~��-隧�٩�����n���  @�1=��v9�`g�0>Y�H���     P}�2���A37n����hJ�      �P��=RmT�QqɈKR}�P���=S�N�y͋ƦeV���ظ����|[�D"�zN   @c2��� �}��!�ĬU�     �?�4��!3ɾ���FP     @-ػ�ީv��b������<��@�6�D�M���������   h,w_j�� �U��     ��]	�ٶm��d��?�炂����{�Lrn]     P���L9cJ�x�qœW�_�c���7�n��^ã_�~�p��:�N2�   ���@m8���5�k�ز"     ��-'''�ڷo_���ũ��dx̦M��.���mÆ��#��h]A1      ud϶{�c�y�7��Ώk4��$��p�������l��[�i�O   h,:��#���ڐ�H�S��w̹#  j[ˬ�ѧ}�]Z#��+���i������    ��������V����     �X�vQL_0���f�FvFv���j��֦[tn�92�j~xeD�1�qΟΉG�?i��	q���FYyY����I��
   �Ř~c"3-3 jK2(�w�~EeE P�F��._T'k�~��   ���      ����3�?_�Ss��1�:����#���QFE�6ݫ5�MN�xd�#�~'n{ᶨk�6,�=���D�s�=�{��~#���3&�X���h�#   �>%bN�wj Ԧ��m�^��c�     ��$(     ����l�9+��䙓S!,#z�H��|}��#+=k���q�/���4n�n�طp���`�qX��*��zN���m�7�zT&�z]9��   ��4�Ǩh��> j����      �NP     �N*//��?�j�>um\s�5q�sS�0UI�n;��X�vQ<�Γu��θ�Ҡ�S�=5.z��ؼ}s�n/�S�Ͼdݒ�Ǣ�  �ލ0. �����1�����fn      �A1      �`نeq����}o�SΘ]Zw�rlZ"-&�19��bH,߰�����9ƭ'������o��2��76�~��Z�V�g�0tB���3'G�'   �O���>��	��2~�xA1     @�     P��/����x���c�.�V9�C�q�)��I��Tg��q��xd�#��!_�P�8lb������ѶG�����4sR�i�' ��!7'7Zd���&;;;�����-ZT�|I�%vƙ����td�#�Sn�XU�*      ꃠ     �Z�|��8�7G��;�r܉{�G8:�~��:ۗdHKeA1�{����Ƣ��je;����<��X�n�� hBZ涌�9-�����	�aeeeE˖?_2ʜ�F����Ǩ��.e�e�)}O����M      �G�     ���-���{N�Yߙ���U���c��N�b�/��6,�m{|�?�H�9Cω���z���&�M���)�֒A5   P�N�{jd�e@]�oL���=QTZ  �������z4E�,   ���     �#�z'�x⊸��[�3l�aqH�C��_��}(+/�)3�ďF��Bm��	q��צ����;��0�-۷�C�
   �O���L ԇv9��=��'�>  ��R   ���      ԡ;^�#�uطb@�U��谋�,(&i��Iq�QWD"��\���1��Ș�`�.�?q��J��Ν�
� ����(���Ԕ~� V�'��>_�ˋj��=��N-:@}7`��     �^�     �C%e%q���c�S�s�>'EVzV���>,X� ^Z�R�=�B휡��RP����^�UZ�wƽ 4=ߙ��h�>��=������W�d`@}ڧ�>�w��c���     P��      Աg?�8�ѡe�J뭲[�}����{���a��I�Ŝ��q�����wj݉�&Vڿdݒxa�   �i@������%C��~Y�     P��      Ա�Ң�:gj\x؅U��꠯�iP̃s��N�-r3s?��2�e����q�kw�x����8���+��;��(//   �O����0�����[cݶu     PW�      ԃ��}j�A1��V��ߴmS<4��J�]�v�NŌ0:���V�?3e֔   ���:�u��� h�i�qJ�S��5��l      �%(     �<���(+/��DZ����%�ԕ{g�[iP��^ã_�~�p���7q��J��?�uK   �S2�!'=' �i�O�IoO����      ��b      ���m�RA,:�����}���k��><��x���3�����DL8pB\����^+�E~���I�֒�4   P���c��	��ԱE��}d<��      ��b      �ɜs��I�ߣN�b���b���q��*�&��>}mjLu�?`|�dT�K�����y   ԧû][v��6n�8A1     @�     ����c���e[����,Y�d���m���>L�9)�ue$������#�����Wk��C'V����ck��   ���f h����n�x{��     P��      ��2�e�i�'�m�h���������.���_��
�s��S����;��8��ڽ3�   �O}��; ����c�W�     ��&(     ���ڲj��V9��e?�a.�Ō<&.~��شm��O:����k�KK_
   �O���D" ��1=���޸-6m     ��$(     ����"�E���ԹS�'�2��>ן��c���^��ʹi��!_��6i�(//   �/��Zű����$;=;N�{rLz{R      �&A1      �d[ɶ�[d�OP̖�[��yǄ�*��v��b�:�ѥu�
�e�e1y��   ��tR�����4@M�06������4      j��     �zR��cG�Dԗ{f�SiP��^ã_�~�p��J�M:����/�{,۰,   ���%�bl���u��_���x��g ��]2�8�K�ES4�i��g   @�     �����W��U�l�s����c~�INF��ŅQ_����dݒ�ݮ����a5�='���U��m'�}B���;��   ��4�����- ���.( �ԠN�bT�Q�}��    ꎠ     �_��[�}�����ɏ�-(�Ef���3(���<&Ϝ�}M�����<uM���}���!gFVzV��m�G�=   MI��O���+�W���z���y�y�2�忾mض!��l��E[S�%�[����X�~il(�ԝq�@c6l�aѯm�X�aa      �A1      ��cˎ;�o)��i��Iq��#�H|�?y��~#c����8lb��<0�((.  ��UzZz�6$��9,��94�v{�Wd���)v+6����gƌ�3b�3��_SKz���qP 4vc������I      �A1      ��k��;���èOK�-�,�G���
�s��󹠘}:h�2�θ7   v7�:������/�-�k}][w��>1ՒJ�Jc����?o�O<��c����GyyyPs���|
�����c���hS      �*A1      ��G�;��wPLR2䥲��1���ŏ\����X�?��J翷��x���  `w�:�u�6��T8��#�=h$=-=�~`�]s�5�t������)����_Q=������ANzN�������     `W	�     �'���a}���Q���P�~�푗�������;xl���]���gpf��'͜���  И��72�q�7�}N��-���ծW\9��TK�p&�<�0�QP\T��>'F�̖��8}��q�{�GYyY      �
A1      � y!��N����5��mپ%�Ν�;�BmⰉ�����:.:�u�P/-+��3' мL̞m?y45+2Wă�<��sp��qI�%��?yܱ������_���Ѩ��=���О�����ߜ
���[⃍��H$b쀱�;��=�rX����  Hz��Gbɺ%�;��̉�:/z��   @�     PF�iU���bN���DCH^�XYP����c`ǁ����L[0�E� ��&r#�<7���O@������'L���D;+%�:/<����W���t��M��6���ߎ� �{㾸a��h���:�ˡѳU� �݌0NP �/O��T���i1f���q?   ���     �zp���wX����h(�/~>�]}���P���ߍ��Z��3   �Efzf���q�諢k뮵�fQiQ�ܼ2�oXo�8
�
��� ��l������r�`����h��:ڶh��tKԴ�i�K����N�z�5䬸뵻��g���VDs7��� �����պW,ݴ4  v���������ep    ���     �:��`p���w8�!�X^^�
}��1?�P��!߬tΆ��7�   -�Hę���Nӷ}ߝZ#�2gŜ��r^�]17�\�f����x�ǩ�L;#/;/�?�t�'uA]���m��ܪs��I��ǡ��N��_�=n��M��p}4G��ǡ]��Q��Wc���[f�  �]2 �Ư���V�y�6,�?��s    uGP     @�ڠ���(_����L��4y����k"-�V���~ �� @��27Z�����e˖4����hݺ��K�'��V�����w�zG��mk[ɶx��W�E�ų��W���K�Gmڲ}K*|&�����S�:�#��j#���Ny���^nfn�`�bⰉq�㗥?w6�fwu��ӫ���1:��	q��;ck��  h���0ɀ�dPLM�-X�<{K���m���   @�     P��w
�rԕ;�w��ѐ��[��@��~GVk|�D �yj٪e�g�GS�v�� VNNN��W�|�V�-b����䴉�z]|�oEFZ�N�K^�6�i1u���˛�M�6ECxg�;����
=9��qN�3���;�����`�{��vQ|��oŌ�3�9�Iω�{ ��܌�8��q��� �1I��^w�uq���R�7�kk�ָ����'��m   ��	�     �Cɓ)�q����ҝ��;��j�$/h|���  �!�e�Ż��{���ǖ�����=~������5xH�++/�Y�J�?��ԝ�'�_��h��z�s��94^��/ǩ�N����k4u��9>Zg������������w  @C�ަ{\5��8��ĚTTZ�:�x�S����+   �?�b      �H��;N�c�c������pz4�{8�8��h��j��&͜   %+=�Cb����s��/_�e�_9?v�P�ז��j���wㄽO�o���T�s��ң[�n���� h
z���qP���  h(�s�ǥ#/�o�v��lQ�yɰ���>?|⇱x��    ꟠     �:�<�����:�p��O]���1�Z�5u!e�UI������   ���uK��n�߾��(,.��ն�m��g�6���l�eq�^�E"�����E�����7`�� �A��j����ˣMN�͝�`Z|�ߋ��   ���     �e�,�?����|;����Sw�kL�q��b�~��X�ay   4&�>�?�������hJ^\�b���e߸�K�Έ���u�_2P�)�ux�h�#�m^  �!+=+&�?>��ѹU��}i�Kq���K^   ��5���      u�O�>���Ɓ��ḭE[�.���ť/F���UYO��  ��X�aY�0��������hʒa8�4!n�~c\w�u1v���ti�%Ft MI"��1���/��E  ԥ�DZ�<&n��M��5��z���cꜩ   4�b      jAvFv\��R��j�����⭏ߊƦ��<��  ��l]����ٛ��n��%ۣ9yg�;q�������[N�%����Ǧ.lhjN�sb�zޯ���0  �¨���g'�,��_�潻�ݸ�oWş��9u�   h\�      �Ny��ϊ�|�;ѽM�j���s?��3'   5�y���sc�ظmc4g/��r��cD�k�.�����8��I���j��:6^�p  Ԧ/��r�丟Ĉ�#j4���\w�vw���   �8	�     ����ط˾qD�#Rw�;��Q��V�C.�|�q��\   �����XڼCb>����ڂ��T%�d�	��j����ȢGR��  �j����գ������Ѽu���goN�,,.   �q     4+{�W\6�j�M$ѶE��#o���)�v�}���Q0̧�w����?��z��   �b��?= ��>m�ā���� ��ի]������#�i՞��hk����q��o��   �=�     ���]�����6��[��/~>   �/6�Ӑ�?  ��q�	� vJ�6����W�y�W�]��=3�k��&Vn^   ��EP     @),.����9~��OS�  ��I' 4�w;<���+�� ��h��.~0����ߎ�-�=���,��P\���h�    vO�b      jٚ�k����~��Í   P}[tL' 4i���L���� �i��2.�����#m[����i�ť�]�W�   `�&(     ���o=�y0��(,.   ����iNo��S�������V�-  �]fzf�;�ܸ��k�K�.5��ϥ��˟�<�_�|    M�#�      ;a������7S'W&O���|�p   �EY�Yqrߓ�9i��:��yt�u�_ �Si��3xL�x�ѯC��MǼ��bꜩ   4-�b     ��I�l޾���܏���~l-��L���j˪�^���_�5[����Ҳ�شmS�y�u�^�=�/������W���ߏwW�[�kX��]\�k8���ј�+X���wYy�N�����h��V   ���{�r�@s3~�xA1 ����?*n9�ؿ��5��t��������;}�   h��     @3����,߰<F�ft����G4�fNJ����Q'��k��}  @�;}���h; ��_�Y3' ���О��O���8���5������n�_��WQTZ   @�%(         j 737z���[u��Dz�m�6�D�n�7FIYI�ܼ2��_�A��08���K�\�0NP 4S{w�;�}M��ol��+X7?{s���_Faqa    M��         �B�6�cԀQ1�ې8������[�W{~��Ϗ�?x=^�����޴X�iEPQ2 �9;��Q��N��pU  �C���q�QW����i�՞�%���;n��M��pC    ͇�         ���z�;7N��ؿ����V��v1���TK*//�7V����h���������-:đ{ �Yz"=N�wj�zޯ h�:�u�����d�%���]�yť�qό{�ڧ���6}   @�#(         >�>_���8f�1��H��m$��mH�]=��x�'Rw����Fs6�ߘ�L���.�yx������( ����c���������⡹�O^�,   ��        @��o�}���n���j�n7=-=N��	���[��e�_o�v47iqrߓ������sT<�� �?��������Y���a�EeQP��%5��b.����nݛݮ[ei�kj7���e�e��i)nY�"*����"�o�����?�����03g����<f��s��sf�0G��: ��~mv\~����   �(        �6)]P�|)�q�7�0��YK�,愡'�7�f����7jjk��8��qQV\ ��s���( �w6��;.��D2��1}�Dk�f���ڿ   �4�         ���l�3~���Ƹ�㢥(�+����1q��8�3��-�F[��! ������w�?�Y @�ս�{|��Ek3c���r��    ���         ڔ�F����?�u�-ё�s�}n��ӓ��w^�\6��8����>����kk�      �HQ         m�=��>�Xt-�[�WTWĒw�ĊM+b�ƕ��jkl���5��.�]��dF�g��1���(�+l���:(����}$^Y�J�� �u\���{�~/֔�	     ���        ���:�E��n�kV�^@�*))�n���/�5�K�>ҥ-_�p�Jb�o\|��ؒ��eO��k^��ښ]>>?����C�O���)��=���ٗ̎�o9<�\�f��E���~� u$�����O^�I      l�(       �]��=*�h�����$~s�ov�����:�YtO�䩟��?���ݾ�t��＜w̿#�yq���Ӈ~:�qf����۱o���_Ǆ[&DEuE�3���� �~g>+��8-�o	     @��         r�-g�#z���ۤR���ٻ�~5�X�F�<��ښx�Շ3cp��q�Ǯ��F���ǌ�;&��/ߍ�ͿF��K�ř�� �\��nq��G�Co>      i�b         �i��{l\x��z����䙓��%�ƞ���%1i��8q؉1�iѽ��No{�a����'�x2rA���{q� ��}|���      �S       �.��[�����#׬]�6��h���덻��W�Vg�[�W�?��z�9oΉ3��+7�������A�=(f]8+��S�m�D���Ę��DMmM�v�� ��Q�F�����5/ �;��w�W=pU�ʚ�    ���        v�����&�f��W��5z��1�c���t��ן��o?96Wl��������[��?�`��?��ی�=*�}N���]њ������9�ǡ�b  �l�ښ    �(        ���H$�G|a�믮~5N�vZ���l�~��8�'ż/̋A]�{��'^3ΌT*�U�����o     �)�         '=���kd�k�5�q�gf�YZ��[����ώ���T�'���_��9b��
       �E1         䤳G��ӵ�~�ㅕ/DK�������9����w=�q)�      h{�         �s�yq��׻�nۺ���%����qE��u��qF�������       ��P        @��{t���ջv�[cSŦh��o[�ν5.;�:k�:�zϭx.       h;�         �s��Nצ/�������-�I���      �6FQ         9�~��;�x��xi�K����x���cX�au��E1S�N       �E1         �!eC�b�њ�i��-�ٷ۾   -M������w   h�b         �9�:��w�鷞���eO�E�.�3?���   ��b\�q�c�붭�)wO	   �i(�         ��F��=�]{m�kњ������+
�
���*   ��l/�9y�ə�3�   ��(�         ���+�D"Q�ڛ�ތ�dg�7�HFiai��  `O�{T� 欑g��98   ���         �SJ
Jv��ڊU֗���ZqAq(�  `OR   �KQ         9���h�k���њl�ܲӵ��   @c�kd|�د*�  �f�(        ��RUSU�|*���(���;	og'   41   в(�         ��W��;�>����$6Ul�֢��t�'�m��   �F�W{��   ha�         �S�o[�T���:wjUE1��[��Tmlض!   �]ú�c�=&�����^�{Ei��(�+�<�]�um���՘���x���c���Y��в�q�I��i���[1��   4E1         䔊�xw˻QVZVgm`��������ا�>�ί޼:*k*  ��R�WS�N�;��bd��;�]ג�1��8x������̥cnz��Ţ_d
T�G��������O6����}��o��/�   @�Q       �.;���(y�k6�o���]���?�UpT����.OV=��7׽YoQ̐�!���b�n��;ߚ�n   �5G�sdL�45��ݭ���=6�����	��)wO�7־�O�I��\v�eq�1WE�v�|�邘k�6~���\N   4��        v�ؼ��)�)r�[���@3�;�w�O��3_��ޭ���W>�9A��wH�䩟Dk1���z�[�\   �;��.7�zs��%[�<<����8�g�Ŝ7���v�:�����Lh�}<���񍇿��x    {��         rγo?qp������&;{���/
   r�g�6n9��F��^�=��q���WW�Zg�̑g�m�n��ŝ��.����k��/�>   �=OQ         9牥O�;?�lhf����h�u���w��7�   Z���?��M�ݩ�S���{������_v�eq�I7F"���y��ŵ_��@    �GQ        �,��4���"?&h��g���;��ɼ���{�q�C�DKwށ��;�f�X�|Q   к��O��i�'����z������鉛2�?s�g�['k��O?�����W��*R�T    �KQ        ��[�nѻ�w���� �Wǎ�_�~u��k�#�4</}�ڬų2'�}�'�d�$����h�
�
₃/�w��/�>jS�  @�v�aǐ�!>���<��v��_9�+���8F�?:�G�t̼e�2%���`    -��         r����ޢ������G<�\pg�T�x^��ԯ޵�?��   �u�K�ťG\�Oo�|��c�1������b��5QS[��ѣ}��0`B�8��8{�ٙ���t.���8=�x�#?�᧓������_�{ߛ)a   ZE1     9�}O�k&\�UƼ��?^������K�|)��G�=����0��џ��G_�U�C{(.���.;�8��Y�����Ƶ�v��?rc?���ro[t[�p�w���q?�	}&d�����;�z��f�4#F���*7��M��ѯO�u�4(���>�٘�|�s�?>;�w�*��.�E�,�a�)OE�d��rO��)�֦�޿����S�G����X�u���{��3�0�YeV�V����an����ݧܝU�-+��_���\��6����%��Y����ܱ���oO�vV�/�}9���9;�M:)�r�W�ʭo��������\V�.}0���U;�5�^v�KwǍOݸ��uG\':)��?����[w�����㨽��*���w���ɺ�����q��e�{�S��/^��s3O�û�*��=���2  �����k��>]����壿�x�QUS-M�ľ����޵�	��_�   �nG<���ۥ�`����q�7Ƕ�mu��s[��̸뙻�k�Z������X�y���7wZH���bs|��/Ǐ����}   -��    ��.�(�+�*�����(��oA� ���^m-=�mn}����7?Q77��mn���>�]~���L$��&!7�cn"��:3��ޥ�s��$߻d��.�n�N���"7����ސ�{|����^��ɺ���yS쑍��%��s�oHk�� ���M��-�%��/ߩ��_���s�?�9ᮥ��_��eC�]��_�"�m   h�3F��ӵ��I�'Ŭųv9/]��/?�����[��.���a%1O��dL�99�\�f    -��         r�O��4�|̗��^��]s�5����/��b@�q��W׻��bS�:��   ���8x�N׾�ǯ5�$f��ښ��o?#z��	&��1�������ʚ�    Z>E1         䬍��Go�o���:k�:�]��G�����t�-�Hƴ�O�E�]��7�   Z����=�׻�x����c����������3��?G"�����\83s�T*   @�(        ���ÿ�0.9��mp���םx]\��+��]����#�>R�����'n
   Z�a݇e�B���(jS�Y忴꥘���8n�q;���5K�S����   he�     ���c۶mYelܺ��ܦ�M�*w㶍��n�'wk��鏹Ir+��nښ��w[e��7o}����irKR%Y�VTUԙۺmk��e���յ�;\O��d����r�j��έ���3WQ]�un���A�c�߻[�~�n���$�M�Gn,o�=���M���s�5�^��i����#�_�:���#K�f/��K6���  �}���WH��G�}5�+&^[����9���/��'^���Kg]�y�  @�7�렝���_6�}ܳ�-��ʃ_�<_   ZE1     9&]^��+~���dM�����8��ߢo�=�1�Ϛ,7�ڥ���$�5�ho�ֵ7�#[~nS�e{r�l�� ��<���1�;��0����tqgsZ��1������\���    7t.�\���5Kc��Սr����Z�����   ��Q        @����磥zn�s  @�о]�z�_X�B��ǋ�^��&�:k�_����   �>�b             ��E�_�uM��Gumul(���;�Y[�|Q    ���            �=dgE1�76���߶�ޢ�e�   �:)�            �C
���W�T6���,��i   �=GQ         9���,���1}������c���   DTTW   �:)�         '�1<n8醸��k��W����o��mT�V       �6�b         �i������OΌ��ǌ3�'O�$���$       ��P        @�ѻC�b�����b�ܩ1s���\�9       �%S        @�4���[��So��_�?S�ȒG"�JM�6⡇��7�ѣG�5* rպu��駟���۔�      i�b         hӊ�cҨI����W���ϻ=��_4�DM"n��z�q��)�r��o��K���Dt      E1         ��в����~=�>��xtɣ1u�Ԙ�¬���       hN�b         �95�5QUSy�u|2��c�=63Vo^w>sg�>��xa�       �AQ         9g�ֵ��q�����1����D"�ح��Ҳ��_̌W���O����i����   ��r�����>6Z�ޝ��w��N�����K�)�~uv��؍   4E1         �u��eJ]�#}r�#Έ)c��A}����=��'��m�n��bƂ���DMmM   @6�w�Mmt��M��b�    ���         r�[�ߊ�=���ؿ��1i䤘<fr��u���k��.&���oox;�|�θm�m����       ���         ڔ�+g�7�F�0>S�r��s���l���t�WL�".;겘�朘>z���]��rK       @cQ        @�T���?���̸�����a'����pz�%���L$c	�q�I7�ϟ�y���że�       ��(       �]VZR�E��k���h^���QZZwɯ�3�VQ]��pof�����ѾGVy��;�%�]�/��rL{zZL�?-VmZ       �;�        �ˊ�����(rM��h^�����/��D�vú�N�!�;�x���b�ܩ�B����       �]�(         v������^�=�=���Zҵ���%���}�͌��V�����gO�,^~��   ��H?�����E�W.   ��(�        �]�h������ť�.���&�E�.�S85
�
�ճ}ϸ|�噱��bƂ��v��    ����͙   �P�b        �e�+VG�K�YW�.�浥zK�*_Ug���"Z��ښ�+��G��Nq���c��)1���H$��wLf�p�q���b�ܩ�ȒG"�J       l�(       �]v��k#'�@3{`��g����m�3�.�1���8g�9�Ҙ�]68�(�(&���o�+f.��ι5�X�F       ��         h/��r\��5񍇿����c&�y���J��w��㊉W�eG]�.y4f,��Z���Z�5       h��         @#�M�Ɵ��sf\:��8y��1e̔8q؉���kPV2��c�=63�w���E�dJc��       �-�b         ��l���\����ש_|b�'b��)1�lh��:w���]�Co��~5       h;�         ��l����#�̌1}�d
c�}n���58+��      ��EQ         �a�� 3.��8~��1y��8��S�0�0       �>�b         ��T�T�}/ޗ��;ǤQ�b��)1a��       ��(         Z�u���mO���~%�y�7c���       �)�        �f֯S�8��s�3�>��
       � E1         �:u�S85&���>&�D       ��(�        �=$�H�у��)c��#Έ�
�
   ږ�z�}:��3�z��X�|Q��M�-�yf��{��'.��%   4E1         ��F��� �;��աWVYsޜ붭   Z�/���������Z<+N��iYew*���.��rKT�TFcI�v.�\g���$   ���(    �����K�5����a�غukV��'�07�thֹ]���ݧd��s������+�un���ur��w�:w��}��vNv�:wX�:�%���sGu���G�5�Y��<6���G��TlMe�;���_�����I�d�{dّ�������_>��A��cKՖ����f�[����PV\�un�*Y'���Y禿�>�;�Ӡ�s�j���o?�I���%���M�<4�^ַ]�:�=
zd�;�dP��.�.Y����`n�DǬs�+�/�zW�0W\[�u�莣c��^;NVFl��r�rh�k�/�����1�ݹ @v�'�M5)���L�*k妕qϢ{�O�4�[�\   @}�~��3%.t���㗋~   @�(    ��]2�(L6�cذaCVǗ�w�ܐ�5zn߼�M��/�_����n��wȾ��{`�3��s�w�;��>���?�;�|/�2��Sz��P��Z"��3��Qgn��-�����_g.��m�'~�Ir��g"�ʃM�[�ޥ)rK߻4EnS�
4I����1|��F��~Lf4v��N�3��s��rDf젦i���m��e�/ۓ^���� ���.�]|t�Gc��q��EA^�ng����c�?S�N�{_�7�j�      ��KQ    �@�;���zC:�D��>QZXE�EQ�_�lK�.�T*m����cŊ ��o߾ѣG�hKF���?�b�rU�VEEMEl������77���xf�31����� `�ڿ���r��s����Ҳ��^Z�R�1���6Z�ڴ*        MQ    ��z��S���>4z��3   v� Y�����#�F��V^]ϯ~>�������Ǧ�M 4�>��Y#ϊ�0F��Uֆ��g3̈?���       �R    �h���b��S�̡gF���  -A"�Z����8����q���������/�y1 ����=e�Sbʘ)q°"?���W���9oΉ���]��[*�       쌢    h���q���a�D�v  �)��k�<>>:���7ϿYa d�ʣ��;ϻ3ڷk�U�k߈iOOˌe�       �
E1    ���OҼj�Uѽ�{   �	�D"�{x��3>�}�޸�cS妀ݑ|����5�D*j߻ �'���%��̧R-�����������q���b�ܩ�ȒG2       4��    �C����?r}���   h�D2�rF�����+c��9uI�%�)�)r�[�oŌ�.@�7!�(���|u�:�U��=�8ڷky��7��91��i��g�7       �.E1    ���>*n�xS�.�   ͭ��,�?5n{���3?�T* Ж�%�b⠉1e�8��ӣ�]iVy+7��{��ϻ=-_       ��    @;�����ߎ����:>}�fmm�����[  h
��7�����+�Hd�����d�3�'�_2���ip|��/EU��9 mϘ�c2�0�>'��v�*���&{���:wj��½�m      ��)�   �&4i褸z�Ց����WSS��r��1�.�| ��.�{����g{aL^^^fl/��g�plL�����ß���[ r�����Qg�'�|"u�u�K�^�;����O�U�V       4E1    �DNtJ\3�]:93]S]]�y  �;҅�ۋ'�ҥ1����Tsh�C�o��0*k*>L��K^��56l�yG�.u����.�"��>��Y#ϊI�&ń"[�7���.�ϟ�_�       �'(�   �&pD�#⿎��z2f����*sB'  ��RvH�W[[���[��.�)((�Я����L�N��#��9
���(���\SRR@�*,,�����/�廕��̏�0�?��8b�#"�Hf��jS���G�g�~�}ᷱ�j[       ���(    ـ��;G'
�;�MMMM�M'_  {B��2=҅1��w���G��|!n�s @k׹�sL�45뜿o�{���]1u��X�fi       @sQ    ��0�0�3�;�W�^����a�1�  �=-]�~>�.���˫�6���xz���� �V�W��}��f�/?5��{       �OQ    4�+�2�uV�Z���tI  @sJXVTTD~~~�0惒�d\����_��*7 �%�� Ss�;c��5       -��    h$�w�?&�T�Z� &]  �R������F�v�"�H�֭�[|��/�5�&  ׭ݺ6~�ܯ�G�Q,Z�(       ��R    � }R�5���d^��������	  ��&]S^^�)�I&�;��5��������W? �kjjk����s�ƽ/�U5U       -��    h'<!�����	��/  Z�T*�)��`YL2��K�^�z�S ���w^�iOO�i�ŪM�       ZE1    �>5��-��   ����b��#�F�s�� h�6�o�Y�g����c�k�       Z+E1    ��#�û�a���2jjj  ���^STT�D"3�~{Ѩ���? ��l���������ɼ       ���    �Ҥa�v�^]]�   ��?��lw��GD�α�|] @k��bs���]       �BQ    d���4�s���kkk���2   Z��󚪪�(((�\/H�)�O��/L         ���    ����������+�  rA�(&///��d��	OP        ���    @��������Q[[   � ]�YT��Ř�w�?��c[��         �y(�   �,�����T*UUU  �+�E��B����(H�!��'�z"         h�b    `7�ܫg�ثG���ɓ�  �\�.�LŤ�� E1     M�#�|$�_:?����z�o��q��+���20   �=OQ    �};�����  �\�.�L?�I������    �R��N1��&�ާ�>   �~�b    `7�<(�6}�d��I  �\��(��� �IQ~QL;%r�=�����       m��    �M}J�dަO�  �U����ѣ�G @kҾ�}�z֭���x�	E1       m��    �M{����	�@˔H$�C��QTT�ڵ�d2� 4���P555QYY[�n�M�6eF*�
��I��         �GQ    즒�ɒ@˓��={������� �<����� S�.�J����ձjժx�w��5�t����s����(�+�ʚ�         `�S    ��(��	��u��=z�� ���Ϗ>}�d���~;֬Y@ː~�J����DQ        @3Q    �)}�dMMM -C2�����G�.]�֭�� ����lٲ��]@�K��$޻     ��g�~&~�藑��-�   @�Q    ���VI�������FIII �;�u��ڵ�%K�d
*����    �qL�;53    JQ    ���� Z��*��Q�۷����z �KQ �M��y隥њ���;��       ��    �n���	�����ѡC�  wu��)z��+V���T*�A�/ hm�n]���M��Nq���c��)�O�}       �S    ��6U@�*))����  ���b֭[���4E1l�����&�Lм�D��K^"���J&�q��3�0g�<3J
J       >HQ    �&E1�����9��ܗ��������z �CQ�u��%:u�\Ӿ}� �Wqqqt�\w����\5���8g�9�Ƀ?�;�       �0�b    `79I�Wii�9ژ�;fN޶m[д��3
3 {��;�9����8��!����|cl��{1      @[�(    �V��W ���K:u�(���L �=�D2�|tL;%�yf��48#]�6��91}����pfl��       �-�b     h��E �=��Ŋ  ��в�q���c/�]�VƲ����w�ԹSc隥      @ۥ(    �V�]�vQXX �=%%%���555@����(�/�\�i٦ ��_��5��2��|Mm��ݯcQ�8��Sc��q��c"�H48cc�Ƙ�xVL�?=Y�H�R��%��T\u�U��v]�v�\֯_�]������     @Q     �O�(�����(�l� 4��6<9ic ���o�Sk���(�H���3�0�t~�U�W�3jS�1��9�r��g��͑��vX �u:tإ�p�s�      �b     hu


��+?��� �eR6$�;�`�1�ˀ��X�~Yܽ��:wj,]�4       `g�%     �N"� ڮd2  �\:u��8-&���>f��;���1k�>z<��H�R       ���         ��D2��)�9���c�½�Q���9o�ɔ��\836Wl       hE1         P�~��Ź�vq�2p�2��_w/�;�ΝK�,       �]�b         ��ס�C�v�i1y��8f�1�H$���|c�Z<+�ϟ�,y$R�T   �v�=>F��h��q���   �4�         Ц%�?`|��ϋ�v�ΨM�Ɯ7�d�af.��+6   ���N���8rь3�   @R        @���#��>�ۻu�w������,[�,       ��(�        �M�O6�O�6�o�Y�ge�aY�H�R��y<��c������M�4)�;��e�^{m���K>n�>}�m���=�P�����+c��ё�������n�qݻw�[o�5      ���?��ή�>����̝=�d&+� �����BYd���b�
J}���
�>�}����>�"}Ԣ��He�� �
��HX�0�d��r�9c	������~���5�s�����ef����        `zs�qϳ��q���N�v�c/������~���1ٵ���c����dr�����ٍ�����     `�	�         �nԵ����4��qC       �X�        �ݨ)�������o����uK       �X�        ��p�㊷^�=��~W�{u���i<       ����������Ҳӟ����۶m۱.7�}�         � ����I��������o�W�sU�y~M   �@}���c$�~�5�
�vY~�΍U�
   `Ϻ���zihh����?�^vD^����tww��c�        `J{���hlo�����gz�����q����?������       ��+c/����V�%	��r���b       �I&�	 �����^7��)�ZzV����8uɩQ�7����X:�p��'��$������� �{G�jq       ��Pc/MMM�����P         S^gwg�zhU:�V̍s��<⃱lβ�QTPgxF:^l~1V�vU|��_��^x(       ��W_�����Z��dYr?v&         ��B��;����V�����z^Ԕ�x�9s�c�~,��[�Z���v��Q�V       ͫc/����V𥡡!r�\0<�b        ��d�y1ټ�})~�w�΁�9E�첼��vC�1V��K2.��8s�q�����%�FA���Kb3ɸ�W��a����[���;       FK{{�N!�$����Kss�n�3>�        0`��GU�*&��0����軽Zwf|�T:�;b�C�ұO�>��C�<�q@�1PEEq��s��|��q������Z<��      0P]]]��2�R__�,߱mr?&6�       v��� ��K"/W���t���".8�x�!�iE�<G���Kұ���q��W�w�|7Z:[      ��v{�1�e��KB0�񚺄b         `���˅߿0.���8s�q����%�E~^���Hb3_}�W�K+�?z�G��ߊ[�%zz{      ��{ijj���2xB1        X~~~d3٘l

Fc-///�ى�����#V=�*�*��y��~�����x���8g�9�x����ߎ���?⩺��=����e˖�v���>uuu1-Y�$jkk�]��|�=������c��]�z��hoo���������~�566��?     L<�|���Oǫ�'�&����       v��d`w�Ϙs��d����ؚ6mZ̝�����ގ�'cBI"/W���t���".8�x�!�iE�<G���Kұ���q��W�w�|'Z;[��%a�O|��]�W��w�S�����8���]���!�.�:���?��ݮ���?<eC1]tQ������m����]     0~$���k���O?7nL�.���;E_��5��<C�㸭��$�{<�c�r�ܘ�k�یB1         0B��˅߿0.���8s�i4���O���Il���j|��/�MkoJ�1w<yǄ9P      F[������;����a�?y�o�ʕqꩧƼy󢰰0���<_CCC������*�3���ٙ��&��e�nݺ�ߺ��b�s뮾�?������O�����        �����Z��y���Cϋ��X\�x�s�dK���cɕKb��u      ����E|�k_�@L"��|�#����aT��\.wP��W�X�n��o�8��^��P         ��皞�+ve:V�[uA��!�E$     ��q����5�\3b�_z�q�I'E&�	a�r�܏���k{{�_�{�=�B�         #��[~�����2�8��4s��':�      ��k��뮻n���+���e+..������d29�         &����XX�0&�ј�5��}��/޾��Q�-	      ���׿�U�V������Eb3�L�7�|�}�~N(        �Igz��x�o�
      `r������\.7"�WTTĻ����������M7���                &��n�)���Fl�O~��f�XA.���b                ��~�ӟ���˖-'��               `�y��c�ƍ#6�������DV(               �	g���#:��0��                0���׏���f�
O�b                �p���Ft���Ҁ�D(        �I���>��☬66n      ��r�\�T"        ��������       LB1                 �P                �8'            0J>y�'����>"s�dK�]~��W�%'\#�Go��n�,   ��!            0JT-��V��>���oT��v��    F�P       ;�d2         �/B1     쵼��Q�_~~~ 0u���?w         ��@(    ����f'�� _��         �"�     ��h�@_P��m��l���         ��h    `�������JKK��k4d2�Q�9         ��     �Z6�MO�ooo�}0u���G~~~������M�yyy     0\x��X�Ъ��~���   ��     �Eee娄b�� @EEE444��~��\.     �ȸ�ޫ�   0XB1     ��3g��͛G���d? 0k֬����GMMM ���i�QY<��eee�����~�E=E       �     0L��l����֭[Gl���QRR ��̟�D���4b�H�dS�-�L& �S�-L��l���|O�P_�_z�{       �    `͞=;��룧�g��NNX�;wn ���O477G.�����g͚  L\3�gĖOo��jɕKb��u      ��!    ��),,�}��7�|��a�{��Q\\ �CIII̛7/6n�8��&q����/���         `��    `XUVV��ٳcӦM�6gmmm: ��fΜmmmQWW7ls&���� �k��Ɩ�-1�lh����ܱ9j|h���{�            ��g�}"???�����+	 ̟?? `w-Zyyy�u�ֽ�k��1cƌ `����WbR���}��/��2�~��   Lv���(*(�eyWoW�v�   �G.�K�H���M�x�<����0R_���w��<&�     F��ٳ#���ƍ���g��O�LH�3I( �$	����!�qZP.����      I�|�?ǅG_����1V~ce   0~l۶-�l�2��ihhH�5����eee#�����t�G�LfP��     0bjjj���2=i���^�����c޼yQXX 0P�f�J�$������'y�uƌ1w��Q{#         `(�b     Q�p�3gN���ESSSZ���r�&9I���$��$q���� ��H"c�/N���\a%���;�����K�:�De����         ��    ��HN�Ob1�HtuuEoooz�~6� NItl����H"1����ϝ���t$�2  ��/���x��a��c.�UvY�?O�Oܾ��!�[SVs��       $�b     �0 ��$
��  ���������a�����7s��wŕ?�r��.�Y,      ��    �M˟۷o��v������#���'  0��-;::����[�����~JJJ��wٓڢ�h��         �>�    ��Es���u�ە��G^^ވ>����hii	  Iq QDF^[[[���#���s�Fii��[Z�4ַ� �������û]___S�UW]�\sM��z{{^��[o���k��7o�Sե�^���f�~     �H�         &�$v8������!0PI( ���h*Gr     ��'                0�	�                 �sB1                 �P                �8'                0�	�                 �sB1                 �P                �8'                0�	�        0`5y5��M6�3ۣ�����Ly�Λ����\ol�m	       ��b        �w�+�rU1�l,���c������첼;����|       �T'            0��= .9ᒘ���Hܴ��    F�P         0!UVVƒ%K}���ژ�-Z�\n��+**
��9s�鿧����2�̐�.ӧO ��:pցq�[����[��%  ���������3`<�         &�+V��]}�#	��+W�����?��     `|������l�0��        0`�Օ1+;+&�m۶0����b֬]��t�vF<       ��?�������[���B(       �+,*����l
[Q\�����       �עE��Rl޼yD�_�zu�r��d2�@N(               �	��o~s\w�u#6����c�����/�b                �������-�����#2������W�0�z{{?%               ��TVV����\�;�O<1`}��ϾK(            `���ȍ��+  ��;��Scݺui�e$|�k_�ŋǢE���=���%��                0�}����������Gd�O}�Sq饗Ʋe�FK.��qIIɻO>�����B1         ��mY����,���       FG�������={v|�{ߋ�۷���\.���1�>��x����l6`��=����ҧ?����b         `/����?"���z�����u=��       v��d��|g{����~7��a��x�q��7ǻ���8�裣��2�o2`/u��{��}ϧo�y晻�a,        �����W�{u��n����O���{z       �3{�����������7��M<��3�aÆhmm��hii����]����;����t$���c�ܹC���#���9��5��[^^ްϛ��ҿ�+���D~~���+��)�<����e��|�3�'��}�[N?��=��-        �����~��       �����8���w�����јm۶��IF���uMMM;�\:::b����u�g�#               ����f���:�5��LCCC�r����               �A��L]]]�H`���9�����M(                F�P#3;3��d^+2��������'                ��P3��Ff����C(                &������ECCÀ3ɲ�~/�                �_C������y��LSSS�����                ��P3��Ff���7&+�                `���LCCC�r�τb                �Ia8"3uuui8f ��dYr��                 LyC�̴����I�1��477��I>&c��b         �t2�LTW�d���=�=      ��+))IGmm����ޞ9����         &�ڲ����-1Y-�rI�ۺ.       �:�b                 �9�            �Qr��wF&��e�C/<    �E(            `�|��o�   `��b        ��la�d��f[����~���       @(    ��~s}ln߼��jjj"//oDKkkk���K�6_rB΢E�  �'�|2z{������a�]w��ڢ��x��M�P9�2*�+b�)--`lEEŮ�_�z�       �   �!�޹=��n��v%%%#�ٶm[����|N� ��K~7�PLggg���HK"1]]]{ܮ��0         B1         L:�:�ť7_:b���������<�������m?�;�s���5   ���]�,:f��\����]_   `d�         0�u�ŕ?�r��?�u'���m�m��{�:l���i���   ��U�*.<��]���ȍ��+c"8r��q��svY���qW    #D(       ��������1�tn�`lݾ����C_�eyOoO    �����l�.�?���ƭ��   ��&       ��m���RG c�i{Slض!   ��[4}Q�����<   ��O(                `��                �b                 �9�                �qN(         )/�       0��b         `��
�       F�P         RUIU��K��ö�������w][W[       0��         � ž���w]eq���z��:�      ��E(         aٜe�����nִYö�Y���՛����       `j�aB+������ƥ�E���촾��+�z{�Ϸ�tD.�   ��R1�"�+���]UUUd^���p+//����a����K�  0T,����a����=��l��Y�fEII��{���  "ޱ��]�bފa��a��wyKgK� `�)��Gq~a�yq^6�y�;�ߞ�Ξ����ѝ�	    ��r��Br���ly�.��ŕQ�-�i%Q�-�����c���oYyAq��y_=�������m���������m�Ե-�ƦΆ��ј��   П���(�+��vI�%//oDKQQ��  �555�6W[[[l�>��Y���Fii�OS[ �TW^T�;�}�]�|��t���ֽ�����w���M ��K�c�]\3
+�����Ƿ��ǸO����q��?�}o�v�GK�h�j��Ǹ����dy�������;�?    S�3G5I}^IM,(�s��cVQU�J>W��g�F�队�{���{� ^���ѐ������x�����M�:        `����bNŜݮ/�/���޸Ɜ�j?ӊ��9���w݃�?  �䂧���ba٬�ST�K��ܫ�e�q�{s���z96Ss���q۶�Η/��٘뾩�1^쨏g�6�ǻ    ��P#"y�za��8�|n,(���>/��y٘h��e�x��y��K��϶o�'[_�g�m�g�^����+        ���������?���.>����o��ݝC��EtQ��Ϛ��  �SZP�׼|l{r�{ɌX\>'*
Jc�I�.�̎��f�.��<�Qڶ��q�m[�m/FsW[     �P{-�W�+�o�XK+���O�*SA�Y:mA:v����/�?��l�m���qCl�Te       ��,����Y��Lf��.��$>{�g��?�sT�?�:0.?��ݮ�� ����������ba8m~z�����
��L�IƉ3��a�����yC�m�k��M/���    �P�V�-}9��Da*���$���3yi�=g�92]V����l�G�6�ھ�Om����         Ʒ9s�+o�J�<h����o��h�l�����G.7�p��Y���-Q�-�w}GwGܷ�  ��e������x��I0��5�dz:N�up��־�+M�1-���gc]�󱽷+    ��M݃=����/��T-���+�Mc(\MQE���xS�A�[��������񩸯��4$        �y�>�;�sQUR���~��O�M��)
�wZ��d�ӧ|:�^xt|��O���V���ʋ��c�~,.9ᒨ(���v���-�;o 0��:=���鯏C�Ga���Q^P�O]:I$�����ǹ?��B     �WB�WE�4�Wp~������i��VP��.MGbC�ָ����E��5=ݹ�         F_xy����gO�l�~��_s۞ޞ��M���O�<�^zv�ۼ��o�S^wJ�����O��l~$��EGwGԔ����ih��'�f f���*  ����lX� ����5o��%���)����|q��}:9^�hH�1�X��d�uw    0��b����iql��xӌ���i�#�wct,(���s���mq�K��/_z8lz:zs�SYr@��N��^����MM/���x��xtˣ�ló���      �w�#*3�1�l�n���n��9����@�vY��w�f�7G|�I &��\v�eq�>��>����c��k�x��B1;�^>wy:�F�����  SEI~Q=���ڃbE����s
�h�S\sf��������և㾆u�ѳ=    ���U�)���4��y]W�4�> �3y��J�MN��"-�������Η��4<=�1LA�E�q�Q���[Z��ϟ�y�����G~۶o      `�f�͊�\UL6]}7`l���f��^�;�=�����������~������������؏�'�8q�fz���o��q �I�0/�V����Լ!����U�)�?���HF�Y��T�Y�H����h�   �Q%3���E�f�1�X�(��aƭi%q����h�j�_��H�d��x�����3���禣��9������?�K�^
       `�J1+����N�lP���w�|7������>����}�/*�+b$$�3���� 0%<=|�����㈾�Ey�`|J�1GN}:�b�3��u�?[������c    `d�L!�ύ�f'�X%�E��R�-�3���m[�[�oZ��m��@�KN�$>t����q���       0�$���������b��僺oGwG�͏�&����\.�ӺǶ<��?��C��y�=t]|��O �dS[X<sy�1爘YTL,�El���,u�[�-�-��M    ���I���(��]��9<�/�LJg���]xB�W�.}1�����|��������8f�c��/����       ^VXX%y%1��������()�����������G ��S.�7�y���ȦG�=�~O�����v���9�����_����5��Kw~)>���GOoO  L��8�z�8q��qL�"/�L|5����y��9�קǸ�S�Xt��    �I(f�گlv��{t�y�AQ��&��LAW�4ڶ�M/�:n߲&:z���>t䇢��"��Wo�7    ���l6��l��藗��.����ttww�����{+y.&'�'#�|���y��ӓ>';;;�?�TR9�2fΌɦ��9��UVV3g������#�i��&'�m��ⲓ/R ���9���+�w~1ڻ������q����_W�k�����u[��_����|  �AMQE�=��8e֡Q�-&�L�퐪��h�j��6=?|���    ����d�V,�s�GT�n��3�-(�-~k���'[�Ī�����;����Gkk7���v��Ҩ.�������GIv`W8|���Ƿ>��vY    �gIp���4=�o��=Ib۶m���6a-	�$�����a�3y�':::���5���  ?��ޱ�i fٜe��WOW\}���|&��n�}�x�8��;-N<�������б
I����o�kW_����va `RH.�zƜ#�Y��d�Ζǻ�)�9���ևc��g�m    `��:	d��������J'���҂�8{�Q��ه��b�sw�3m[&���^|g�wu����x��7���]�/9}�a�O���������    v/	qTWW{ f�d�iӦ���$ʑDc`O��󣲲2���FlI|&���Q `��-��U����8˪�V��]붮۫�p�w�#��,��<��اb��*��l~6��Ե�ņ����G����=� `2pTvH�y8q��t<Ҳ!Vm�3�kx<r�\ ;;pցq�[�ث9����sޡ�Ŋy+b�<��    F�P��AΜ}d�=�Ș^8-��v����3������U���� "=��'��$�/>>�s�wbNŜ�n��ɋ9�_�;.    �_iii�I0���"466Fo���ӿ�9�ċF������f�Q__  �ē��z�7�e�]k�_3�s�w�ǽ�ޛ ��,?�����y.�J��N[K</�o�������ߥ�F�e���pɈ�}�ҳ�   LlB1Pq~a�:kE�k�qQ]X�Z����> I}��g���W��S?�C��и���;����n�;v�c��Q����   �Β�hEb^���ӧ�Q�^���$���F}�;�{hjj
  `b�@ �T��[{`��b����=ٯlv|�u���q\�ܝ����    � �L ��8e�!��'���i����?��������3?��[� bS˦8��g�}�����n��C�+   Џ�����f�XL]]]zb$���X>/KKK���#:;;  �vb.���x�� ��K.jyd�����'��������ϊ�s��om���U�Z��    �k�� vbΛ|�U�C��!/N�1_{��xrۋS�Û����������6g-=+.��   ��UVV���c��(Hyyy���$'%TUU��R�� ��I  `x$�$p�Sb��9{kA��Ԓw�3�6Ƿ7�\0    vC(fK`~S����SbfQU�pKޜ��p�����ן�Il�l
������������Olڧr�XP� 64n    ^VRR�A�hkk����`j+--�������0�(yN ����'~��|i�~nu  04o�6?.��X2m^�p[T6+Ƭm�W��5o}>    ��5�G�ү����ŧ�AFR$:a�㘚7�/�����h��0mnٜvĂ#v�Ͳ9��:STP��;,�ZxTP{@,�^�Q\P�^����1��n��u�������;}l��}����{L,��4����&�K��u�����6<�my,�~��x����w���<�?>��c���d撨.�������F][]�w���קG  ��$�/f��/��ʢ��9�ڒh�x��b���  {�{�{�����  ����"Λ|�6{Ed�n0��X_Z~A��nm���?�-.�
    )��q�"[�-8>Μ}D�e�FKa^6Νw\�8cy|c�O�-��
�j�|����,�z���O���Xy��(/��*���<{O\���q�o������[7��5m�.˓��I_=i��N��������MM�>��{̛�9�p��]w��W�c8$A��x����k��}7�l���.���/�/=�)��&_�����s����wZ��NqƁg�ǎ�X��������ۻڅb   �$3��LqI�(/o���2��?{wUy�}���d��6�$a'움���REVAl�V�^�*Z�k-�����V�
EѪXq��\pc�!�=d��I^���Uf�/'3�o>�#�3s�0���<��    T}����֭Z��V   �c��%m�iz���E
h*�{Q�&��Pww�q`�^����*���1'<�8G�������    @`�b,�fӄԡ��a���x��c���~�&�����\����BIV^V��I1I�����֟&�I�:��}2���i��=p��ݲ��/���§�2b-�z��;�+����Z�}O�5A��Wy��)�����F9Ʈ�]�/#��ŏh��i����Km�ژa����lF~�|�N-8���%�K���3����7�����V���'���    �.�Ŧm6��v��^&�*��!+�$�   4;�=��O�����ۛ�V��L   ��a����x�D%h.�����H�m3X���(*��/����     �������'�]T��@c��N�S�h�^������BAvQv��?�pT%���&<f�B��f��ֱ�����u���5��iu��,۱L�Ϙ�wlt���
ŌN]�uN�>��@�(񖘫�ՕH������؇��`��!�hb��L-ٺDM��7��O���6��    ��	��f���!��P��0I   h~���c�ǘ��R����3_=�uY�  ���:ݺ��dH�,�*��^uT�z2�.�      j�5[6��آ4��(MJ=Ka��$z���rB�PO꥿�z_+�o���U�h�����~�	Z<{���z�Ð�C�򶕺l�e�l�g��}FfF�1#���O��~��m�������q�'W<Y�c$E'i@�~Ǿ��ˋ�߸�8-��@���D���ֻ?~W��}{����������m�w	    �6�(KDD���� tY��'Z   XK�3Q���ܶ٢�腕/�x�q  ��laᚘz�fw�(�C�J���\/��D���PEe���      ��PL3�w�h��s;�to�+�͉����w�]�/ X%�$W9^T^T�>��������:�U�c�*|����D#���K4��q����>�[��w�KR���.�z�y?��S[#����
�F@ǈ�x+j���n#���Y�c���xΖ�t��w^����C����K�0ߐ�k��&�=��:Gb�_     ��iX���ń4�=�>_�_c   �4z��֣�Ճ=�w6���ּ�%ۖ��r  �`�9&E��_���X�#<B?��#�ߪ���|[�=Y      B��&���v�H�[�Ҝ��g�;��=j�5���l:�;W9~�s��q#����Fb����v|�׿}]+���a�a+8��h�%�)=9]zOЌA3p?1��}��:�3�y<S��,s��PL�3A��k徕����kt=W�KC���{�n�cddf�z�C���j#1F��>0�����u �U�+Sld��ĵшN#4��xM�;��o �O~\�ٙ�׶���;O_�t���q�?���y��Ϲ��b���Jo�n�#�S��     �x�^EFF�*��	��2+=��k�V)   8]�=RSL5���,���e���ig�N  �
#�qE�9���y��Y+�T�kL�O����ᕚ��c���      3B1Mhd������ڣ�T����&iDro�i�[�.�&F$�*{s�V9~��;��KUV�_��޼Ik�9m���Hۏm7�����{�ޣ��>��ξ)`���,��HC�jFKj*cG��;�:�c���n�P̩�6d(&�$O�������2�/:��Ǎ�ʳ_=�?~�G�>���u
J�Y�i�z����fph�6p�����mzi�K��߽�XKC2"4��i������/�Vnqn��O�N2W�  @��<���j����,��q'Tz<=z����t:ճgO@u�/_��K��*�v��ӧ����L��r������7
@hZ�~}�ŢJKK�����v�����R"R @�j�j�9#����W{�҂��p�B�
   X��K�=��]T�����ɩ�48����Mm/�      ��4�h{�~��"�k3D@�0^Dv�-�s����F���c�h�#ั�uǻ%w���_�1^]��f�cv��.'�N��ެ�W�a#0�π�t��;��Ǐ��223̿�� �c��1W����I]���vy��DQ~"iF��6���!��ғ���}��S3�R���T?�����j����ٮ�j�_#(s��W��4�O
;}%��d�q�5��YjH���ϝi/M3�.5�]���w.   �\MN�4���P'�Vu?��}��p�\�zk�;yc���B�M���b\\� �����yC�[���	S�  v�{�#:�0�����z{��f4fY�2^7  A��r�a�i�ek�E/����L���N���T���**�u5      ���idFa}N�˕�lb�Q���T=�]O�|W�5_ Vu�{��vt����q�����d�]�kT�+��}33q�qzf�3~�.�_������y���>�����?��ic#:��3©�����Q�F������hJ�)rE��w��N����#}T�1#|S���z������٫�^���?O|���ʊ�������4C�-L�oRcX�c�&ϛ��v    �F�v[�����|!4����J   �y����|�0,�{�Չ�����3�m��͚�j�^^�r�ߛ  ��֑.��}���:	6��p]�a�'v�c�-ҡ�      ��PL#1^\��n�fuEaAot���A�mS[��	h�&���i�Uyc��@���K�]p<�x��.�Z�H�)�}��z���m���w܈���_h��sj�O#��/co��������^��w()&I��L����H3H����j~�n������15>��X^I�ƿ0�^��S����tn�s�I�?d�B��~���������]2�"1    �Fg�0l6�|>�����Xeeer8Bh�Z$�P   ��<�s��	���g�9[���������~��|�r�}�ś�k.   @S;7��n�6I�v��`�+����3=��=e]/       X�i�Q���c�zƥ	mN~�?��Z-؛�7�V���R@KqV���ʌW�hG ���j~����P��o{�6������>]1���������:����ψ��׹��w���4�b��6�ۨ�.77cr\J\�i��SǨi(�8F��a�am>�Y5�p�Q�@�Yz��\C�u����Xi����f�i��=��E7���@     4���p�\.�8qBVaC�������xd%�b    �ؗ�OO|���������!ר��S��g�iL�s;QtB�6,�_������S  `]N[�n�6Q�Z�*�푺��ru�ӻ�S��L      @KG(������9=.����d��ǝ~����z�7U�-`e��zέ�ݸ��a�z��n���;�]��\9�ʀ�]�u��5���|�z�5o�<��I�I�k�yk�ӝ��[�=�����?��O��>j���7ڠcǔ����v�9F�ֽr���&P5�����~Ƕ�n��֐r�s��W��Αw�6��{^�|��;޲�e�p��    ����nB1hv��n%�b    k21��>zH�;7��ꌫ�S��#����v���9�F/�y�܌�  �U�s&龞��1���P4&e�zƧ顭�j_�1      -������ѵ��(��ʆ&vדn�C�^՞�#��X�k@� ]��"�l�ϔ�J��6E�E��;��0L�b[��gՐ�����I����M&��X�P��ԣ��V���~hp�`%:�S�S�~F���,۱���#[t(��i��Ai��Is5� �����g�8f� W�+WC{�����b��cC�b^��    Д�P��X-���O(   @-TTVh���v�{w�����c�c���0�g7�G�?�w7�k.Rb,�Q��O����x�w�^����DG��{�`ll��?�|��aI=uG��c��Ҝ�zb���㎷���      -��m�ԯ�/��^�om�n=9�z�y�{���:����w�ڡ�V{�G�=i�j��ȸZ��ެ='��}L���ǵt�R5�o�^_���Ym�?�~C1FT炮�MoU��@��w|l�ט�fgƠ�Z���5��H����:�`L��)cB��.�;fL�id��vߡ����>��ic�:k����k��    �)������*�v����vb)   ��W�-ջ[�5���f�b���I9#�u�_�=ʌ�ۮ�]��z�毚o�g4�M�6i�ܹ��f��������b �1��]��|�h��(* �i��==�����w�9o      hi��S{g�~�k�:D���s�G�闪W\{�e���V�4��m��[cy裇��ZU9��YǌId�r5�EŤ��� NV^V���l�2�;�^�cF���P�=ܮ�>ɣ�W��w}��oDc~�1��mt��#Z�����;���Ј�#�Iy��ܷR�=��X���x�i�wo�݌���k�1cB     4���DY	���d��n��'^    -SNq����y�v�o���O]��衋�>���~����5/���H   �%���zNՠ���}���W����qi�ݶו[^���      @S"S�&�1#Q6� 6��3����(��$��
��x�=����^�_j��cF��1T�����k�1&�Т#N_���TgH�!���?���~���IƎ����1�V�3��XF���2�ݠ�coTc:�{�����-�ܝ����z��>�     ���햕�	=^�WEE�y�9!!A    �S��T���Z��x_xD�����G���W����6k���d��/�1TVV����v�$V�5����=C�#]XWg=1�=�u�v      �R�L]��l��e���j�@M�su���o6����Xٷ�Ս�n�7�����1���op|]�:5�E'�7g�:&v�;޽Uw-ݶ�F�2&��ؽBv�𴱞�{���]�љ@��e;�}�����ӎ�;���~�}m��^�s�>F��1��:U�}�ݦ�t��h��v��$�ر     �ILL4W_4N�B1����X���@(   ^W�|�
J4k�,M�?��,�It&��7�ۖ#[�`��[5������jݺ�fϞ-�1�߿_�/6����, �opB7��s����BQJT����:����V�l      ���%ce��u�	�C�vR�����顭�jc�V�z�j��?�����W��m����	]�e��MC1�ݯ�ؑ�7c0B0Ƥ�@E\�\��~�9u����>F��q�OFf�j#�cf���kuqϋ�?��"���V�����f����l    �ԌՂ���,h�'r���d%�b  ���r��l��6�$>>^ �����}���_�����B����ny�M�;Y3�4�;7"���;������>��C-X�@om|K�
�   j㢔A���D��lPsN�C��JٵD�Z)      ���Ԃ���=�����P7qv�~�g���c��� �9/<�U�W�]�i���vt[���:�u�1crX^I㝠r��D�����Z�kY沀c�d�@�g�Sgw:���=�����eF(�Ƴo�{�@��({�Ft�wlá:VpL���J8ַM_sk�c��K8    �<���,h)**Ryy�"""����xd%�b  ��f�)<<\��.� ��:����&k��l�	0�O7�	4���n�u�Ե��r���{���?�76���y^m  @U�C�h���0R ��XP��]'�}t��ٹT�'?       �"SCI�8=��ju�I�������S�Ι���-P/�|A+�U_�/�)�8O�%�����u`ğhGt�1#�RY�xoU���|��Y��N9�9Jt&�66:}t�۝��3��C���T���._����o���ƛ��/#�����Ֆ��9��OcƉ     �Jbb�v��-�0�5F���*��S��    �e_�>�~���mp�`]?�z]9�J�G��z_����[�ḿ5z�����W�y   �ɘ����KuA�~P�S�))"^�mSe�      ��PLt�n�G��RRd�ߴ���0V.pG���;ߣ��:�ؑ�Wֽ�lǏ�G�/iܓS�ڿ3�Y�}�*|�d�'��不��s�S��^�zd�ic����e;���<�([��V������$��)��������T%Pt����aV��Vx    @sp�ݲB1��j��˚�b    MÈ�ܰ�ݶ�6M�3Q���؞ce��t=#:������ɏ�-�јe��u�  �2�ڝz�����  ���Jt���-U�-      `5�b��-&U��{��#���K=S�Q��w����'���j�UxXx��.R���]��1�������+3p��8�C1���/��r}��3�V]&�   ���ƨC��'^���+<�qG(..n� Bc�_ ��j���U�C���o�á��m={�l�����:tH�-55UNg�!��7����J�HT�9|� 4�]����N���W����[�7ֿan�"-3�0�1}������c��jnۏm׼U����O���H   �$DĘsܻĴ���'��~�������+��P      ��p�t�Ƕ�#}g)�^�d8 uwAr?9�zd�k*��
hIJ��'��G�7�]Q�W%../�����K c����/���e��D���Þ��txS�ǹ�;���+���ˌ�㐴!~��j�*yJk�1/��w�Xy-�8G�a]�:  ��	����D����F�'���� ���B1yyyB����r� 5�=�6����،�]�*�0�σ�����
@3[��F��zF�(+/K�-�܌P���35{�l�ĥ�z_�[u��qs��Ʒ�ݱ�  BKbD�����Nѭ��t�i�?�����8_���      X�� ��:��3�E
@�;��C����.T��L@KQXx��XG����UQY�(ǎ����~���6sb����]����m�U�N��223�\%��]����H��ƞ��|����V��	恎a�*lS���"�E��{i�KZ�{�     @�Y-���>0��+?�:�    U�|x��z�.ݳ���:R���Ҕ�SQ}�  ��֑	z��l�uZ�5y X�w&����6�ס�      ��P�g���7=��! Mg@Bg���L�f��*�
h	{�;ڭ���حb[;��N�4"/ƪe?��L���Z�o��]6:}��}Tp)*/��{�6�0���Ґ�C̱�a'�n��C�CWd���L(    �:r8���Qaa���!//OF����@V���     �	c���w|ln�.�U��L2߳�m�9�   �?�9�5��5j������?������w�-<*      �����s��hN��e�	@����\���M���:#�b��h�V��~Z���Q�m�;����:�ӈ�����h���mT�}T{��e��b�c���Q(�Tl�.���������     Pwn��2���#��6^��
���4    �^nq��^`n=Z���3����wI�"  �N1)���%:b��qz��l3����      ��D(�?���I$�����h�k5g�<��ŕxK�'gO���$i�PLJ\��Ʒ8����:��X�,#�27c��g�ؽRz�v��w�!��1��.z��ct�G>~����w����c>���J����-G�hr��~���r�     @�������
����`��:!!A    �-Z  BK��$��{�#�� ��5���lݱ�E�+:&      ����_g$t�ݽ� XDט6z���������W&��6�03���F9��ϬrܸOu�����Ƕ�{���<B���ˋ�h�?F �&V�[)O�Gq�q߻|x�኎�VQy�Ƥ�	8�-#3Cue;��g�'�    ��3B1VQTT$��+���B�]~~��$11Q    P[	�]1�
�2K�;'  L�#]�ۏH`����s�~��*�      ��}R�����t9�x8 +��^���ڼ�B�UzX՗{�Ԥ>�����5^Q�(�xK���L8f�^���؋�P���0B.�x}C1�
�>���&����#�f���<Fm��ϊ�+���~z�as�iцE     �g�@Fee�<��v?�y���%    �	�}�]G�q���_n.�  pJRd�~���j�  �q�k�W^���\      M-��(=���H����9�z�H�_��B������>V�����\f�!�#1�]�����Fd�>223t�����@����
}��Z燡�S�0�����{���\}{�[Օ��|�纠�~�猜�77�i�L     j��v�J���ń���|Y���PLL�    �*}�����35{�l�ĥ  ��\1����F�7`E�#]����j��)/      ДB:�9&E��3SN[� Xװ�����T����`5k��jω=����w܈�4d(��C���؀�7-����g.7�����O�m�z��4W�ic�֙��
�1����������_E��Q�.��~�.�y��l]"     P;III���#?+�b\.�    ����T�4C��F}���׾�9
�W�ׁ�  �'��G��R��V`]�4��5�s�<�{�      4��Ŵu�5��l�ٝ`}�$��Ͻ�d�;�������3��㣺��e�.�?7����J�I�>p|�~3�R�E�����n�ic��kJ�)~o�lǲZg��M:�9r��h��iꀩoW���c<_��{����r�ǉԊ�+�_b���     h	�N���
�A���˓U$&��/   ��/���_���g꒾�(�Q�}�xK���w�Қ��dےz/�  �)���#}f�[L� X_��=��j��8O��      �BH�b���z���J����c\�!:R���|.�j����1�9l��Fx���;<�71�yşUQY��2b,�B1�p�~y�/ަ6�����~���]�u9�?�����O�[s���;޳uO-�j�&ϛ� �'     ��e�AS�x<����   ��ˬ!�4c�%E'�k_k�1�0/�y�\�  ���wv��qi�r�<�5{O�iz`�+�9     @��P�=̦{zNS�3Y Z����XY�2��`%�h��y�����wrw�;׾����،��Žc��5C�	8~���iF����;�/TS�-Պ�+�t��bÐ����}����g���a׫�����	�'��i/�7o��sV#�c�7��X]���     X��n<xPV`���#��   `���3��O���ғ�뵯E'�h�"��˿�ۃ�
  ���^��I�����]�u�H��Z*      ���T(&,,L�H�D:@�t��8�,_�sw���>�OSL99���Z4k��/������fmE挜���>\���z�.yJ�#�R�+����������ʋj}�e��jw���~UJ�%����ʸ1C�p���a�mh�KӴ���9n|T��x�~y�/սUw�?H�
    \eyyyBp+,,���U�   B�3�i.Bb,R2��hs^K]�*|Z�s����9-޴X�r ��1.�LMN& -ץm�����}�k      �)�B1�;�֨��e���tO�i����u��� �8ZpT��s��~��^g\�qZ{�Z��_��-�+W�WJ/=w�s:��9U^����U/�����_�.�������bω=ڙ�S]�������T�]�����o��6�u���wl�?��C�}�6�X��$:5��$]��r����i�     ���v�*��k�E�d����   ��f,�b��?s�L]u�U�������ݦ���k���:�9"  z�&v�ϻ����Ʈ�XY����*      ���L(梔A��V���X_�=Z�����?���BV�`�sB�ug]�:F��k�6'{-ڰH���ҡ�C��v�v��G�NӰ�կr ZxU�љ�Z�cY�C1�u�s���b2vd��=��#j�j�ξ!�u��v]=�js���wf`f��ڟ�_م�:QtB�p��	�ޢԳuO���s��͜,    @(�R(���@>�O6�MN�GV���(    ������>�J���J歚�o�}#  ��c���=�`~$�N~���rݹq��y�      h!����[�M�����{{]��6Η��'�*n���j�J������!�{��[�c-8���c���223��EV{=O�G�����q�v}��3-F�1��ϛ̉xw������h��ܪ�    ʬ�1ºFH$!!AN����
�á��h   nu��TTV諽_��,\�P�e,� @�Kr����3es@�p�G�^W�o�Qv����      A�q;�tw�����Z(���w�O;_�gv-`�rM{i����y�<�ю�y<S_��mG�5���U�
J[���g.���[���㤭���*��l�25��sޟ�=9{�ǉ���o     ����X3�QVV&+ ܬ���   �p�.�q�b1���9{5�|�_=_{N�  ����~w�+̹� �����^W�W^dAT      4���/����@л����YpH�V�U���4��YZ�o��h�M ;eцE����S���bo>�����W��>��q��s����Z��mVy��Ŝ��/��Ow~��N����r^��S���}      ���MLLԑ#Gdyyyj߾����U�   Z��i�5k�,M0M)q)��W��T�l~G/�yIK�-���C ����e��X"���3���?������      hHA��Y�q���@H���D�.<���C��/�һ[��#?�i��+������u���{[�SSX����PLC\2vdT�����';?QS�rd�������g��y�FtѠ��Vx���aN|k�[*,+     ���v[&���//#d�b  ������N~�[�v�� �|ڄ���3N��w�c�wC��WJ/3sՠ����^���9��|/��5/+�([   ��j�_S���7���zf�A}xd�      �����ѭh\���M����g��-�GAi�������ٙ���9{u�+W���5C���P��=k|���\36�p�B}��CUVV�����]�h�#�x��D[�n��q^��U�F�?�9�E'Ԕ�����h;�|�&����m�����F���|��8���t���o�돶�������    �)++��ÇUPP��"^?�!�ݮ��h%&&*99�ֿ����P�Ux<��=�f��P��
�h��s���D�>��a��IIIQ\\� �%i�����ٷ?|?���u曆m�v�7��`����m5u�Tsk��C��h�X�����_���o  P��1)�-}� ����;

      hA���F�u�$ �%%*A��~���*�t!4.c��ݠ`�+{����~sK�OհÔ�*]:(�� ��a^/�$���_��VmTEeE����w4��z�js���כ�=K�+ʥ!퇨{�����v+љh^��[�����)�0[��3�@���f,�!=��3   ��(..����a�3SQ�<�_�4N�S]�v�g��.]���+�b�������/� �o'N��ڵk�e��Ϩ��W�^�Ϟ֭[   �x�wr�ɚ����+{x����*|Z�s�����M��=a  �b�N��k�"�# t8���M�+�scA�r�      @�](&�����./�!�,w]�v�^;� +;�HomzKhY�̲��    ����i���Z�l���ʄ�1;�6m2���d]t�EJOOj.11QV��x��TTT��r뜌�r�ʌ~�����UVs����\}��W�fD�.��b�j�J   ���h-��@�{�W�=����rd�歚��׼�Þ�  �)#J���)5�:�u M�ud�~�~���
��     �ނ.��n�&�:�4�YGi}�.m�     @�����+���Ç9Y�!?~\.ԙg���c��f�	�s��3�=//ONV� Y)�����ݫ�^{͌���v�ڥg�}V&L���  �����є�S굏��|���m-X�@�2�qR'  ��	m�j��� �.�{��6g�C+      �GP�bF�ꯑ'7 ���9=.����UžR     ����\�����'�U�V)''GӧO'S.��|�|>_s��'���"�a,�p8���V(������[��=�x�^-^���<?�� V�n�VjD��MII� 4���8�k���K+J�=M{_�X��~N�.TaY�   �Ct+����뻌զ���SxD      @]M(�U�K?�:^ `H�r��c�x��     eeeZ�p!��F������_�&M�fDY�����wE��E||�\���d��{(:r��|�M"1�h�����W��,��Z�(��4SN�QH����������6�����ڗ�������;  P_�v��~�"�# �0���1U��{Fe�M�{      �OP��	;�qG��kw
 N�f�����g�7	      حX�Bǎ�ڵkկ_?u��Y����D(Ɛ��O(&Y)�����P�t�R3T��SYYi>����r:y/  �1�zK���w�Қ��d��*! ��sM����* 8�Stk��8Z���@      @]E(fz����Ť| ����Dm����R�,     ��������_M�/� SF(�*�P����W�˥P�w�^�ٳGh|���Z�f��9�  ��l9�EV/�+_����  hh�\�4%m� ����kr3�.w�      ��j���4�� b�N�"�Rݽ��檛      �h���*++��G�z���[�K��J���<B���J�������[�
M'33�P  @�)�����3_=�uY�  �X���wu�\a'? ������~�n\��<�b      �Ѣg����u[�I� ��	]tQ� ���     ���,�锗�����jӦ�Xbb�������J�+}�7~�4�C�	   uSQY���=��sz{��*��  ���))2^ H�#N?=���v,      P-:3��y��* ���۪��.�Ή      �ĉB�2sB1UKJJ�UX)(�����'�p�\
5��iZ���***Rtt�   Psy�yj�P;�  @S���[�! �����c�6w�      ��j���v�$]��<@M�آtc��ȶ�     lrrr���c^������������
�� TRR���2YEbb�B����4-#�C(  �v�|eDb  @�r�G迺M6_���+n;�=�uO��g��=      `m-2v����K�k�w@397���'�җ�[     L��Ѵx̫g���r������w�PL�x<�
��!�өPbĲ��
5�㞖�&      X׬�#��� �TJT�f��@/��P      @M������3�7�� ��~�u�6��Q��X      ����TEEEB�2N�G��n�%B1FTĈZ��k�R�'11Q��XV��q     ��.1mtI۳ �uY�����&�(8(      �:-.����c u�>�=��'��<��]     No<�5c�����SAA�����`�PLBB�B���2      벅����Kd�	 j����Ku˷��[�      P�����8�ڣ uuq�!���:m�     @K����#//ό��lL�����Ux<B1A�PL��gO��q     ����g)=�� ��:Ǥ��^2To�J �+�2\EEE    �������6-*�'���I�- ����03:u������R      -YNN���וrss���$f�P��iۖI����X���R��gO�      `Mqv���p� ��ft�e��+��`U��g    hP��嵾M�	ń�����83�  ��3.M#[�W���     hɘ��|�ǞPLլ�����������D�~�4��������p   Թ��zm�k�����Z�P��LԜQs���6�_5_  �y��4F��h@}�ڣ4��(=��=      ���P�ؔAJ�e�O �'�/����W&     ��*''Gh<��3B1F ������<�<��IHHP(�����c��III   �1�c���VkцE�k�]ڕ�K��as��7���7c1?���  �G��V�2X �PƵ������#      �i��-R�:� 4���x]��-ؗ!     ���ĉB�౯^DD�bcc-i!l\�	�4���\3��A(  ���8��S5��$�훿���A{s�*XEGD��C�;Gީ�	�  ��].�-,\ �P�O~O1��ܵq�       ZD(��(1"V ��.O���Ց�\     �4^�W�/��q�>��v�-�����Cyy����e�CN�S��HV���  �/������~6�gzsÛz����f���833g��Ƨ
  X��^��M ������c���*      ��,�i�tkr�a����Џ;^��߽.     ��&77W���B��d��1B1{�6�j�D��������D�"Y͋�  �j�a�:`������ۖ�ٯ�ՒmK��%�ۦ��v�f�9ی�   밇���N	 �u�/����l���      ��X>3��h�t h,�%�ћY� K      -	���e��o�z����P�x<�� a�PLBB�B?{��?  ��UTVT�;���k���;�W���yA�r���#�u��+�@��Ϯ�m�>�  @��f�� * 4��(����C+      �'K�b:ƴ����
 �1ihF�t���     hI�P	����UAA���Xѻ*������***RLL�в�i^�J�?�  �-�8WC���/}ZC;��i�4�����mˑ-zc�ze�+�~l����Ԙ�1�:`�.�{��"k�Z��8<����j�  @�q��ue�� ������#�TVQ.      �K�bfu�0��'��w���zƵ�6�~     �������PLլ�1�B1-���E��y�������f�	   ԭ޿Zß�ϾQ�}X������[�_x���9�Fn�P�d~�/�|�²B5��p�K�]Gjt�h��>FQ��߾��B�W��]K�ұ�c  MkBۡJv� ����m�譃_	      8Ų��N1)��K �Tfv�{6-     @K������t��Q,))IVaFRSS������*\.�BIee�*A󩨨0��Y)�  М|>=���zc�f,��3�U�-�F��6���u��}��f�7���Fm8�A[�lQ���A�g'w'�O�on������*9&�N�2�6�|��}  M/����v� �ʕ��ӿ��Q��L      �����k;�Q�� h*������6��     @K`DJмx�%�ө����+f\-_^^��"�b*+c"zs3Bq��b   ��h�Qݰ���?���Դ��^��q�s:�cn�x+��}b���?w��߃��xL~I�|�>��(��H{��"�d��M\��o�v�vj��ތĸ���\��N���^-ٺD  ��LJ=K��X@SqE�hB�P�q`�       �%C1=��t����S|��.�/�-+�xʋ�T�(��=�e�U�T�|�^Q^�<|�6�p��",9�����w�m��0{�3��6&���e�Nt;b������fv�;7�     ��UVV*77Wh^�������VVVVs�y<���󘐐�PB���K�.  ��vߡ�^�G3�Cc���k��OF�%=9�ܚӖ#[����o�� ��m���i#���2��DyA��[�]�-�*��.�,?R��ey}���u��+�l��
��>[xxDEX;��v���=,�m����fK��;��G8���1��8���5��9z��*�J      X23��(!ty+}�_t�s�8w��[���[���2����.m��^g=>��#��8��c�N��������f;���������T�ӧ��V�@A���c�i�o��>�Ev�&����V� 	K��"�Yd�d�$��m�~�3��*$�����s������dH8w���;��~�:'�k^6+�>���b���wJt���//&w
     ���PB�\��h��X%�L&��*����K('!�e�{   �mk�V��΋eA���W�eg^&a_X�Ov�D���^{�@  �igI��X�)0ujc���P�/?�k��y1].��(���\�q�˻��h�'����,��ϛJ\�9R�(2�����ϒ���"      ��b��dE��sTkUٓ;��;z�C�콅b��w}a��S!���G��ݨ��ޟ�xከ���3�h~S炸�yr�BC��s�      �c��5M���Tʐ94�T*2::*V���i��X�  ���1�C����7��\����U����\��L!#��t�\��k�  `~��i���凋�3/,��KW�w�sw�Z��W>�
�7�}�����	�n�G~wns�i��_�jt����X-	      ��r��O�8[`�jY�H���=���R��w]��M��o����؍�Jww�����O��cW��2���D@`k�Gȼ�Nٕ      �b��5�r��5
	��P�J:��Z�&V���i��X����a	��8`8 `6�����c��������z���3W�%g\"�:�S�n���l=��i������?�v=  �����$�k؛:��st �+3��p9}��k7>!r���������W�̵矓D�0�����M����fX���mц��      �f�PL�?"�/ؓ:p�=�;�c���C��?�]9��������w߾�e߸��]��_,��Y�5���r���ϖ����     ���$n��Äb��*��d2)hlVZ�NŨ�̧������ `��p�4�7A2
 s��~ijz���[��an/��P�~��/��.���a�Ȓ����l�%[��#o>"m{Hx�ٟl�aT  8��o||�{��[*��޿q�8�w�y�a*w\�ȓc7�*���+;��>1:�C�վ>1��䡾�&ֈ�     ��
�\<�,�<{�Tr���=��d��Wm�(~��!��l�����]�Y�<�����r^��r��Gd���    �51Y�:Ժ�>}��Ȭ�)�˒���4�t:-V���i��YC�T�l6+���  ��˕rr�+�կ�Ү�r���e嬕��¶�S������<��9yrד���'�P.  hg�.���6���ky9�{מу�v��7H�{;p�1���7�����/.�̞�s[j��ӌP���X,Om      8�e���<����}($K���@-uŷ��x@l����G�n�R]/���f���uyl��~�O��T��c�Δ;vo      +b��u�.�M�^��X,�}W$�L�i`j�YE4')
���AE��   L�W�_�_���|�r���'ssen|��k�'a_X"���Ai4K�R�L!#�B�ٟ�/��vׯ��v�+�����  ���8[`�J��5�{�|���W��[�<x��͍���4-�z����s[�aΊj��y6�      ��L(��]+��4���p��#;n}i ���ݛ�� ��ݨj"�}���6/�q���R_o|�Z)�����@H      �FM�5��D"!���f�I�R���%hL�tZ�"�������>f͚% `�Z�& �SM�ow���lޱ�~  ε�y�,��4�ty��BrǏe����?: p�U��:vsޟ�ta�O���&���6�Ė��-�#      p&K�,<.�\<�,Ac;TL�6��]��k�w�g�iaMp�6�8vsڟ]��Ýw�[�D=�јT������O     ���r9���k �3>V	�X)4��S���F��$�b����lW�x��Ć��� �}��{�wO��;�oF(  @�Č��-_-�~:���ʡ?������߷��x`�����M��������<�b�j��O۾+      p&K�bV�IG &hL�JI�~}˛����_�0�R�ܹv�c7']zÇ.Z�<��%��킆��i�����x     �R�n-���Q�+�Rhg��$
��Ų� ���Omm��4�}�֪  `q��ݶDИ�{���v����{w�ѭ������৯�`���+�OusRԆ�[�K���"�EN�      �D��\ԵBИ^J���Fn�ŷ_����p���4vӱ�Ə��{ZO��V�#h(3B��,2G~��-      V��pkI��R.����!wˊ��b)B1�*��*�g��bY�     �xt,�����h���Co~���=�m�;�u��7�nN��u������	w4	����ǶQ��yB      �<��Zo�Gde|���3է���u���K�1]����ޒ������j=�,���Ý+�      KX�:#�������,�H�$�IAcR��L&#V�F�i�X�8      c�\.�P���R����m�葋�w?\�
��]��i�;�i[�����4u��{z~,��      ���Ṗ:O��兑�o�����ݫ�/��\�����{���#W�Vb�u큨�?��9�K�Ɲ$S�	     �09�z��UB1�TJИ��T�U��x<.NC(�Z�٬
	     ��wJt���
ǎl�š7w�U���ms���f�?�>���؂�4M�´`\N�͓Gv
      ���P�K(�7��J����+7���?\+���Vo�9}K凋}���/\"�<��+�8U~���      X����url�HD�^���eS����e�u���I��V�z`-*R���%      �z�:C�*��<;��������4*����n|bG�y�+��󾎥��uy�wQ�
B1      dj(��	�p�@�F�+۟~6���Z��s�����?�7vs��7~�t�rE��Xۇ;W�     ��&��ZX'��r�$����M��bQ����AAc�R(&������H�VX�      cD�a9;�� �p1]�r��+o^��:�q�ܽ��Y�������e7��-�b,Nm�"���J4�      ���P������m��[�~��`J]���Wf����e?����5��SNl�)��=     `�R�$���fhhHpl�D��P���#�bO2��P�#'agM�      c��y��ܦ��8���%�=�ƹw�ѭ�)��;����hY����̄��Զ��������      8�iG�[�!Y�X$��r�"��z�]��s�՛6Ԯ�,:%�����3Z����     f�Z�&�&돏U�*8���!h,�tZ�"����}���     `�v�&��g��غ��s�ݟߜ��ᾳ2cdh��3�NX�      �1-sv�I�uy֔�j��^���>��	w����|�����p��U��K��޶�r��R�U     �,L
�&Q��%8�D�'��Rp�J��
����B!qbX�488(      �Z3Cm���K`M곘������������!�S�������;�����X���m��p��=(      p�B1�-X�`1Uy��/>q�ڇ(������ϺO>򾶓?(����IN�Γ���      �0Yߚ��r=b�FG���
���Xe��b1q"e��z     �z�3�ݪ�ղ<r��_�ƕ���V�z��>^�����;���6m

�✶���      �`�Q��/,�F�	��P1U~��/.�c�ÏL��?_~�����<�]�ه�F} H(     ��P�u�uC(��Z[[�
R�bR�P�i��XS2���ʼ^&f      L������B�$���7�~�_�P��������-���;� w�y�)�b      ĔQ��V�q���[*lz��o�����T�v���vK-w~�i�q�Z���[����r�"      fX�Z7��I?��x<R��{|-�NK�V�L&#V���I�c?22"��nT,�*.     �F7;�.s�:�2Z��xi�-k�Q`���n���F)^�qڍaO�X���
�շ_{�      �gJ(�Һ��GJO��r�7���E�%����}i�)_ر��.�8�UD�a9-6_�~S      �044$�&�ͱ��n�F��?VD/��訔�e��H$"N�J�,���T��P     ��x_��k)TJ������e�"1q��7�n�/�8���;� w9�m�|+��      ����b�f99:G`��Teˁ��������_�ߗ�oqG/�8�����     f��j�L&�4D(f\���U:�4+m��s�I�ضY�     `꼷u��:�Ւ<|��knZ�����|�Cw�nt�?�q�MA�_`�S��=�b      �@{(�춓��r�a���>z��q�#O
,��.������$��v�K�����=R�U     @����T�?&�r���sϭ����p8,�@@<�1��T�V��ǡP(H.��r�|Կ��+�����_L��D"!;v�0�>��y)���3x�QX)����IԾG�U�V��+G�^����|��~H��Q���P�������۷~����      �on�Cf���P�Uec�����5�.���Vo��{�g�E]+����K�j�yM��+;       �7�U�EkP��͇�^qǚ�X�W�|�����X�X�L`�foH�Df�/��     @']����y���577������k	�0Y|Z[[�
�ɤ��3�Q�R)�
��btF�N8���ZZZ���THFG(�H     ��X�X,�������<�-���V��w���s/�\~��V��     p ����+'G�
�W�lx�_o^��:ACغ��"�ٻwitv��tg�O      ��5|��F��7:
�f����$8�x<.V�N�	�4��� ֯N�k����,��]�B1      Sce|���:��3���{�@�����i�m��Ӻd��tg�m˾��c     ��iŜ�+!�}x6�'��������a��^_����B��D@`�3���ݏ     �N�b&GW(F&s�DB� �L
��ȈXA,�a�39�PH�r�~�V����      LN��%�Y��;�����
ʖ�������'������li�%[�      �Kk(��u+x%��?��E"���?/�/xm��=c�!O��&��V��q[     �j2�v��Ũ��̙3G���A60S*�4�t��b�Ѩ8��}��B1����r����D" :}:�i���j��^�g��<gzϔ�>����.7n   #,�.��#0סb��ux�{7wo.�Zg�����oy�#�	L�q���|���      �����1[~��rvߪ;�o�
�mWo��1|�G�����4j"ˊ�	�q��     �����`���:]A�F��z�����P�U�#��E�>*t�$�\N�y=g�[������b�h��Ծ�P �®��k�����. ����ma�������  �8��|�jI6���w]��MAC���6�
]���G�����c&�M#     `o�B1����
�	�S�U噑mWܹf�>AC���^�yG��|2e"�"     t�!�[(&�7��P��$	��)��G0>VY_�hT�DW�L�[(FQ?��P�ZOs��      LΊ�	sm9��wo[��{��v��~�>vk��>�~��L�2��~R�Z�&      �'m����Es���+o��;����w��B��@�/0���q��&`���Γ����7~&����j�v�eChÄ��2�2Y=g�<��3R(&�o�=��%�eB���������'^zBj2��z�=��O&�o>�����"����w��y>�����%�K��)�ܶ�&��W}��/��    8�L&�e��b�P����߯���
��޽����L&�!��I�T+����$:�Wv��(*��1$R     0ys��pV �j^K�;��w��|_��½������ޓZfw
L��ȜP��=       �'m��Ӣ��ّ�K����Ʒ��x t�w���W�s�����!9�y����`�x�.�GZ�.��m��W_^��bub��Ү��l��E-/Z�N�LCՉ��X-���I�:���2��\���Z^�    8]�������v�	��ZB1###�c�Bl#�J	���U,'��1�ɲc(&
iY��� ����qG�n����h��D"�ܾ�.�  �)wZl��<�R��ud����^�Ym����z��?+��R�/� w�,۶�     �/m���"��(U���?^߽Q�醡ͭk7�6m]�����x��K#�	�      -tMW�<�؍��#��d�A��/8�D"a�]�\.'�RI|>���ŘGg�D��FWl�P 34�4I�o~�o�
 s��w���y��  0��8P��'ï�t�U��*��ۯ��r�-�uu��\`��ƶm?�}Z      `OZB1ӂ	I�[�xj�M���x���ި�~hAaZoG �l��2[�/O	     ��tMoi���P(�e9�ZM������Spd���b*@b���#K&�bj;�&�:�ڞ��v�m���3�     ���Z8�Y^K�;���p��������n�����|hf�e�9      ���9)�t�����/��w.�|(~C�?���U��F9�     �C�d���f�#�?��c{��Û�PLcH��b�hT�FW����I\.�؍�PL>��\.�-�     `����"�
��l��w�{%����4m����Pu���eZ0.}y=�1     @/-���j�f��������Q��ݸ恿_�ͮ5K"��Zq     �s���<�k]5�@ P�e�YS�
�������8ҥT*I&�Ѳ,��{t�b��1c�      `��n�g�_�r������k7>1��O�i]z�@�%�ٌq     �)=�����^I��a���,p���{�paˌG�.�@���9D     ��s�����u�\��U�K$��b�ɤ�����F��$j[V�մ,���Y�Hg(F�/B1      �4�w3ӕ}��%p�����g���#r�Lm�;�      �~�4{�2��]�W�V�W��>-p���nzt��/��X|�@���g�#/
     �Q
���������А�����۷����N��g�PL,'���k�,���J�b����      Lܒ�Y�~:���ߺr��#|��͇�����F�'|    `�2���w�}�T�V'|V?�C1� �k��^ٹ��5�H�(;������R���sRt�      I�d}B1�O��jd�D��`� 	��*�Iō�DgxĮ���U���R��     ��&OP�;z�凋�
���R*V�G��3�����Q?�s��     0>�`�T�M�c|(fa��^�ZEve�.8�ݟt���;���ĉ+��	�K��|�(      F`������x��mdd���<�B1�dR`m�bQ
��XA4'ѹ�k�L��ѹ�      �`A�4q���^J�顫��A_hs��:�����/�vƕm�	�ն]      {1<Ci]��w���M[��w��%+����@u}v�]���      #������tM֯V��J�$���
��+�|b��8���e�=����     `�:z��
/���$p���:5>|�`ܾFZмp�      2<3��K�O�V���_8�]_ڸm��/�L,Z&�F}`H(     E��簾&�3]�E�3B1Gg�P��訔�e�z���d��O(�`0(N�+R�r�l����Q��g      �7/L(F��S��ks����Ժ_qK�ӂ�?hC�zOxJv�v���z�]q   0�*��Zt����v�ev|�,�X$'v�(Mc��y\	{��$�	H����C��7�'�������y�UsՎ�Wj���;�����]�v�ԕ���D���#�n�L�?��I^������8������6����At     ` ]�������t��:�?���T<A�7���i�A��S��%�5xw�dR� ����׆��^m<�ؕ�}�Zg*R���.      86�	z%K�ա�N��p���ڑR�S1_��5�� S+UNI*�X{   !�wqc��/k]V�.m]*K�K$�3�e�JE2�L�$e�T�~��h-*��q��|�o�YEc^u�\?�}�T*=��/~�_p���m�BzmO������]�i��o��[�3M�     #���:���A�It��it*����k�}Pp��.�x<.N�"1�C`��	�BږE(     `|\c�9��z1�s�]_�<"p����Ԝ[[��۾��-ԶNm�jR     `>�91~�,I,��m[����V�U��r����@�A'z��j/�\��Ǿ~�T*=�v��A��343/L8A���H���ʯ�<(������E���@���.q��]��2+2������ߜ�A�5�:v�T+R�U�������x���z����7�SV������]B���y��ӟ����k��c���>3��(d׮]������ۂ���^^8�/o2�#�ˬڬ	����&ٳgϤ&��:YN��0��%��'�3��t���k'����/;]���>Y&��J�U#�L̔�`�/�<���ͫ���73���c������������b���   �Jj�����Css�ؙ����O�S��C1�^_���bb��8��ؕ�C1:����|�     0�C		z�=*��(}I�1���k*m՟{8!�j[7=���y�    �[{��ׂ0��0j^����0L6���aԭ��T�Us�[�=�=����^���Δn��hL����&B1:��ڻ�k��ㅃ���_}O"�������s�%�K��"CŴ8էN���w�{�ԛ�N����M�m�������\���7bp��~�2�;w���m۶I$1t����`P�n~��q�ݻ��M(   eddd����C1�	{N���B#kmm5�.X&D�w�N[�+���}�3�h�d)     Ƹ��Zz_��W>�s����M/�r����Zf�B�d^s'�     ���� ��&�	×[.���_UF�N���j�*Keq��z�'?v-��`�]�7����Ѐ��0��t)�*ҟJ�� o�ܽ�|���'�۶�<��ƶyN�؉zd�]�`o�b����!    Ǧs�~SS�ؙ�P�����r	�,��},"���JȇP�q���Q�Ǆ��     �c��ڙ�E�_�3;p�I-��J����=)�
     8~j,،��(�H�׃0*ctF�?+
��QW5�t*�VG�1�����0c��B�kS�?CC13B�	�)�����K�	�+��#�0vs�@�i��������L&#�թ7�R��e��$    s�����,v�3�~_�f��L��B1V	���%�I���b����-���I��-�`�����t�7     �F6�1�ڤK��h8�/����s�m�+-�0g\Ѐm     ���k�b'ԯ�b�~�u�k�xd5�9����9�(���?W��)]N���݅ݲ;��U�a�ˌAk��b�.���[z���o~�k~���Z4:;ܮo��u�5Q      �kҷ��m۶�K��@@�R�ԃ���S���]3���J$�=��xX%D�wR[��D�Qq�����^��/v����b1:��Q��Ծ      G�`��.�e�m��3��q��qk���sn���"q�"��:�    �Qy�^��2KD����zF�No��e�j|�:9��
�Lu�X+����zfW~W�:X4.�B1큨�]z=:]�Z�d9�O�����ͳ���3`�ُ    ��蚬�&�X�R*�Ď�^��A��rZ���ݬY�G���R��̒J�֤֍���фB����ItE������]�=jߪl�|��(��_�b�   ��СC��A
ٲe� FPg3Qg����n�]��X!'|M`�.Ƹ    P��0���zf^d�,��u;?:_='�T��TF�'S���T��+T�S�=�=�[蕾b_=S���aX(��>۳}��\�q� ��@~�ڱB1t��!     0�����'�؝�P�N�!T�������!��+%�:��qZtC�&tśT�����'TG��!F(   p<���|����x[�n �[�.�$���e*�����x�P��l%��&O�%0T��\���    p�X &3�g����̼�zF}���7^M}F�Q��TGaF+����O����0{�{�@�������X��b&�t�	����6m<��?�����rz ���"     `j�j5B1SL�ϩk�5�D"aj(F����4aR�ڬ w�g^:#W�{��Z���      ���`L\B�B���}���R����g��K��{rt���ԉԶ�'wH     ���?"3�g�um�!b~�i���0���d2R.Om�5W�Io����Ga
{���Gơ�tP��H9}� G�{t`[G v��PoX�ހ���D��v     SK�+��C�#q�d�P(�mY:c�L�b̖J��X��ZA4'��
��:N"e    �ŋ˶m��_��a�?� Fs�14.��P����F���0���2�O��$    h�GZC��l����׷��w�C0ӛ����7�>
�z�pF�N�x��Ҡ�/엞BO=���{�aƅb��:��Y����n�$�Q�'8vC(F��@\v��ŉ:��l2�����R���\w�u�3Z������I�l�rܯ��˗;�L�   �/����~�>0�Ig����c���T(�c��ⴈ��ȕS"e:C1D�    (+W��_ ��w}��7p��z���@�q    ��.�w�|��OJ���? ~�u�3�y�*���������멜��A�z���˯s՜ Gc`(�Y�f�ғ�+�1d�;k��_�\.��:1ٙuf(&�
ϱ����)��T��zA�x81,   �b����9Y_�~�����v�Z[[;B(ƚR�bL�3r��:v��l�b��e�     8:5��;P)���M/
pw�y��󿻼��6�o�"�    ��E�E�k3�>�j��x��Q��a���U�����_����/���`}��Dv@-�k�P!�� �p��y�w���qm�x�m�x�8�����d   �[�L=��#>�OJ�����BWW������wA���zŘ�}�1B���P���     @#J������P1N�F���#s�����    ��*�1\�|�����j�:%�PA�����[蕾b��ߺU��jmj�(��b"���x�������Ю��ĉCE�l� �x�P   ���k������%N�~���Q�P��E��z��R��vFFF�c�P�z�:	�c��Yՙm��l��      ��Z|7�a��~F�q,��se��PQ�}     )���qT�"0�+�K�x=s�*����A�C�C2P��aTf�̉���!���#a�sv��X-Ir���a��ya�P��"^�a*�xh�b   �_7<���'M�W���tZ˲t���b14�>�z>`�T8(�͚}7$
9�x�:[���]��^��ia9:�Gj�C(��\��$    {!��G�4�#�!]�o���Cq2T    �ݨ��v8��VA����M�BFb�ظ���ZI��d=�W쫇`TF�y�4$ձ`&CF_F|aG�}�,}������E�![��x��SC�1��9��b   �_�+�>ٹs�̚5K�:�,�+?ذa��r9m�Ե]<75�J�֢�=V8.���N�3n�֯��,Y�D�-[��   �cIDAT&v���'O>���J%m�T�q�̙ FjK�I[�M������\*x�����K�Z�.   �-B(�p�ZU�J��è��`MjDi�6	     �BE`�x+}Q����χC0���B-�0�JRR唌�G޺�����åa�V�?�p4Ƅb�kq(��/�8e���j���D��ř&�^�H�(�b   ���b&��&�?8Y�t�L�>]�R���Ȉ��:�����U�o7oƟ����n����F��$:�V�5���H$l���x<ڣaD�      �,�	�_)���a> ��|�ʍ��βRg0��H    �����=���H���d>)�BF*�ʔ/g��v9X>(��Q���PL��H�G�	0N�y��}��)�V�!�{��� B1   ��0c��݃j�~KK�� ���'���|�d2�D�`�P���M�̈[�b1�33�CD�  @#R���3�+  �Q�.�4y�d��|� p���ƺ�i��3���&w�u     ����s�+��1$%��E�VxM�	.f2��{��6ۿ���� �G(   �L�7��u(��d}���K��h���w����X�UB1vh�&3�Vv����~	�B���-�P  hD.�K|>�̛7OJ���޽��  `ʵxC���X�rn� 0����!c �;�����     ��g���P��J�%& Y=8vc��>&ja�7��8K � �k   0g��SB1{��ն<���
����
��
���I���'l����:�@�
�Ř�����s�D��ۆ�
 s555����eƂr�����#)UJR�  �xE�!����n& S.��Y.0T�&     `��b���x�j�& [����,&��o�U�U�n��~��B�    ��鞬����vgF�AM�'stj��M����� c�p8,>�O�.�K���e2)���l `��<.�tH XDG�C.=�R9�����O|]ny�  8^!o@`�|�� P�^����P!�@      �0$�s�ů(VK��m�%�䫥}Cy\nq�]�5�& 0Y�`�P    �'�B!GL(�D"ڗiF���x��z�hddĴ��J��a���NQ�T$�Lj]�SB<fE�:;;  ��͉ϑ����5�F�}˿׃1�r^   &�'��JR$�	)Vʯ�u�     �cB1n -]�U������Sы�b���g�`��=)	   �"�q����9�d}["�05���b��ᔀ�a����x�SB1fD��   ���]�|�/�W�����M�'   ��0�]�bMv0�jy��p��     �CB1����-�LP�Z�'0�O�b�$���G�b    �+�˒�d�.�)����9uG�
��ܹӴ�R)�5�c������)����V9e�c�s�}  ��r�,�lc,  ��ː������M&�]�����<      � Ӡ��b^�	*��{��{��� `��    "����'<E"q�h4*.�K���d��1;�A(�:��T�U��F}{�$jߣ�Sc3�8f�O   #���ox���_�l1+   ��u��*V˲����`r���ؽg��M��H<�      �aȑ��P��ʵjI�	rWj�t��#|�8�8�<�b    s�"fLb7��땦�&�d2ږy8��582�C1*N�z��D{�~N�fFX�)�3�8D�  ����)��s�lޱY `���yٲe���}���ŋ k#�`�R�ĠOLJ�V���ˇ4��      �aL(�H��V�e&�䩎
��SˌP��������իWp�-Zd��53�-�b    s&�;)���:C1�r�!�D"�#kmm5u��j���hii�K�^��������8�1�B�P(h[��%   ��/���u����(�������޽{��bV�ZE(h �q7^�Z%�I)�*���qBh      �0�f�%�`����$�<�]osDo|*�a��3�8C��e�	��b    &�M�bzzz�.SM؏�9*u<F�1#|X*�"cj=X��Z���=v
��h[��ȈT*�x��  4�]C���{.�Ƿ?.   S���N�U�B(�R���1'C     �C�����0XM8�	�U�%���.�`�91�9�    oEEtsR(ƌ�U�̙#82��/MMM�ɘw��d2)3f���*�'EL�qX���P($�@@�B�{t�b��j����  h|�ZU�����_�l1+   S�%�q׀A����0`�hn��      �aH(�R���r�H�c�j~W��p�jY0u�`v ΢&��n^�   p4�IM�W�����F�H$LŤ�i���觞���c�N
�)f<���	B1  ��l?�].��Ryb�  `�r�1�Fs��&���p�N���     ؆!��R�H��<�2d���<.O��p%bYS��� �
�2::*   ��߇GFF�.�I1Ō8���O�R���{���|�J��
��p8\��:��(��{�
�,X�@   ��Z��uO^'_��-�!  0��y]B1���Ȑ�8*     �}�!�`8��C(��H��p|� ǏP   �,�LJ������3��q��$3>*c&�������1־L3��f2c_k�z  ����;������   �1��x>�L��Ȑ��     `��F8�d���`���.0����Π��T(   p*3�"N"�1Y�P����I��s�c�VXN�.����D"�$D�   ~]�V�o<���%�%N @��U�NV�Z ���w��~�'�?�_߽�(�8}��w��O`,bY      �aH(����y̞Ƅ��;K`8bYS�P�\�b   �d���ڗ� ���P($�\N�2��|}yj�82�C1�dR`���Q)�͏q;m�Ⱦ�xfD��X�   �sp�\zϥ�y�f �>�O�%�\2����}M�z�)И�D���چ�}�� �T��O���6     �>	�p �x;�!���u{fGm}����P   �lhhH�2͘�n�x<�5��u;c����PL:���b0�yR��X��"&f�{��755�CeŢ�)���6  X�zo���ur�}�H��   �8����!�	py\�+���     `j!�`�&O�����	��}�� ��z��R��*R ��!   '־L�M�W����۫u�j��9:��`(��9�R����h=� s�1�=T�����ږW*�$��Jss�   �m��N��=��-;�  �YJU"	:�|�yL�W<s���      �aL(�Ұ�\c�Z"�r�KFO`��� ���*���c	8�   8��А�e:u��nf�Q"��������d2I(�D�b������L~���r����QԾ�P  0���ݳ�����l1+   f*��" ޥL@���9�A�y>      �aH(&]���.�b0���4��Res�tlW�b �"   '���z���ï@�jD�x��PL:���*���B1���ڗs`�L1#R��=�f�   3��!��s�l���&  `i�xj�
0aw`��p��     �CB1�2�t�'01_�3G^k�� ��"8�   8U6��b��u�jҺ���1#R0<<,8���VS��L&����Y~�_�m�SC1D� ��*�*i��Mқ���] �Y���=(7>x���ny������,�]~\��   �$c<�h�(cB�� ��     ؇!�j�z4yK����"̺7X�P֔"8�����+�rY    '1c2w<'R�ݘ�?>f?'���<Vx��11c�d�6�
����3<gH�f�}�>�>B1�qR�/��^ٽ{�,��{j��e�  p��ՒƮ�O`�x��K�	�{�Ck���      �`H(&Y�
��7/`�Nh�?�q�P͒��>�� �
���y   p3&s;-�p�?��G1UG�H$L]~*��'�L�}�]dߣ�2  `g����^6l� �bQ   �J��l83d�KW0���v�]��z�L���b�;     ��2=U�	����;Z%�^ 0ѧ��ق� �   8���#��8���C]����e�c*����.82�C1V�8����qq3�=1"eژ  Σ�S�{ｲ{�n  �:B1�k�]=O����a_�S��9�%0T�1�      �bH(&W)H�Z����)�o�|���u��78�_p��p�2�, �*j�&   �4fL�v�d}%�j�(j����knn��o��S����\δ���Զ�I���8�1>Lm߼^���em��f�R($ L%����7�ˎ?`$D}���eÆR*�x ���*K�!$��B1�����pi�}      �bX�%U�I��E`�fo�Sc7�Cg0�L`8j�SK*�\�b   �D*"�[<�R������4c7�D"!����,[�b�q)&8�g�H��Z*X�N��/ש��]Q����A��U1���.�����&����n���z��e����iӦ��|5/�]   �[�X�Q_��n�F�cHZ> 0\�ȶ     �N�ŔF	�h�7_(�bp����v�-!0\��LB1���  ��Q֝ʌ����cS	�B1*����$�2#X�n�1Q�$��a�^��__f�b��B1  `����۶m���~��� ���w'pr������VU]���{ $��5��uT�GQpA�g��ܙ�;�2	$( ��@e�fS�%l!���tWU�յ��4����T��T�߷?��,Os��9�O��w T�47t�غľF`L�y�Pq"Y      5�b��̓ݚ�8F��1u	&F�S�����"����S ��   x��s}o���@ �hԻ�o�1�j�L��^��i�q^*��U/�lī������+�2�=  �\���G}T�7o  @���:OGLn�|�¹M�/h���YpzlR}kL��M��     @�X(��$gLihm>�y�o��\���c'8b� w�.��b�}�   �kl,��b�^��H$�F���xm�̈́bƎ+8+������بp8,��q�Jq���{  ��*
Z�l��.]�|>/  �j���<���T��JO	؎x��Ű�bKZ�.�X�     PK*�a"�!P�B�����.`;&4�+T\��Wg��B�Za.4�m�b   �56q{}��	�8���{8���@�H���X߄b�T���|�񸼄s��l��� ��a>3>��ڼ�{X ���5��i�4�]��v�
����"Y      ��b�&��3���"��8�y��5�����#6v�X� �G$^8iP   ^`c7�����7w^71�o��I&�V�'cG&c?ĝH$�%�������㟍��   �~��.˖-�ҥK��  ��+q���ч؁�u�	���     P[*�a"�1�������/=
�J\��������.�e��C 0��p8���A   ^`c����n���8�sG6�ut\j&�C�XL�`P�\����b�p�v��{�s��l�c&Pf���
  0�sb{{�:::  Pk�C}���>*kR����/�7�'�?�T�_9��yGN�o�*�?�>�     �vT�j@�	�i�ă����Y��?�W&ֵ|Fp��Y�D(�Q__O(   �a�!Nk&V2,pz�y��O�.l�����s˖-V�O�����K3k"N���Ǆ������cc��Z���  `G
���-[��K�:�y  �i�S��0Z�,3�?�����O�+�#�6�*o� k{      jM�B1=�~��� ��qu��E(��+�6��0Ep�&B1eE(�QW�gI   x��P����c#c�̎�K&��B16�^��f500`���T����\��q�=�1�Ѩ����0ߜ{�  �1����� ���k��{���~���P�̍	�8cZc�)�azØ�Gp3T     ��S�P����K3��	�73:�ж�6�Q��H��R��8�$: ��   x��K��0����D��1mD���͠A&���N��6�	�؈V��H�י�ӡ�=  `{
���-[��K��O @�{��� �m� s%N��86��E����zJ�_|��y'L�om��k�     jNEC1��6�qHK8|���o��^!�/�5�����U����)� B1   �
�X�韅}>�b���.�;>��8C5���f����W}}����bll�1�s��:�6�=  `[�g���vutt  �KV����)f>�5����ӓ��غ�0W��q     �=A��W�����$8grc�E"�����ysf5M#8"W�km�P>�b �b   �6oG�Qy����6��(�LZ߄K�8�����F��ay��s��c�q�  �
-[�LK�.U>�  �׼��5�N: 6�s�=7t�W�<oιsB��&+8�c     pHQmbq�C��M��Կ|%J��/:y��>y��>�\����~�_pƚ�-ñ�� �   x����,�����f���;���%	��g2�C��)n�x�h����;ہP  x��\�裏���C   ^��o���/_���G��������?�;�q�4*�n1�c���,      �n	���V(�Bs�+��8)�jB�ea�驂�������cS�
�y�w�P^�b �b   �]]]���L(f��h�y�	��	�����;�ېJ���q�2{lls�1��>��  �*�ղe˴t�R���  x[>��]W��1�a��D(%3��/�q��t�     ���pPPeU�k�;�J�)j�qpb�Ig_9���o�w��4�?�%Li�I+{	c�� �   x���ijjR0T.�st\�O�8Q�>�1!!%#���!��n���̹g���`�s���  ����裏���C   x���P�sfE'�~���>������Y�.���}�&��5�     �1>B1N
*W����`&�j�&8#j��'~Pz���fŧ|Fpԛ}L��� F(R ஆ   �y6B1,�����tvv::��׼%	k��T*%8�P��z{{500����x��������<�9�r� �[
���-[�%K�?  �;��ݨcZf�0�a��\VzJ(�æԏ���p�J�q     N)*+8&X�2ϛ��b�v@|�g�l;��m�y3y��}��'׏��$: TN$Q__�   �Ze��a� �B(ƽZZZ��oX��/�d2��O�bl����wĄ��Ѩ��s�2e�  �7�s{{��l�" �N:Ip�c�7N �7tށ��3��蔣~t�CO	����wP|��Qo�r�     ��h��TAY*7�=g��K�'�y����sOikk�w~[pTz�O��,)'��
�����	�   ���8B.�s|\��ƶ�i�66�F�b�c��n���K�E�*s��X,&���oNg8�  ��BA˖-Ӓ%K���W������o�r���B���ԍ���t_�sf���8���l�:     ��'RV�&����y�&�>�̅s������3:G?w�Q�5�z��\���nuuu   j���`���^�ZZZ���J�g�X�����F0$�*`��̹g��Վ�ɹ ����٩�����  ��m�R�P��C��si�>��N=���|T��/^}��ǧ�en��~�ya     �����c����� k��(��S,H��I�±��`�G��+x��7έ;�n�E��^I;{!7 x�   �:��
���؈C���*��*ۗH$��m^���AE"��2����jD=�~��.��e��C( ��U(�l�2-Y�d�9   v�ī�Q�N���4#:���i�g�l�xC����rz��y'     pLQ=�c�j�Vedf|�`x=�FG&��ut�>������ߛ���kB�k����IV,X�bj�P^�R���  @�c��}�����3Fؾd2)��gm�(�N���U��T*e�[��q�s�}6��  j�9Ƿ��k˖-  ��y)��P�ŧM������Y$Լ���cS'�{���     '��!8&�6�t��K�+v[NS"&㼦@�ojc�/JOj��/;i�-{}\p�P!��z��E(���  @�3���X����M��Y�G(fǂ�����p��B1ΰ����׎��{쳱=��߯��z ��W(�l�2-Y�d�9   v��"
6�@����ߟ�6������P�J�q���W����     ��M���v�����([sXr�Ͻ�g^���5k�Q��A�`E�e������ x7B1   �u&�4뿗	���yGǵj�F&�c3���d2��O����������XLx��}�|�0a�  @u3����vm��uv   {��(��00�
Κ���0g\���焚5gl��)��q3T     `���{�۳�檁�*5�����
����6�����3������Y��w��i�1K���*��� x7B1   �u6b!�x\x������tww;:��HP5J&�Z���<�g�a;{)c�=6�`M�	�0�bs�q��0�;�  P�:;;u�]w�P(   {Ƅ����~�ɂ�m���[�����,j��W�z�1�f��`�9��c     �c|�N'z;�Y�A��!��Y�Y�I��L�{ڸ��KO?&Ԕ�,8=vĨ����a�K��B���n�b   P�������^
"���&�b�ɄblI�qD*���-x*bb#Pfp�y�`0���F���8:.�  �_GG�  �2z9��P�%�:��Uz:Q�9�'&����V��5�     �y�b�v(�����*B1�2����?�c7~��_	5c�����G���b����@(����~��ae�Y   ���܆x<.������XC���qC��2���o�S�E���s�ys�q:ù     �^H��3''�q@|�o\�����+��P��X��E�ǧ��1�6      Gd��x�z+�+m�
��_ڵ�It�"���5�����ы/hw��ST�W�>��j��P��W3��ʏP���D�   �&�Z�m#��v6�Iww�������}6C1n�ԺB��x(c[�1�q�ihhP0�˜{֮]��6BA jSSC���Tk����](RSS��v&���$  ��e�75T�)���-'��w~z~��7|��'�����'s|�~�	֘c��c     ���b��֌vA���@/�W�??��@D�crCk��񏔞!T��/�7����k��	{�t�& �3̅�,�  @-��X�|�61F���H���R)�!�j`s���i�������э��
����N��H$���)��P{���UWW�Z���^&6Z�￝��F  T�@>�ҫth����@�oN�޿ɴ%Z�-�nbU�����uoc����0�v��     pؐ�	�y+�ӛ�(W��O��::9K����>�_��#�_p��/T��ms����x"���ZҵB��C ��/v  �7�X�m#�Rl,�7L,�P̎���	y���:>v���,�+�1�EL8�����b�L�\N� w�     x��q ��f4��m���X��QB՚\�،Ʊ1�*n�
     ,ȩYkǼu`Q+�@�y����X���tҘ/X�m���#T�&�}|Vt�(��L�_�{�U
� �P   j������(ngk�����	y��&����"T�B1^:.
+ۼ�s�6��.f�ݜ{Z[[     ����¹�>(�utb֑-��\p����s�5�/sS[�:B1     ���jSNp�[���V*P���e����ߑ�f�1p�Ќ�����*��k>z��-�)��Ү* 8�P   j�֭[�����ņC�Nlm��ȄZ֮�s��T*E(���8���[�|��q���~��=s�!`Ouv�_��5]YB�p��|�6l��  P)��:�y�[�#ޙ+t����=�}Wg�х��J��.���F���.s,3�4      ��)8�P��[�REg�ߞt������M�o����B��������w��g����/f��t��$�dp?B1   �E�\N�L��q�	�lS P4u<ZA(fd�����2�enؾ^��tu�Y�ιg�l�{�{ �ÿ���I�jU��-O����   �k���tƸ���QOn=������7]���}���r�b��	�qsg     `EQ+G�������J���5B1.�w��D*ۻt����j_^p�}�Mu��`���,�Z!TF�P �5B1   �Ef���Xj,�̈́��V؊6T��A'/qC(����4[�B1����Р��>G���     �~&�@(��h�����5�i�|��͂k�s��GG�z�%
�`�W      �qػ'�ސ��';_�'&#��aɽg�ˏ����~���W���|౭�?5�Wx�g���=Be�X ���   ��Z�� ®2!�իW;:��� ���,�H2��6v*�*���x<.��!�}f�8���     �͞�~]�����;Lm��_Ⱦ4�p���sѮ��pn�A�I/Onhm\��̱     �q>�)8�ݡG*=/gVk�`J�#޹���k������{��ˋO\��<n�q�f?=�.\㱎 p����Y4IL
   ���"m�o��X��Аzzz�F���qCȤ��޾f��K�E�����l�9��_���1m�      �l�0���^��Q�0;:iT�PX�x���tN����/8=rX��WfE'�\��̱     �qEgZ%x�;��^��n���';_�ߌ?Zp�G������;>)��YW͛v\r�����(�����P9D  l�Y�UWW���~   ���"m�P�,�ǶيE�}�P̎566�\80��u�iB1c�M(ɦ���B�i��8�؈pU��������s     �;̍	Ÿ���)�r��W�l;s��m���u��"<'���A�iW�f�     ���Bb���	��̩A���9e�A�_x�{���$��s����-��L�Ū�y!��:��r� �B1   �5[�nu|L�P��&O�,�X"�І�PL�HL>���=���Kl�b���w��s�yߥR)k�=      �Z��5�����qp���!ߪU����Ӌ�e�ޢ3�m:�)�ʁ��Db\�??�%]+     `�*]���wB1�,��ո�J�瞵�<��������?����w���+�^x��'$|b\]",��c[��-&   ���Y�c����}�%�I+����>�r9�A��2�Qn/M�'�u���͜{v�湇�     ིŜ��zU'�(��~�)c�>ߊ�N���[�;7����<::��}��F�󇭯*[     �/�{��+կok���]�A�Ţ�xQ��x��>Ǎ������s��Z�u�umw�	�9wѼ���r��p�.T(�d��Be�s l�   ���oww��� |���|>���[�r=�H�P�-�t����*��	/mkb���}��c���M�&      ��c[^$�R�c�[��UMN>�Ƌ�^}���f1z����S�K=��z,     `�����(jY��f�P�{�i�kf��s�;��X#T���|�Ni=�@�Op��S+Օ�*�P��!  �Zb��|��q�	��P0Tcc�zz��"32�bj�ٮ�5���D"!l������%      �ߒ���'ׯ�`��>��65����������o������>pBr����%+���\��     ��'
����M(�;1�k�뵾���sa�[���l
�/\�����*��?��sG����/ �W;�u ��P   j�����87��� �N6C-&���d2��Om�A����P$��pt\�=      ۖ+��d�+:m̡�;���C���sOdQ���	s��������3l�F�.�d��*�     `E�P��ŘZOљ��Ţ�ߴT�L=Up�	�-uw���"W,8�����+�6όO~���^{	�֟��-/	�W( �B(   ����l���Fk׮ut�����@ ?��X"��6��&�(�N����WN#R�^�ܳq�FG�$     �}�oz�P�˙pɇ�����>�غ�Ƿ��S�(���6��ė�9!���~�_p��6.     �%�Z�������998����?�)')��U��N{ط��t�+NY|A���ӭQ�.���#�g�fb<��oyA��A��LH ���   �%]]]V�%�s��f�7n��}�hT�`P����z�!hR�R����}>��"&6�=�pX������P     �{��^�U��5�q��^f���Q��iZ;���ܛ�����=v���f�F�m?*z���̱��     X�+/8�+�NkU��'���3[�똖ق�O�'g9�tG|A�g~t�}w
���{�=���[��l$�ý�� `{�   ���X�m���ي�}�P̎�y�D"����Ƕ4�U�L����
yg��ƹ�@����N�lV���|6      ؎�6-�W��.�߾��c&ԍz)�(�ݫο�߄�v�5����~/n�N�U��ұ
     ���+������C�����"�[�>2��;��5�r�z��^ܶ8+���r\sb�/���"T������g�  v�E���   �[WW��c�����v�V���>Q��ɤ�P��I-2��t:m�{�R�dppP}}}���L(fDl�{�      l�C���s����/(�_<��?c�a��zC�+7�v�W���]�kN��wx�}�%�ޟ�'V�l1�G6?/      �~/X���뢞�O�q�XڵB��5:��"�փ>����;q�i_��k��Lء�ms���K�xܨ}?S�0{^e�ݸDp�Y  �SWW���   ��V(;gk��֭[��ki���N�RBy�h����"&�bT̈́bF��9ڜ{&N�(      �_&ׯ�oyEs[��	���g���V7/j������{a��_��;69�_Z�Q�HU���9�#�      �??�[�?��דrp�~��u���t֔���2���~|}��o�x���O���GV	���E��!�闚�%T�laH�t,�A$���  @-��������Xdl-ַq�6�D�ʸoGM�A��.�L&c�[��q�V��H����9�      ��o7.!S��&�����F���՟��>,�����}�&�t�ؔqBU�o�R     X������￢�I/*#skLǮܼ�s���s�����t��Y�f��������;#]_���A_��q��'�v`l*�b�b�oyY=�~��b �	�    ���b�fB1#����0q�����$�I+�y+.�}T>�t��� B1���{fDlE�8�      ���7���S�[��|��Y��M�ѨgVv~��X#蜅�&M�kY|x��G���պ�N=�^)      ���y��^�
�����>��7�%���/i�(���*���:�O�^�3G]��}Ն��-�ʃ�^x�����^H��L�W����^  �   �Z�b}�3���P��f�r9��)P��J�x��B1�c�L�����ʸ�gF���~8T��:��5B1      ;f"�w���.��a�:��e��WM�>��������`�Y��=���aɽ>5p��*��uOq�N     `�OO�l���B�E�9�1�\�{B15`T8<e�!�]�z��k?�����_��#��SO��8f�!��$S��zC+z7�� v�P   j����^
"�)��֯_��f^���[�F���D'������cg2�|��I$�
"e�g�=��i�3	���/}�|>՚���B�p3_�+��k��ͼ? �n��>7�$łB���G|ǌ���t���1��Z7�:=�Rp�U�M��xhb�)���@L(��zp�     `UQO
�l�f��C��N~#�{��ԛ: >U�~�뒑��ܮl�3�k��`��Z�L?�ӿ0�~l���)��>��k�k9?9�P��	�B   �����ֶ2���3���������ةTJ(ۡ�/y)�e�����♑2�"�C1===�f�
���]u^�yj.���k�ktK�p���;���kr��.�L   N,�7�է'�(T?J��z���B���~ܺl���o�p���S����N�T7j������õW{�0sL�g     `�]�?�l;Ӥg���ҳ�N~3w�{�PL�I������1TȽq�O&�}�o�U�7vy[[[U��眅�&��7�i�''7��5���jI�
�Y�b ��   Ԃ��.������F����
���7�Q2����6�5��gSS�g�r����mB<&ȃ��.2�1c�      ����O��U�j�	����#4�9��H�����U�}__������L�\8�i���;�G��t�Dn�Z{�
9�z��     ��^��m�V�����`��g��f�޺\k��hR=wL�5!PƦN,=.ݜ������o�l��ݷXU����5���	u���':q|��/{jٝ�$Zb���   �n�V�/��bñ���P��}�%	+�f2�|l�bl��mH�RV�^m�W���H�     ����#�����j���5�ql���l&����n�����wt4,Xܶ8�*pfۙ��־���'�0+:aV4�@���=��yu�     �*����Q��T|�K_w���.��B�i�G��}���fW�m|�c ��w��ڛ���-�ҢS�jD/I��WӸ�u��P��f3�]���� ؙ`�P   �[6�U__�����qa�lm/�X;g+>ab(ۡ/mE���)"e      �v����1����Q�L`��^������־K���o�v�f����[���J��YW͛��]4:���^M�f�C�1��u��X     `ِ��`��W�f���*��9:i������)'�9�(Ծ1��p�a��s�C�r�>���^L�ޛ
�n��+�op����է�4�m2?n|Cr��H2"xί�?��BN  �	�B   ��Y�m#��b�]�b}wkii�2��I-g�d+8d��cK,F�H�j�E�$Uk��D"%����ۙl�K�^E  �^��:�L�r��G�}&�2'1c���o��os��=���o�y8����o<����������|�%=eL8�ϔ��&��6��<]:�c     �eO�*qQ�e��\�]�%�gG�A��}B_�v��-�@H�4Mh)=N,���b�y��7�y ��=��zfh६�����OO�t��mmm����+�6��c���a����x�ဖpt⸺D�!PG���ҹ>ݽ�i�� T�@     ���Z�O(f����?L��I�����#܍t�l>zzz����ٴ����q�V��s�.!R���5�)���444p;sc�h���;3Pp�gt  �m�ٚG	�x�	�Lk�TzZ�S���3~qXa�`wWg6�F&���`n���г���37�Ӿ[^Ͼqn]�7|D�:<6�5MiN$�MTa<���g��     ��
�w�W}���l(Ƹg�3��c�{���,�i��Kjǿ�׆F�t���!ߛ�/d��������|������B�;P�������Hc0j
Գ���?k�T_nP��P��	�   ������f7ntt�\.�L&�X,&l�	Ř�c���x&�ǅ=�J�l�zm�@lE��Ucc��ܗ98�P     �Ƚ�Y��������x^s��_z������o���bA���Bo~`�??8П��T��|���3O�l��}�|��@��>�k�GB�P���L��t�س�g�      �+�q���b~���M,��k�Wg�!`[B��ᦀy������jc��P�����`� ;c��X   �����q���l3�C1��G�����l#��t:���Lp�6/ELlE�x��3�e�Ygg���ci>�W       v�U���L��}+�~~�_�P�����<�(�3�K޲�     ��J]��v������z��lo9췛��S�Uk��Q θ}�c����FF��?L��Ĉ�������[��/�o�}i�   T�������®����>2u�Taǒɤ�P�������rx��x�ƹ�DG�Ѩ�k̹��PL�P~O��*      v���Mzr�+:nԾ '<���^�u�      ��s����;�;|�E��g9l���mk�E3>" ���ٌ~��YyY����ޏ[�̢۲٬�l�R���ܙ���C7�|��ϟ/`g��'��Y�a5�)��ټy�6��̙3]���,4ړṖz?���m����ڵ<�\   @�lݺ��1���XL�5�B16��jd�+W�t|\B1��d�����4����s�����N9殼&�HX�Ą�      ��-kѱ�f�'�� TV����5�     p�p(.��`���|(�x`�s:s�qWg�H �qۚ�4X��� ��	��!����"����Wye!   j���ڈLx)�PN�b��VL!�J	{��v������1�K۸�l���~2c�     `dV�n֣/jn��Jj�xA+{7	     �������
;_p�^��z��l_9,W�׏/��o ��y�[�mZ*��H��D4n�8=����� �����>��n����#'N�ׄB!   �Ȅ
����X��\���kii�2n&��������]]]V��ܳ{lm7[�	     @5�e�#:~�~
��{�/ ��/t���	     �|���#��lQ�(�pm��M�G����	�J��h���6��'�M��O���[KN   ��� ����H$���b�������ia��ގ��8�T[�&�2     �]���S�lxF� ������     ��b�dd���n/�pm��X����{u�_d�>��{%�F�myI�ϫ� �.�GX   �ml-�nnnv]CC��ᰲ٬�����_�����%����8=��J��=c�Sf��K�=��־I�     `�ܲ�w�@끊� �ԓ��OW�     �%��+ł|�*��������ӡ����j=������ �\L���K��%x �T(   P�X�_}̂�����5�ʄ	��3���F���8:n&���"l���6�-�H�+l@��)�h4�@ �|>���ñ     `י�í���g|H PN?Y��ҹ>     �BQ�
�2�P��ӏK��1�[y��H�T���` ����?jy�: �K08�   ���X���Ȏ�P��W�윉}8�1!:��b��I�R��O�l�{��)'j1�m��rCCC���USS�      �k�����{��6� �����tl     p����Ip����ꧥ��ҳFY�1�ҝ�~�OO:Q �����ɪ��0�l `$�]�  �j����y)�Pn����}�ڴ��h͚5���N�	����lz;��������m�F��c#c���     �]W(�Õ���� �õ�cJ�tl     p���J�\e䡘K����E��9���5����kt�����JǓ�ٌ��b �T(   Pm�Ͻ���V��J�lm;B1#�H$����0��'lo?�G��jf�6�H���g3R6i�$     `����=��U��G �'�����v�     �ku��:�v%���"�bC�����}>% �]�:u��?�B(�Hye1   jKOO�������Q�pX�=��ۊ;T�d2ie�T*%�t:mu|[�klE����+�f(      ��7��!�
���	���s����     �"k�F�
��k3ї��Xϗ�$K~ױL'���(��&FrՊ�5T�	�B(�HqGj   T#[�����X��n�B1�C'�.M(�1��S�DB�}���D�      �����m��秜, �?]ծ����     ��Z���:��,��^̢�ˢE�ߣ���T�N� v�}��ӟ��܇P��
�B   ����ׄb������ӣ��!~��	B1�����R��Vt*�	���>J�     `��b��:�e_�h' �+{7�uO
     �E
2��Ү�b��EC�^�Y�,�<��ͫ�W��. ����x��;�0R���   l����KA�Jhjj�$��9:��'���Vkk��}���Ï��~G�M��#����"&�"e�����)#     ���ł������/��� F�X�ZP:v�ܜ     �ʽ�B�W��U���K��&�~��)?j?��, ���ߣ����F  �   T[��m-6�>�oxvvv:>��g�윉!��&����g�{�R@�ֹ�P̞11#�߯B����900���:     `�-�Y7|��'&# �;��^�d�     �U|�\p�]�>]������|W�_�[W|��>ر����'��,���S6 �D(   PmX�_�l�b�s�dR�ׯwt�L&3<�eBB�5oo;��r\4Q��mh�ܳGL$��b���ی9v�X     `��d��:�e���y'\`�l�֭�'      �Y���.���^.�J}[w��3eћ���x���� �ӛЂ�ܭH(���Z�   �n���2���`�$v.�&32&�|>���^555	�&�JY��}�r\4�s�^�ƕdb;6B1��C(     `��t������N �=f�k�V>+      W)������*۷^\��㧫�5'��f6M l����ά�;�bd�� ��@@   @5P����Bs�[��V\����&xB(f�e2v�i�k� ���Tcc����9[�"e      峴{�~��Y}h���m1�s�      p�7�������W�Y}K�˧�eQ�������U���?$ x�Ƿ��G6?/ @�`�   ���EבHDuuu��bV�e����
���T�t:mu|/ųlŦ�	���2     ��p�����4M�% x��}�~��     p��T�r����*[��P�n(�x{��� ��c0��+~-�_�X ����S P>�   PX�_����q���U(���������T+�����b�������     ��`aH���X�:WA_@ `r�t��#      \�K}�Ap�=�4�ne�R��~�����tT�,@�����w�'�/��Y� �"
�  @�`�~u���|��j�:�X4U8V6�ut�4��ݒ�d������"e^�ƕdk;��o      j��=��U�S�	 ��J�sl      p���"���g��6tq��b��V�R?�^�d8* �v��G�,�R ��p�   TB1�̈́H�� 6b�f��uܹD"�M�69:&���c{�y��Ĺ���ڎ�TJ�\N����
      ��?k�Ԝ�tp�t�Ro��u�     �u+�+����W�]�;t��Xzv�,K���w���%��' ޴<�N?[�P=�Ţ `W�X   դ���ʸ�x\�sf���b����־SmZZZŘ�v��P��
y��o�q�28���َ����ܹ���q v��k1����������M>��7 ��Q,}}��;u�!�+l o�����w      \���u��x�J�c�����W�t�\`i�
ݱ�I}j�q�=f��^��rE�����G(��
�B   ��֭[�����,���K؈.��w����G&�v����ݼ11��|���Wb<�f~755YyϘH� #��'����㾉Dn�D<��k�0(  �j�9��^���m֧�!*�A����w�c��      Wڢ�U����G�ҳ��7����5�՜��;�����ІbeՆP�]�Ż$  �:�r9ka��`k[���عd2����tzxN���G�m����+�E���8瞲1�7�!��     T�S���kӧ'�( ��5��魯
     ����T���(V��b���r�B��K��?����4����^q���٭� �}�`9?�   �cB��f�9��ֶd���$	��4���>566
#�JٽCf4��|���T}}���P&��f���%R��&M����ڭ��hI������<E�8����   x�ͫ�^M�uxbo���_�OW�     ��6*�EBU)��W�A]��J�N��s}��MW�%��!�m��nJ�N6�$�:�B|�  @u����|fnhh��f(�̛�|>a��ɤ�q3���]�N���o�^a+2E���lD����N��555iΜ9������?J�F��N:d�>��	   ��ͭy_}놨����p���n]����!     ��O��6�	U�ܷN�V��L���޳A?|�^]��G�vm�������� �*   �6�)[��l6���>b$;a^�`0�\.�踩TJcǎFƄul�ݰ�V��PLy�ڞ�� ���ת!D���V����e�e�����5�B^   ��'ׯ�x�6]yЗᆨ@��s����J��
     ���ԵB�)o(�
-�ź����r��n\��M����w�' �-��,�c ��,    ���k�������1E2����NG�M������^��O6؊�yi;!�Y�|v1qw�s v��`���z��i  ���ѻQ�_���a�O	@m�z��z�g�      \˧o�*
U��+ls�N���7�gv�^܆E��F�Z�ol� �s���ݥ���f^K ��w�  @u`�~m�F���m�a���&Mv�����PL&�F�v(�K-"e��V�,���l�j      �䑎e�'6Qw� Ԗ���Al��      \�a]����T�P�|m�ź���?��bNm/�LW�eM�k��pӪ��hǋB�+
�]��c,   P	�B1,�/�@ 0�����U�d2����TJ9���Vt�i����ss�=�e���H�      g���{��똖�P��Z��W�/      ˩�o
U�2+l��\�]z��\"��ӿ�x����/+j��v����� �Mf�&   �vfa��0����lS��X;g#bc�f�L���^9.ڌK5s�)+Jnhh��8��GS�L      *�X������e��Y�IP�^�Y����*��&     p���J� T�ʄbڔ���?�gw�E6l��{�v]����W�?@�-�Z�+~-�wCP�B��    �3��\.ge�x<.��	��^���qmF�I2�t|LB1#g� m�b|>�b�����1�sO�����P���ޝ��Q�����t�}�!	9!܇ x���/tWD��*�?wQ�x�G�@ �,����E.E��k�oP��}O��L�Ꞟ����WOc4H��1]OU��W�t�g议ꩩ�SD�      ܕ)du������U��d��;���ܠt>#      P�~ �Z�j)�u�.�έ��!K7h�������*��_6o�OV�Ny*��P��a��   x��I�L��"�bv�o3��|>om�����K���F����Ɨ	�l޼��q��      �o ;��,�^��5Vs��ܨ�����k     �ӊ�H?Q��k�=+6�s�+έy�c��hJ]�>3�T���LR�]z��ri�r��7��    ��5�ڼ_6Q�/3Y��UMM��s��1qx7�5e�Y�R)��!�HX����[��X,&�?[�.�      ;:Fzt��蒣>�HU0��@%������j�p�      <�5�����O�^�u���\󛍏*m�'�U �/�K��%�i��	  o�D"   �n``�ʸ---�`Ɨ��Y�&M�$�	$�u?��:��� ��ݐL&������}Ɵ�ǕP     �=/'�k����7=SU�*�B���+o��5     𸌳|^sT|����Z����s�y����T[�D�}k �3��E�\Ge�B�y�g ����+�   ��lM�nmmƟ��Y�Ō����J(f�ĉ®��ɦ EL��T[�k:�V*�"�     `�#=/+
��C�Y!qq ���9�?[�G=��      |�ǚ��BE(��[��l}NE=�܋�Ć�+W�AuUQ�<��L!��/�Q+�6��P��a�   x����A
"��<��P�ʱ���al&�v�ZW�L$��l�b�1�d2�2v+��������1S�L      �닪��˳�/ ���������     �,WF�	���c���wn}KS(4o�m�G�����;rż~��f��X/T.B1 �FUUUi)
   �*�[����Q]]����>6���cB1nK&���l?NA�.�����D����k�=�b      �s˳j���gf�* �r�t��'     �U��R�B�p'c�g��s�Py��Q�h�o��#�֛c��}&�tي����+��F(��2�4͕�   /V:��26����Lط�1���F(fppP["��:~�B1��)+�h4���:�R)��&R     �����j�}l�?�7ܶ�)�v�c     ���~���x[a��,TJ�l�����ǘX̏�߬�)�<C �1���+o��K��G(�ފD"�b   �Y6'W�b1�<LaӦM��K(f��X�mP��fP'
���YA`s�C(�|�ck#þ     �;�{��G���o ����^w�      |!�ejҷ���^(Ƙ�E�@?pn�P��gt�+��{G~\'�, �3Ѧ�V��HL������    ��9����E([!#����4����R���M�dR��PLSS�����u�-��=�񭯯���{�l����6�C      x��Zs���i�=�d��MO�W�     �O���Oh�F������M�DI���)��BV�_r�.<��:��pO���OVܢ���	 ��e�   ����j�0Q����	���q���;�D����j��D|�k�TJ�\����O6�������P��=6�w      ر�:R����f�[ ���M��W��      _�H�P�ܟ];G}C�V^/9���A�b^?^~��?�u���
@����`�o�||�,n^�@e1    ��5����Y�pX(��	�N��y���d2��i���
;f;�����=A���`��5�Ry"�     �-&V��g���G�p�9�������O	     �G�W�
�Ι}�k�.��[�ȣ�ł���R4���@�������t�CB1 ��_  �eL֯L6߁�al&
�~�zW�41B1;788hu���A�P��X��)/[��9vo�=&L      ��[�U��׹����� �Rt����;uO�"     �Ȁ���� T,{�����k��sV�Oˣ
ł~��e
Y�1��0��a]��:��"� {��  ��lE=��_^6���C~cB1nK$�v��tl��N���K������o7��o      �tw�s-du�!���P� �/s��y+o��=�     �3��m*��ٵ_v���hy�	�皻�9կ/����8ڒ�w�\�M�^�>S�OT% ~�D����T�*���q�    �*��jxx���6C&A�FU__����Ƕ򛶶6�ǴB���A��e�h3&��-D�      �3n}I�̰.:�c������g���ӟV
     �g�;n*��P�<����
��s�ӗ����i�e����T4d������F�Yz��Y;���zy���7���e��=�wL� �V8ޫﶆ۔�f   ��L���3ok���V���0Y���$ėw�v(&(�E�1�V�=eUWW���Z��i��H     ��-���/�R?8�P�p6PN}�������"      _)�I��B �/���*��O)�;�{U��{��wtPs�<[-��;O�.��+oU����P( �Vu����   ���z0Y��ZZZ������f��	�B!a����]�v��l�t��żf���'(��M�1��!R     �놻����.�bf5N����y-}o��:�E     ��lQAg�j1y? �1�v���������<nYr����5��Q�Ҕ:�O8��-��5�8/w;W� T�H$"   ��L��&뗟�O.�S2�Tss��s555�����Ȉkc��;g��ijjR8V�
z���<�(/�����v}\��i      �g�2I�~��ׅ�}Ton;T ����5����j$7*      �1q����"�7B1F��hH'����㶤�u�K��{G~\G7�����|����?	��\ �Vu�w��   ۳5Y?
�q��P�a�-B1ckkks5�HpU�]����b1��}��������=�����     �C*�ќe7�˳ޯ�Oz� ����ו���\1/      ����	!P�3�v�
:O�R�LEb�<n07�o��k��A��{&�  ;7�ѥ+n)�ց���/�rEp   �����]`3300��3g
�fB1�6mrm���Aa���2�����2�YM�Æe�������ؓ�}      �L�X(/�m)c�C�c�y��zÃ�ݦ�     �S����Jo�X�~]�8��t�6y\���OWߡW���Yg(Z��Z=�E?\�u�휤o#`_D"��  �7���L�v��(���ߘP����P�Ѩ�Z�d����XLA044�l6kel�=�)�y     🻻�ӆ�]t�G�m����$���7k�`�      |�1e��@�V(Ƙ�����I��ܫ�<����u�G|\k9Q����/��w*S�s�: ��UW{�,   P(488hel&q��fx�V��o���u��~�	�ek{�MP��6#R6�YAbs]���Ӂ(      �ϒ�:�ūt��ӑ���U����S�n�     `,WD���ɛ�k��q���(��8�B���[t�KW�ۇ��7��d�BN?_s���^$`W�Ţ `o��a   ^�Ǖ�筌�d}w��Ԩ��V�t���m� ��ḞP̎��e�h3"�J��6�e"e      �֗I��/�J��q�>:�$Aww�s���sE;��     �*�]*N�
0o�b��Y��P����`vD�Yr��eƻu�
��q���t\?Z�[��0B1 �E$   �5L��Xwuu�>.��wO[[��c��x���%(�E��V�=�hhhP4U&�q}l"e      ��/�����#գsg���*λB��]��=��      |,��>��Z-�wC1��P� �֗��@�/�ߧE�՚}��m��.����P.%  ʭ���oe  L6'S����0���PL*�*-uuu�Ι�BMM�FGG]3�H��L&��mb�A�.�	�>����>.�2     ���@��Z1�I�<�,�0Y@P�Ln�e+�ͩ>     �X�Y>�yzZ<�ϮM�+j���{�#/����/�\��!���p�l$7Z
$�����=Q( {����4�X,
   �
���c����a3a�P�����͘����z6:MMM
��
[!s\�<�p��P���6      S��ꋿ�ǧ�K��~�B��R�s��zV׬�O�b^      ��W5O�	�B1W+��t��t�s�d�H";�9�n�i�ӿ�Ն�*͊�Ra�3ŉ��s� ���je�Y   ^as2��@w��p�®�����I&����贵�)(l�{���[��L&���a544      �!_,膎����z}��3�_�Y@��M�����z     �^Hj�~&�/��1*������׹�N���/j��&}밳4�q��J`~It��'u݆�(�c����"��   x��x�PWW�h�P�[l�b������b1WǳD�2��KP�Y�tZ�T���n�΂�v��P     @�y)�N_\�3�{�:y�1*��Ku��;���9~     0�j�~"`;���4�o���!�t�|fc�W_[|�>1�d}d�;T�
���[�p�Z��(  l�����Y   T>D���Vƶ9y<�l(lň����������Z&�j+`be����om�V�=���x��l�ԩ     @�Χu�[�h`��������N�_fGt�ڻ�P�b     T���|�/���kf�eJ�\�GQ=��;R>�-�t��H��:���&N����yݶ�)]��pi}���< �*&�   �R&��26���e{�>��v(�QL%���:~P��6�Q6�YAD�      �t����U:��������7��.����Q��      *įդ���b�+գ��ңνY������K�轓N(L�Gx����t���0� L�  ��0Y?8����F������{��&����.��P�;lƣZ����H      �-��ܕ��.�z�3�������?�ޥ���	     ��ܬ}^�� `��1j���w:���ν��CE���]�����{�:��`^4Z��ƎG���O�Pd_ ��j��  @eb�~��8OO��Q�d2�\.��Cchjj*=F�r���2�M��bʮ�}��]߮mC(      X�ܿR���C��~�>2��
U	�3㞮E�f�}J�G     P1��I���nQ^�N��L���l����9���Ou�t�+�鴉��s3ޭ�h� �x�w�~���f�^���X,
 �U8   ���f����cn#c���um	�΅B!�b1W�#�a�I$��6�ss��������^�Ǽ�����m�g      ��\h�W��׳}+��?�Y�x�ʡ���5wiEr�      *JH�P���9*���b�yڪ���u�s����_��KK���N;Iѐ���ۚ�.]��n��X/�\� �HD   �W���[�P��l>�bvO[[����x<.���p���%.kk߳-Zw�
�)��(�
      ��$١�t��c����X�Q�-���n�xX�v?�B��R     ����<}���l���5��*��z������;M>��gJ.��~^��q�N��Xn̍覎Gu�g9x��#`<TW���,   *��P���g�1�����	Ÿ�fŋ����c��� ��Y[�8.c��H�ĉ     ��):��(�Ǧ��H��\1�����_oxP#�Q     T��.�}K�n��#��4���A�u��"x�|�g4��+o-c�x�{5�a��r�v����i8��B1 �CP�   ��F�����e{�>��v(fppP��ᜠĳ���6��Af�q7�s�      ۶��>���eƻu�~G	(�g�W誵wkK�ߏ    ��d:ͳ����������!��y1|Q`qb��}�*�{����'k�N���2{�G{_�����t� 7�0�r5   �bttT�T���Lַ��d}�-��:���J$���v�涠�}�D�      ���~�x��zc�,}fƩ:�i���t�C�nx�4�     �BeT��@7�C�5�v�r��/�-�I�H!�\�X�}�����/�'�Q��v��k���k�����5C[���PL6���͛����:Ngg�.\��}�s���1Ƈy�<��#��{���}��cmذAӧOWs�w�{D"   ^�d��!�}mmm��G(�o̱���k�e�h3��1M;l>��{      ��̹�f1���q�m�"`_���M��K     P�҇5_�����f�����t^�9�jUrż��zN���B)��駨-�$`O�_�����2�Y ^���W�6m*{$�0���zH��u�9��SN012��+V�2���V�ZU�Xg�1�pX^S]]�og  �?�b������3I.�s}�D"Q:�
���^V�a~�u�X�a�(f}�gU)�LZEe�Ⱦ'x��     ����|a�?jV�d{j��V����[�ًQ     ��u������	�K�{��ݢ�Y!����Ob[0桞�:c�[��)�PK�A�X�W��kyr� /��/q:;;�e���5�f,X��K��_�"��S˗/��C+W'7�@���4k�,����K��  @0X���Ep����Ǿ�����M���b5�ZUUU�9r+n`�w�c=�XLAg�O�������������� ��l�o      ������?�w�>9�M���S�QF��ꆍb     @`�I9}PW�[�>��������PXw9�TI�3�e�����k���蔓4�~����?�_��l|T˓�x�W~�c�����[���ޫ��}�;�QSS���=��S�7o��٬��!��hŊ:��=5(�   ��?W�2Y�����f�>������\}}�@J�PL)�c��8�������ǎm�w<w}l�}3���      �s��/��Wt\�A��ަ��&��-Iv���O�ɾe*     �xE����I�ш�}T١�Z���&U�&���0�BNt���_�[�Շx���:K�T>�����n�������0�;�������f�ҥ�袋t�%����Q��j�*-X��j$f�B���kזb1^��V]]�og  �&�a����؛���3�	Ÿ�f �K��������9�j����v�}��P�96h�9���      �'�y!����0Y�<�D�<��CUBp��"��iyr�      ��\ͺPsD1�"3k� ޫ����"�Ĺ]qG����������5��][���;��P.% ���۫��.yɺu�t���?�����`���)�����
3	ɬ�f�Uss��oG\�   ^���gmlB1��|�mƉ����p����%`bb<�\����e4창�!     �=�zx�殼U�u<��Oz��?��j�
�a.��p�bݺ�ImN���*     ��
�Ӛ�;��`�b^U�<]���y1]�ܯ���L?}��u����^c"7��D��ֽ݋�L�
�y~`b6e�YmڴI^�|�r]y���7�!���s+W�y��]�VGq�jjj�~/�HD   �mf���(Buu����;l4������b1WǳH�����s[ln��{��P�Y�f͚%      `ot��������M���L8V�t�j�$T�5C[tO�"=�u���i     �K*��Z���Y�B1�Z�?��z��͹w�*�9�~]�C���a�z��7�Mz{������$���uw�s�Js�`�K�P��-h�ƍ��Vz���u�����O���'��s�='�2��9���
��}�p�4���   ��m�'mii���<�l��잶�6W��>6#n��{��<�^e����\�      P9�riݹ���rH�:m�q:u±j���o$7�Gz_փ[_Ғ�     �դ��(���b��Z�/���/�٪pE���5��=ڤ�x|i�\��&_,�O+uϖ��\|�
E����̕��pB��W_�c�9Fp�,�\N��կ�u###���Ԕ)S�~����f�   l��`��]6�&���q30�H$���7���477����)     �x[5�YZ�]���5��g�	:�i��?K;to�"=ֻD�|F      �RQh��K@3c�\C��O�|ݮ�~��D5�/��o6>ZZf4쯓ڏҩ�G4��L�gir��Y�G{_�@fH��ٺ��6����L&�k��V^x�,O?���n�*?0��	&(�Z��   �6��B1v555)+�ϻ>���h)�Y__/����<On�KL�8�̱��!{Ǳ��]d�\D�      P�R����ZTZ��iՉ�G�	G騦�wu����W�p�bmN�	      ��(��5_��YpC1�,�-�@RQ�;/�� ����:�!�贉���G�=�$���8L����Ae��1��l^�xO�`�ҥKu�G
�q�w�/�빳�S3gδ�=�I   �M�����f��]�PH����&Λu�P�����];d)&dBAeb9�B����X0��6�=Ay����w����qv�ޙq��      @�l���ΧKˤژ��vx�<��&�m�Øs�7�z      ����Q����p�j��ڠ�t�fh��2���f�Pgi�j�=:�e�Nl?\o��)u�;2��'��O�+�d�R�e��,*��P̶��䦛nҏ~�#!Lte�����<y�jjj��O(   �ي�---�]&�ck0�N�:U�5�X�n�+c��N&�䈓�H��W45#�Ͼ'�L�ʬ�6^k�lV���jll      �����_�13���;�;Jo��C��($��n(Z1�YX�'z��B1      ���
�s�����Y��ܢ���2��c*�z��,P���8���\�{J��[g��rB�����3�RmI�������j��P^�DB~�x�buuuiҤIB�[�h���L�����P   l3�m	r��+l>6�=?ikksu<B1�B1&`b"�.�J)�N[�P�}fc�f�=�b      `����Z߱U7t<���z�z`������h0"�nId�K@5�?ݷ\�!     �u���>�+EY�cV�ߛ��u��QH�w���W*���]0����+-��j�<C'��1-35�a�¡*a�ų�Z:ء��k�h`U)��Jؐ��522"�1��C=���>[�|�?�������32W�v�   �d~f�����o%c��`�� �w�ۡ*�6m���f�9(���>kc��Ԩ��N�+�������&3}�t      6�F�x��r��t��;Doh�����6v_*����F��X���Wi�H��s}     |�\��ۚ��X¬�Y����[��~��~��>AP��+N�b�TEtp�:�yzi9�Y��99x{&c�0K7hI�C#=4d/344�����O>I(& �-[&?�d2�SCC��c�  �M�����rV���jj�ꈶٌ�،E��ۡ�]�d2iml���(e����lml"e      ��gersi�ɹ_�Ҵ��tT�9�}��v�����^&�UC�ZR:ϽC+���+�     �1�t�F�o�R=,bV��Ջ���)�X�;��3�=l��}5��,����l�_G4O׬�I�퉚Y��µ�t�]���ֺ�n�Jn���FfG�;���j�ƍ��Mcc�P���x����Wf��1�c   [��x[L$&
	v���X������P��P���%bbs��J(�l>6�? �M5Mj��w~�{�յj�oS��e   `G
ł6o--ww=W�ڤ�X風��K�D�"��٬/����9�]Z3�U
�l�      {d��|I�t�  3�92��B��U�j�.a�L,�Jq�����Kᘃ&iz݄����pT~S,՟��T�֏lպ��Rf�s;����)
V�M�R�+��Y�b�N8��r� ��ي�D"   ��u�b1�>�σ	vf2E��;��&�����[?�&	��PNP"&6�=6�X���"e �����Շ�������>���^����   `�����!��ׯ�DJ�X�8�H�\צ��:�����t���w��0k��4��§      ���&�TH��<ٙ@	� ��ݵ@+��'k��PQW8�vKw:^Z��_񚯷F4�6�I���X�|�i-��߹�\]��H���t��ȣ�l� y&���x��{�}���Z���}c�'6��S~�f�B1n�֭�;�P���--   ���w�n&�{CSS�B����f��ĉ�]kkks-388� ��	J(��'(����|`s�      �S";��kJ��µ��N�i-]uR]�纛���R
������s������o��ʏ
      ��a��5��bì�=5O�yz@a}EE]�|�I�+��piY�ܴӿ�\]��H]�sK�ܮ/���T[QuU��i��-��HUu��E��P.]��90n0�H~T�bQ�|��I�K�KK.��_���5q*��w�)���Vhe��z������   ؞�t��d}o0?��X��8���cB17nte� �b�q���!k�e�hs�C����`+Rf�a��i���
      �D����w����ה�mo�4�.����hU�_���{U��ҹ��a�g�*8��_�.�����|�s2��y�۟�n�}     �k֨�ok�n�Q�b��B�����<ݠ*�Ĺ�Ig		�n�t�{D��' �W�BA~�L&����PL>�/MN1�T�T]�[Z   ����oml&�{G,�����	Ÿ��1ǡ���4�؆���y����U�٬�����>s<�����1c5�4i�      ��J�GKKW�^�      �nX!�S�.��x�j��Bmv>~Z��ҋ^z�  c�q�S�P�nttT~gb1n�["��    [�����*x�y.6l�`el�렟��1ǾL�#ђ��H$��m� �y�k���U�H�w����1c)#            �B�+�]�*}Ws�%�Ō�z��x�f�4u�s�� ��I~�(RSS#T�Jx�C���c��   �I�RJ����	�x��p������b1W�d(�f�8(�D�q(s���^���oڴ����{             T��B����-�J>¬��4O8(c
���0/ �g��a�Y'Mcc���Dbl�����  ����Yۼ���D�������vW�3�� J$��J(�f��<�6"��1�=             �W��r���;������rx5�&���ď��o ��X,Z��1���&���=c�*mC$   `��I��g�0�Dϰ9Y?�+�ϳ>�������R)W�j(&�LZ�PL��b1�;ZZZ��ms=            �}����M���|�PL�5O�ݥ!�߹�-�k'
 �f(�����d�}5y�d��M�6M~VSSce\[�   ��$i����z6��B�P��p�y�ŔW"��6vPB16#e��͂w�\�m��             ���
�v�5O�'�Y��6G��J�:���Ug9�Y��+�@2��l�����v�aBe�9s�"���٬�����ʸ�0o�   `��I�A	"��	ńB!k�\-"3���6uvv�}�.� �3�<��������v�f���}���|>L*��p            �eI�ߊh�.S��
��{n��E��O��Xy}Ź����j �HCC���|�S�N*��Xab1�V��ي1����L   ����DA���\b��d���f]�5k��kn�n��|��ӣ�!S^f�2�[Z	�x���ٲm]loo             xL�B���u�.��+�eD(Ɔ�Z�|���ՏT�Ϫ�/8� �͐C]]�jjj4::*�y�ޠ��*���-o�e(ƄZ������KW1   �40`����͂��	��B16�E?ikksm�L&���Z���q�q� l��81�U4-��GFF��o"e�b             xD�YRHרQ�k�2*���������r�Np>������� T(���\9���K~s�i�	�p�I'��o�ߘ	�����Z�  �۲٬������d}�1�ɦM���m&�cln�bL�!���T*ee\�	Bd�v�����}��P             X֥�~����\��b�b�9����m��)��9�r�  ��L�[(Ɯ�����0e�r�!Z�j����Ճ#��FGG   ��LַC%�=6����p3c+�b����M:l�9L����I�����26�             ���^g����G�W�G���2g�^QZ��Q
�,�q����
`s�QWWW:y>�H�/�������]v��y智��K�555֯(�k   n�9Y?
Y�׳�����s1�v���Q�hT�L��c5f��c�#A�g����m��I��>   {+����gv�5���������~�5����g����Ƈ9�k_��&�;mڴ�ޯ��Rmm���^CC��f�����g.hd�5       \SPQO+�[T��5W]��^�PK��f��]4���� >e;cL�4�7�3�C��,'�x�f̘�6�8� ���   �m6'G��חNB��؜���fK�L;g~v5�Swww��"㮠ĳ�e2Ծ
J��ol��6�G   �Oے6E�_T�ºx��;���TJ������9�dG�
��~�6s,"Dts����>��r�Y��X���8�W�l�%;{��}d�0��}m�cG��R���秿������h,��#      �R�t��t�.W� �T�o�oј�5[oSQtn��Y�u~��7��{3i�Ll������	�s��g?�Y]|���:�~ڜ�M5�   ���������b�IB1ckkks%�N�4�x��cA��،�����$�����<�^  �;���z�^��W���ÿo�
��a�Kl�RB=n����}���՞0gA�v��V	       *HZE=�*ݣ�n�e���aF��5OO;���m���*�]
������Lm ���ӧ+�L*��˫=�P�~��B0��Mo�)����~X^eN2�%/�,D(   n�9Y��F��툂Y'�M�&�[�3��f8��Wj�v�f�,(1�����r��1���f            �>X�,���T�{u���K̨��y��|����q�ϤNTH�9�w:_{��4 <�愑�+O��S�ׯ��+��[�"~p�s�/^���>yє)S������V   �6���mI�c�hT����2��x������6ֶXLPd�Ykca�8<<��+I���}�'����C�b             �-��Bz\ݫZ) {���d�r�����Hg)��:\Uz�s�*�]�s� ��]A���]�TJ���򒪪*�w�y�0a�lMMM��w�[���iy���2q�Dy�   �������mO
�Ι��V(�f��O�Ř�GMM���g��KB��v*�	�c�1���֎��rƌ            �]X+���P���PK��ޚp�3j+�-�;��e�����t�Bz�����g�c��@@@M�2E�������3��+_����0f͚���?_�^zii2���Wt���P   �d"1�|���---�7�禳���ض#~�f(&����SP<��V�5�)�1�Jg�5ξǻL�������D�             l'�,��������T�E���`\1�6hj���,���k�T�r:FEg	�h�pLH3��& S+ 'Ţ��P��X�v��X��^���/��SO��������7��y��&�����T�ט��K�   �M�'E�	��X,fm�~B1���.�ϐn�|m�0?G��1�`�u�&��qs(H�ߘ횭P�             �̉C��z�F&
Sp�a-���
@�1��eJ8����Z_�dU��1:���)�W�sn��|n/�~�s� `^��b1����=��������[��V;�w�C��K�J��|���O��H�A(   n�=)�L�7�|nFFF�N�U[K�{W�ϴ�y��+��)���$���V�J<�f����Y�pX�&"e             �I�Y�	�=
�>���|~5c�u�8�_m ���ص�j���,O���}Y��S��SAag�o֭m��lp�u>W9_gP�"U���O��;^�f�Ќ3���X
�
�ƞ6m�.��BM�:U��w�q��+4w�\�Z�ʵq��ì�&L�W�I(&V�jr4�  �8��c�,��csRt]]!�����4i��kmmm��bL�'Hl�m�ϲ��iH�ǯl>?�b��ЦC�|�_ ��������AC��������W�OG
 0�jj�H�Z*       ؑ�rz5 c�J������R
;�S�ӕ _ ���s�K��e� R���+T�#�����Рe˖�=�Dt�Yg�#�H�6�;&O���/�\�^z�+�+FO�>]555�=	ż�o/\��  0�n��!plN�J��l�̺I(fl&� �b�q4[��րDL��;����;[��t)eBv���������W��w��"�}T�M�-��TX}�� @Y���zO����        �P �5�&��)se�P(T�1L�Ƅ>L��S&�b�-�6u�TM�8Q~�'�   `_1Y;��P��V(&�˕*UUU�t�l��ح�d2[�5 1���bV�7��              �f� \�P��������z��b   �&��ۓ��k555� m:��2��u�O�|�XL4U�K�R���v�v�P���z Rv�              ���  ��P.�b   ����!e2k�2Y���s���eel�1	�hoowm,
B(�lm��jnnV���b��muuu�팭�'D�              p3j �!�\�   �-�'C!��w---�B1L��-&z
�\9V�J���2�yl�sY�lG��v�f�k[�n�2v?�2              \ŌZ �k� (sq   ��'C����6��Q"�P.�#�9�3�	_���e*'NT����2nP��6#P&�C(��l�b��             �.� ��P�r���*M����   ʉP�b�92�^L,���]ص��6WB1A	(��X�HP��6�=���ħ|�f���{#              ��3;  P̤%B1   (7�чh4���z��lN�7̄}B1c��b��344� ���I(��loӰ{l��ɤr�A!              \�{  ט�Z@���a   ��d}��v���:�'mmm��322� �d2V�m@(�Dq����[��;�ϓ9�oBz&L              (?B1  ��PN�HD   @�ٌp0Y�b�����d}�ͭP���*�	����V<�z\�}�?�~-��G�b              p�   T��j��  ��FGG522bm|&��C]]��Ѩ2����mƌ�ĭPL:�V��f��ƶfr���SK b<���k�}              �a6- �6�z �   �ܘ���e����+c�^O�bB�PُY��~.���Ym��ᰚ��U�l8���C}}�"���p�              �S�g& <�P�r�&  �2c�>vW,��1�aL;g�
���J&�ektt��fu�1��	�zξ�üL��������b              pO垙 �B� ?���Q>�/�����/J�YW˥��J~RM(   e�d}�.3Yߖ\.W
w��v���͕����`�g�J���ieܠlm8lnϰg�k�V(��{$              ��ٴ  ��GQ����G-`_�y��k�  @�1Y��v��L�'36�ٰaC��I$�<y�*U<�2nk@B16uuu�F��?�|�`��bQ�PH              ���M p�9I ʉP   ���d}�~���Q��Q5�9s��k&���aU2[�AŘc�6#e�XL����|>_�b�$�             �M̦ ��P�r#  �r�9Y���Y�PH���mF��ĭ��Ȉ*�9�g��/�d2�\.gm�V��b�5a�=�3              ��i  P� ��k��c��Ď���?���ۄ@s1�k'ΏK���t(��DT�?Z�R�*jz��q�����J�;��rIU��Q@>(��,���@�c��C�������L�;���@�=3��x���3�̰_�3�<3�|�@#�A�K�.���������fԨ�4+����:U�ĔJ�T��f��ӥ}ꆟq'ɵ@�lǎ         h,Ӵ 4E��� �$ @#�HL��m뷗����g�JC�q�v111єuC�J��[�ZiG��{�Kڏ׬H         4�iZ �B(h4�  )��F7:I�$Ձ��/����P̆���������u�bꯧ�'����N��k9������X��Q,SYƹ         ��4- M!4�P  �4cX���>i�bVVV��A��&&&¹s�����z�҉�[RY7��b�����Φ�~�9�>�D��zϒ��         �E��W�  t����   �277��������v�'��\[|���;2�����ʺ�.	��)�
Ŵ�)K�y���         ��P MQ*�@#���  h��/��~�������[�l	\]�Ph�:��YXXHe�n9&��SZĦ�P�Ǚ����ndd$          �#@S��� �H���� �8i�g2�ԣ#\��Ci>g�I�B1�����F�I+���P���JX^^Nm�\N���Z��#         �e� ��  @���i�э����K���333�kkV(��Q_�|>t��"<W�b�R��=[�n         @㘦���@@����$I  ����|X__Om�l6h?i�7j'�
�P_�p\L�5��iK9�         �xB1 4�P�,}}}  �mff&��s������X���	�b1���~޶�������VWW�#�χN��k8+R֖�~�f�{         ��b h8��Yz{�� ��fggS]_(�=%I���S{���χ��5A�(
�����L1���{���dB�TJe}�         h<��  t�8,  ���гa����b1�;776m��:�����f�!�N��Í�������4��         @�	� �pq0	����  �[�C�1�@{J;���B1�C1��\�LҊL]��Ӿ�c�V(fqq1�������          4�P '4Ko���  �_����E�Di��~|>h�pL\__����2<<hO�5r�̙�֏瞷���         h�� 4�P�,B1  4B���$I���x�=�����	\[�P��\�b�y'�ߩ�xR<�Оr-p��        ��1I@�	� �" @�-//W/i�>���=��f䨝Ŵ�l6:]ڑ�\�x:Yι         :�	 N(h�  ԛa}nFڏ_���v1>>^�<���h}�|>t��_����di?~3�=         �P&ih8��Y�b  �����T���okccc!I��~7277W];�xs���#�����/����=9����)        ��f� ��! @��=�3���zzz���x�t�R*����ڞG�V(�b�@|M� S�s��f��\����CG         ��L��pW��� �!��2�L���ۯ�' @���f��0�PL�ÞGז����J �ӥڈ?g�ו�ҫ������Ce��         ԟIZ �j�������� j�� �P  ������G����3gR[?�bv����B�h}�pL��KM3.�{�^����)�J���*         4�IZ  :�P  �#i��޴��ôcG�"��Z_7Lb`c}}=��c�wtt4���k��ٳ���=B1         �&ih��Wp�!�bs  ��8������!+���[�;j�֗�PL�q�x�I�$��r-p�ٹsg          �O(��*�J�Yb(fmm-  @=�a�4C���á��?����O;:�.�������b�u� �vܩ~�� ��         K(��Js��>}}}B1  ԍa}�!�ͦ�~���v��d����Wk���ӥ�H��E}d�{         �c	�  �1�_ �z���Ku�B�hqX?~V)������������P���kNܠ�e� b���gbb"���~�~        @'��=��S�7��\.�f���� ��I�3�;��@���S�m�N�>�ڿ!�b�b�-��ZW.����N��C=��Y.�K-ز��         ��0I�M۳g�?�l��v�F�a�h�84�$I  �zMm����p��:�{����B1�3���@��&&&�+��v�g�4�=�6m
[�l	t�;�3|�{�Ke��>         h� n�׾��-I����|�4���t3=���[\  �c�Ν�a�Xl����sO	t�ݻw��{.�?��ko޼9�-��ZW.��`׮]�?�a*k:t(�v�{�7<���aaa��k�z�         hS� ܔ���?-��qJ��o��Z��8���� j��P�P  �244�����6u��۷���?�9�g��}�c�_�B���6f˖-�ֵm۶�b(&F6N�>��u����w�+�9�O<���/������#{         @c����MMM}�\.�j��V(&���7� �U<���ᥗ^
�Νk�z1�я~�:dMg��r��ѣ��_�rx��W������>��066
�B���	��P��w"G�	_����ڳgO��>�<1�Ce�<�LXYYiʚ�
         hS� ܐo}�[ٕ��?������7�  ꩿ�?|���X���['�T�����{O��n����O�cǎ�S�N5l��طo_�Ї>�>1���|'�Z�򖷄�[��n#���'�W��p��ņ�300P=��߿?йv��>��O��~����ٳ['F�z�p���          4�� n�����l�\��ҥK�I���������������˕����os�L& j$IR�p���?�������R�~�̙Ϯ���/^�_^ݼy���]�o�PX
  p����ѣG���?������ٺ}��y������j��7::�x���/�g�}6�>}���ݷ��m��Î;�/3�㲼�h>�`5��M6m�>��O��~��azz����x^۽{w�����$:_�}�?����s�=Ν;W��_��s�С�y��          4�P �mjj������~�ӟ>�裏n8� �(�c�L͗�sss~�ǎ  �	qz�޽aϞ=���E��/~��_����I����^����Q��[��]�vU��>�|�;��������<���K��ŋaqq1Fx7�=2�L��4>>����W�ߖ-[7.�F�9�y智|�q1�/�(��b�)��N�:U=�\�p!,,,�˗/o�{V��1s�-��m۶��;wV�7�%����;��W^y%���1�\���2=����T�=�\.l߾=�v�mհ         ��+P ���O?��>_���'|���@��.��ͽ�u�$��رc��c�  p��u����C�P���^h�y�{�=��~������G���n����z��!�����         @{����ʦv���f{{{K��600�7�/_~}z*I�?y������_   p������·���@:b���ѣ��?           ��P 655���������~��d~�T*�@����|���r��ym�����?�l�e   ����B.����7���b�yv��y��          x� 6��ɓ�Q��we_�$����w��� �*��b��t{���?������ϧ���9r���   �w�qGرcG��X��O~�����y������]�v          �7	� �!�������[��P(�MeS�0��R hI��b�jtt�,--�T�O��n�T.�yzzz����>   6dxx8<��ᡇ��b^x�p��Yј:)
��[ow�ygu          �9� ��رc�(�˟���������=5_�@�����
�\�/^|����y���ue��   ����P8p�@�R,���\�+W/���������/          ��� pU�r99~���U�������+۞��	� -!I��CR�}}}}����n���3���;|���   pzzz���D�          �,B1 \����'�$9T�ott��L&so�R�$��r�\�g�{&&&VΟ?�Q�k�*�����z��ş|             �-� �����R*��}�$IGGGw��_���9 ��r��*Ǫ��ձ�u���###�-..�]s�{��}���|              �6 ��*�J��l�����t�$��e������T h�c҉���{+W�*��q����������qm��t�ĉ�<�ȹ               -N(�����㏖��߫����{f``��׾\���O����� �b&''�zzz�@�$_���Uvm�f�5;;�`��Ƌ���+��              Z�P ��ĉW�	����+������J�҇����� Т&''���ɓ�;>>��r������}}}����n��ۣSSS�w�ȑ�              ��	� ����U6[k���L&��r��+�#���g@�;x��J�\~bzz��$I�o����W^y��7��sǏ���Çg              �(� ������͓���$Y�f�o�\����{�� �D�V�l��я~�ROO��^YY����-�r����              �(� ^w�ĉ�R����r9S�?��=[�wjaa�<xp= ��}��}qzz�T6�����qm����?~��_>|��              Z�P �+����yO�L&s~pppjrr�@��˾����}vii��ܔ���?��7��;��              �� j�8I��߰����C�ݻ��'O�|�r��/o�muu5W��     ��rE          B1 ��ȑ#_ ]�������y&  �$�  @�)�J�        �T�    �J�D(  �6�         @*�b    ��+            4�P    ܸb            �&�   �T.��b            h
�    �q�            �@(    nP�"            @�                 �8�                �'                ��b                 Z�P                @��                hqB1                 -N(                ��	�                 �8�                �'                ��b                 Z�P                @��                hqB1                 -N(                ��	�                 �8�                �'                �����3��>    IEND�B`�PK
     )u�[����  �  /   images/7de8bea6-aec6-4ad5-83ac-8e47725efc1f.png�PNG

   IHDR   d   B   �s   	pHYs  �  ���R/   �eXIfII*            (           V       ^   1 
   f   i�    p       �     �     ezgif.com  �       �    �  �    �      �w��  �iTXtXML:com.adobe.xmp     <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="XMP Core 6.0.0">
   <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#">
      <rdf:Description rdf:about=""
            xmlns:tiff="http://ns.adobe.com/tiff/1.0/"
            xmlns:xmp="http://ns.adobe.com/xap/1.0/">
         <tiff:Orientation>1</tiff:Orientation>
         <xmp:CreatorTool>ezgif.com</xmp:CreatorTool>
      </rdf:Description>
   </rdf:RDF>
</x:xmpmeta>
�[n  IDATx��]	�U���{�����F7�Ѐ���*h���$I�$��8T��c�ʤ�d�d��JU&��*Sٜ$f☩%JD�
���4Mw����}_�s޻�nO׭��������g������oy1|����߹���hT�.>����v#iK"�f���!�#���8/�`�9-���UaK�q�aN�aIZv�`��)m�rP�U�9��:a��\v�'�w]!74CQge!�,b�\A7���]w#mM!mNɻI{Yc�0��<�c�,
��a��G��u
�!OIsRڲ�|!.�,D:���}��n����:~�_T�w}�i�O�<�8U�<�ن��۾��˞W��.2���p j`�ۋ�� #����]7�F�9]���n����b��jőA?�m8T3z����`6�7@���5�1���L#�a4�*O�0��|w%B���8Z<��"�OQ�##a$�,�{�	�r�c�8�8*���p�ì��-�� +�#Tv[	G�	wc�~|�u6�_	�ǰ��J�W����{g�)Mt����CX2�6�9��g��4$T���;��;��� Ӯ��Q�U�$1N&��O�c*,�
��13�f��b�F=�^,;M�py��[�٤��r�
M����R�Rw�`	Y`�6"�5��J���E�6��z����
Q]�".��Q�����8�`6�-�h�z�l��v� pu��Ը�%#��eWT]6���I�P/��c�~=�fŘ�h�<�������ճd3�""߫A��|�z�ë��|/���@$q���ɀl.W*'R�w�IR��S��NJ9N"L@��?ǸO���XL�0R���ap+UU!�	�7�~�7�A��zy�လ����C5��C>�O�K%\�^q�g�d�R�W�p��n0L�HB�*XC�e�i�o�1�Buh9g��~�%�V��f�����Nt��겫a%��)�'��z\FQ����K��\����h����x�?B>���Յ�����\�%�b��PSmCo_v���V��rZ�v�I5E����C1TU؉��p��s����%�PW�T:�?������}Ǎ@(�h4��f��cH&�C#Qd2�z00��
8���=S��XE8�u�݌r�E�q�Y�v�1NH�BX]��-��:y
�Ch�)��:�FR��[#U�D�jcƸm�?v����l3�usF�e��q2����ߡ{0ؠ��`����Tfc�7h�2�,HO���20i�h���<�0��dΩȐc@���S�@=�ޑr� >��
_W���yאe)��1#x1��n�Mǋ��sT��u�ڐ#��B��[��b\����qS����+II��\��?�&�A�{��%�ep!E�nfB�:��ݻ�p:�t:�*s��r��U�2g�B�U8]�}��`~��26�|�T��>�0C����W�n��f;�C>�ZB����,�K#�����hA����p=q�����Hw'�,���e�%cApI ���<y\!t��eDx^���q�#�at�w4�&^V7yS9GqG]�e5��G{Y��l��� -I�1K8���0F�H�~�?���,����Ŗ<A����`NY� /�6���g��`C^nQL�aZĳI<��"z�c33��s�Y+�=fv��arYT�V����"���G���Ov���H�6m��l6��3��'؀_�]$���`���ǉ��F��R9RF���cu�jx^8MN$������*W.&&g0�2�2��~��w��RC�D�r��X�gj�>������K�c�X�]f"���.��o�\��
eG�T��x���k�rw����%�"�3b��n�%k9��Ʉ��r��ԉ�iR�Ia���COOrd�X���4!~04����Kh�^����X�X2&��,0j�N�+�_9_Ž�S�~
���Y�U�a$8�zo=�c�r�����D$U�O|��1�yꤧ��qy��Bv&�B8���D:��g]��^x�^�3q�n��>dHO���kE�������
�'�b:�:��WͿ
ۻ�#j�N�m4100�w�yG~3�-�v;���p饗J�����:U���3��1���R��'��	p�-�-XZ���c�zہ�Hf����BrG��i`È���R1D�Q!�4�t���ف֊Va �J�D���jTQ�G�5���ar�33wU�@�܁XJ�i�{�|��֭�33�I�^�3�TJ�Sq�	��$(�F�.fÖ�[P��Қ��ӻ/xQ\B�نFw#C��uբ?�/�r#���t��v!~�X.��@�"���W,C�x�0��l"3l42�D&1{f�"���N� aJL��gF��b��o>g�gg"��L�h�֒�%����o�i�&<��9|��Ϣ�]���0�8ʬeⷳ$������p�/���1 z(2��+�a溭n!<�5�������%fp;=6V6�D�x���ܹ���.�"�UY�0�9T�bC���Ð ���PSV�M+6�C�����U"ꨨ�G"#bK����?/b��a�j��K	��C���Рq(<$��sl_�^���ƌ�;�U�'f��-�S�t̛7O���>L�b��0����rfB�94~[۷bm�Z,�Z�n_7�D �ԃ�!z�R�����Xd���L��}gO"�}��>�c�R�I�W{,[�L~��bO��ߝ;wb׮]%�rf&"�;�ueuBtڏ���;�{3�������v4�[G�B.�C�*0�6����q�ݻW<)6�2`$�����Du��3��`,<�߼�X�A������g X��� {�6�#xy\�R�6���IT��mVLf��I�`,h	�������R))��a��!��F�>:���Ư{-���uk�e5���m�iarAB����r���<�~�h����&T<�^L�*Y��w6�z]<
_C�,{~0����Dg�S��>�]�pGBGND���=��@����#抦+Ļa���o7"�Ȝ�����h�9P�^M6&�ug'w���N�������-�>�.2�rX�m,2�*op7`�W�A5.]��˰�gϩ�TH x"���@ޜǜ��Z9âAS�*�}֓w@jN�*�tm��L�afn��������!f��?e�(����h<#���9�4s��+�H�ϐ!��C����x�`l�����	����L����g�!�\R���Ig�8��y΂N�+��M[]��B/�p��ڊ�����6�s�=������|��1���G��f��b�N��#���;wZEBlZjZ��(vD���с�a�@veY�2ll�(㐅��b�;�0��i�x�8ĻԶ�WO���*O"-kZ��6���\��Z�@RQg��u��	Cd��hjIXp��p!�[����f����`����3��C��,�c���D��0K`� ��MN�ӅK�"֚)�����NHp������_�fM�f�)�9=�u���XGi?�� +"�7�t��ȒADZ�S�}�7��o�4.?s�aWT�(��?���ق9x��XV�~��er������)��DB�B��õk�ʴ.K͉��u��ˬ��CNX*l^T9�$z�JN�a�p���S]]��(�!֒������p|�9�Ygsn�#�T�1�a줃Y��9[w܎��v�,�gY
jjj���(L���uR����O�����(�/�Bm�[�H[�3~~jJQ��k[����#5y��
�d>]�GWUU�1�L�ϛ�k��Μ�T�-K�T"��uM�pB�Ф{Lt�ۡ'��Y���hmm�ē�rY�X���.�gƪ�;�;�t[WY����Kj�8'<p��믿�����^��h4����YԴ���?� �R�P���s��(��wvj�	ӑ�6g/������԰*[�`�̭�'�N��5 &d�3�~|�RE�z�8׃��4*�k��Zθ�:��A_{?���%#��y�p�9�t8eĞL'U�'��X:x�'�8�w���H�R8-Pp���Z�p��b�M�J��^/L�Vf���"����'��P�j֭�;h�r��N�ө�/r�礄���9�� R�3����+�wC���ց������؍�7�x���,G�B�i�HR�$��A93q������l-\4fd��:^�x���Dw_7~�����M��G� ��b@�H{�s���%R�ϕܯ�:Cv8uHd��6��k���j�*(�nչШ�����<r�#b@9��#���,��TA���»6�qo�^��z����X�-�[���H����.}���bD��"!��Hޱ,E��s�I�K�R��O6�;�d���i���u�oP"7����r�L�����|�|!cD��w��f���5�U_2�}�1����G�rT�����C烺bpU�*D�D��=����6����Z�x5�*���g��[֣�V~J���TX+িH*b�a��k�5]�����b�W�^H��o��-����?�_<���h�"49��q����4�{ٽXQ����i(�,W���<<F�Kz��<�%'|�po������� >������ JK�Kp�^�VX����tUK��dCq1a"p��N!��n\8�BNF���T�j�"R~��'�2�����U�i�|�����<�s�rO]7��9 �3��]����W�%���G^�;cߚ+�%��K��b�yr���~�_�Jl+���a���*yy�Ǯ��u���tY3�����W�BK�emQ,����?������/�><2��e�Y_��ax��>Z�L���X����zdÁ���.�x�+�U�?b�v�`��y�fܵ�.ɗҁ����?~����6�͞f�}�m�84Œ�3�8��u�2A]{��
�>��o��
&V���$1�d �d�(S&o��j5Ye�ˣ�+�D"�8&���~\U�l<0�ph���sj�\	���l�d��pV�]-�B��;���ϣ��(�����P�W��xu�[�o���W%?�cU=���i(�D�tV�s��1Z=�2�Y���ό���ے�󹔜O�r��b8{�Q��������/���0GGFq��<nϴ��^�Ep˂[D��e������薱��,&����Z=/��\���0#&��d͹�)�+��}4^�ۡ:$$#s���S[W{�tV����sެI1�''��h����9� 
�<L���x�^�=n t��$��:C �:��*���cccbG�˺�(C���;�~o�	����e"���eG�˨��*�P��L-����o�k�����$� ���H�Ux�&�͜-ȹP|��esΑ��d���ק�=�;����"!����Aڢ(���*�K�`U�j�����x��^B������!��Hޯ����!�I#K�n�)={O�'*.�g�C�E���{�K�o�'��oO��x.[��7��M�j(�*fo�ĉk%���\[�+����zo��6sc�*��,�ņp[XR��=�N�S�b�z��|�����w���I6���j,�\ ��m���]�n�t`�{#��Ll�!�SbXd9��$�����K/���.�Hz4�N&c�r�G;�ʸr6���
K���_Jrf����K���>�h#6Ԯ,П~�~�O~	�ӻC$���⭡�^IXдi��ɀ�"	��9Yz�^�rO��t-74�f��	�b����WV���α�׿�W��`Z�f]w����6���ͺ�l�";�0��ڄ9zV�+�-��ό�t�[o�����a��h(���t9��#
��"�ب�wE�aZj�u���ɺ��=N�5���j5u��4�z˻�C�s�}��v��Ų��Y\K����/�Iy��'I]}O���<��z���}7|?��?�QB�zŤ�Q����]xz�ӳ
��HL|���\r�H�T2#$%��[�װ(oܸ���B@q7'���4^��F���֪�}��f��7�w����.�t<dP��Jb����-w]�nA7ｨ�FD?n�1�F{A�f)$,�U�*xN$	�����`j8�f��<�ؼ �y �Oe����n��이��L��S��0�����%K�H*%�f��J��ҥKe�H�'��80Umlߵ�=�%Ǟ�sv��ŋe�Fuu��É�ŬVr����r�U�wl�HG��	�ۻ���y�������3��[�T��2�l�� 1���÷͍\:���x�����)�Q�l���Ɲ����{>�0^3�q&���EOJf�74xN�YGʦ���=���'�.�=9��Ib��c˳�:�߇��~�÷IK�3*L���@:
V����K��C�O=�����'����Zn4�������Dy��c�s��l�}~��L XJFͳ���S�,�ng��b�0�a�>�TUWU�*J�ܭ�[Q���϶���Y��E_Cw���bX]�M�cB'��s��� ~ֳ��s���}&*��:�\���j�Z�y�oO�+6��e��y,�l�::�EԈ1������R���l*��țb&�/�f�y�����%�����6�U��R�4f3���[3�&��6ILVF�Zs}�eq��F�G�F�#��t\ֈiYʹ�/��-�VQ�:	�A�o�!b��!��W���~�wdW���ށ��L1���G�xQ��&)r���/�~Q�\��<'�D�t�u���:����uAk����Be�Z����_'�r�K���x�՗�!�����B�1�y��;v�J����3��y��+����}�髷������W��?F�w��]A�y��f����󹛖�/?���8>�i}���x�!���K���Z�8�;��솽���
^d+U8O9mq�"�󖓷/�!���r8�	�\�M~�;o�5�k�;�;�#w/KPt��:�����r.�+΄O��Ϸ��<�R�223x�A�~\q�B >n��Fa@}}=�7�:c�����o>���#��$��ƫ�'�~q������\�kw�1{��4J]���{����mYӂ�5=	���ţgeϖN�U 52��    IEND�B`�PK
     )u�[�W&��*  �*  /   images/b3e67e62-159a-497d-aba3-70fd70f56319.png�PNG

   IHDR   N   �   5�   gAMA  ���a   	pHYs  �  ��o�d  *#IDATx��}ip\ו��{7�Fc%v$����"�Z(J�,��%+��X�ؕrMy*I�&5����W*���5�Ԥj∶5�����D�Z(��. �  ������{.�`/�~�z%�SuQ�~���{�{�yZ��@L�!�(�ώỵ2�V���<Ո?]nE:��{Ct�4����ɴ����6��b(J�����Fa��#6ء4HZt�el�ȓ� qt����U�DXCM����3�&��'�Δ�`����DM�X��z	?���%�Kd�b��,�h@�����ޛ���H�~��"X�<��ƲM��8��Y\�˖�d���KZ�w��O�o��,m�V�F�/c�1����,_:u���8�2�J����M�^J�4�N++���3j��i��P��g{}~x|�_�`$aș�6.�V��V��������^�Q1qz2t������Ob`{jK�j0��aP�1=#�g`W�b����l���SD�A��"-=�_��������Pf�ä'-��O��ݓf��"
����˦���5�L�8�>��T��''N���U�>F-qI\�h|0 ���qk�6@5{�*;E��9��]D��ES0�T���T���r���[�u��O�V���/�9��j�d翂����1AZBJ���OĲ*"�͘�3*6I��b���9�rɣ�P�tj����Zt�._b��2���`V�,W��рnii�$��<ş�ȣ��:����ơb����Ec���b?�Ť��]GJV�p��o/Y<����.��3�+]�
� ]HVXIR��!���o.7��cL	E���%1Ar(���o2B*N��F3˖�������$� Y��>xf��D��A����B�Nh��B���k�����<���g��D��2Ub�8�H�8ZY�&��u�ˁ�PL�&37����re<PL�Zk�7��\�l�	��b�t9��iJ���=ޕ�o("��(M�o*�2��!K6qdTz�[�֑<
��!����:��,�8��~S�H �'1%ĭ +�)�
q
����{`t�B�A���_��W�	�>~�#3T�e���@�|'jT��(+AMY�l���a�����6F���֯�O�ǣ�e%.�1�Zg+�h+5�V+<�ˍ��8w�7U���
��X6∴m�V�ǟEi�tb0�q��n�V����x_;��0`9�,�i�Nlp��?��gc�������Oc��/q߰�˅e!�2ߏڀ�2�r���!�T*AR׬Y��vV���t�Vc��v���j��G]����|>?N��c<u�Bv������:n��z|���5����r �gչ�a��B���YKK+��Б����i���ذ�6���|[2`���aX�dCډ3�fQWj��j��k|�Y����.xl�%����q:�<<^a�^Q^�ڛ_a�i�u��a�7[`�A�`7��8�.�$�o����gv���}�����E�ǖ����:��Bډ�1���D?_����bA�~#_��i'N��@��!Q�u,���v��v��Z&qI N��.$�	�w��6U���[���Z2�jܹ	�u��A�~#[�Xq`"H;qY?��§���Ƈ׻p�]�ˏ����c���"ژp��}�$.@���ѱ1\�̓7ka1��\���
�c�ej}X.��V�E�jN�;�8�X<�����ܵ�����NI��+��6m܀��ȸsM �j։�&:&���qP���h$�9t� �l��������dU��G��d�yM�XP���ju�f�U�i#���n�84��d��Pn6Ð����!�)'������F�9������ǹ[��e�Z�BC�Ʉ�%%��kqϕ����,3�VVbr~���wz�+u1LLL�w�� 2�^�}p?z�9X,�S�l�c��ɐ�-k*��1���S��w'�Bʈ+g�bw���/JM�ũYFq}��݋��}0mm��8��Ӌm[��e.	�f�9��tH^J���(����%N�,�I�^�csy�{�C�j�K�'�ɺzN���$n�� UH:q�A��&?�Ȝ�S�ԬǕ;���3Gه���?+z<���p�L�>"�TJ^R�J�I����:��HVV~��g���U��uG�Aw_,��愉�[S���><���T�h�����0���SJؼI��i�V�u�B%/H
q4H���K�8���|iw$�4�oJ�΂+�'u�&U���I�N���P����T�?	OOy��ǐ�%�LzãE\�,�6�^:*0<)�χ���E��8o4�g�j����OS��nF��4����E^��Ք�Ĕ� ���0--m8wo-��|�J;�z�� h���͈�>��GnJ2E�đ��`1OpI�p��vx4zhsK�w;�37-� ��MUJS�IZ2EB�Q�N�C��8�h����[K;��\�	��t����9�-\��Kd((� ?3Q$D\h�#�d���т�4�[�a)�bG��Ousn��D��uى��F�ፄu~Zr��P]]�_r@δ}~�3| iKV��8R�d�F��d5)"H�8��� �doM'�AQ�?�_B���OrCc�S�Z{Pɨ��}�e@���\W�>7�&v����g���L���َ��͒�g��1;7�̜bY�HV�N1qd��1�c�X��)yLgg�|�*޻3���g���Xx��̲��&eG�Ur��<x�D��8�B�:Nc�����1���ۿ�?o��#���Y2Mx`�A<��jU��du�̪q�R�JgFrss���]�Y�֚g���{��Jx��%�� ���đu���8���[���ƍ�x~|���>^�&f���ū*���U�Ѵp�lS5^���P���C�öm��mQ�l�}|�9�Y�5$4�e5�G�]:����R+����h�/?��!ũ����>�B��o#*dR��Y!�%/�����%/[�U�J�����.?v�ՠ�@��1�h�i��S�B.Z�M	�#D�rr\���a6U�$�g����!�骸q�q����/I֒PF��,p4Mi�7�̄b r&�f��¤�I�Xzzzq�]�iS�;7�EOo/��l�I���0r�923��uH�绗�8(X��k"���>F�_��5Z��7�A3kw���``7�b�⋳���g^�$w�,$Dݹ`2S$iD��hv�EKX���Y����aq�1��<'���K~ga�ֿt�=��	�Gӳ<���I��B�h������_2�I0ge�g��@ww7�j���J.`HǙ�RI7�$o��ǰv]�>.�$	Gw�^��?T�BA���XU�ɈM����3�J�(��o:?ݰ�λKҗ�:��-Hi�R� TI�	�N+�S�n����7�?����0��_I�,�9�̎�~��vԸ��r@�Z��^�ϤT����ᨆzt#V��a�$�'TR��l�"؏�j��svr|���z���1j�07Ώ��m8�Ò�!�KӥL�������E�D�=�?I�jm��K�8��'D���Y��4�Q_Kk�=E@͓������z�gM�����jaL�l0m��@���M���T2��%D�i�u;PX��**q���fc�(��]f������ �-����؝6�k�W���w��5u����k�(GM�"ISg����t!��j�����Te�l:�\�6Â9g ��P����31���2ŕ��*�)Z^1\�M)!Oq$���ֈ,����+��WH<H%��ء��:~��b�01�e��=(*Z�{:^Һ��
�L3j�J0i����'D�6#'���qGj�H�DEnxF�J�3�j}�:��dY��$�5�36tCuL�<��a�9�Za�ܮX��M�0d֔����E%���䮩�"ˤ%Q�z�$.��o�E���v�?���(��Q<e��xw�^#�I���R�L	��RG���h�$���<,��% Oy4e�z��F�q]�w&B�1��n�+F���[$�x��۰�x`�L���LM�1�ٔ���vM)%��-ұ$�F.Y1��\�kVKU'�5k*�4����f����I4��躹�� %�3�M\d�a�6R�\��/�x&:����T"�>44�{����0'���~TTT`�����
�|Q�*��&���3�Q�y𦒥�;�ʎu#^�$.z�^#�9i��,L�wv����������믑�����Z�ݻW𸾾>~���<<�u뢭���?aN�К�]J+ј�ٔ��"%��=A��4�/t�L������R����5��!��
�X�l7q��}����{�=ޡ�ĉ1sn�W��/�Ӊ����K����Î��\���8�ٻp���R�3ª��㵻��#LŤ<���g���X�"����BgZܣ�QA3|�qt��m�eE�X���Ř��n�P��v���رc���H�h4�ȑ#��>�z�-����a�!� �gE�<�m�n��������v2C����s~9̲��ͱ��[mĀ#v_qCC�h��%��U��v�3�T����=o�H;t�V�����uff&�~�m��F���i1{����w�P�:Q|u����wаg�h	Fq�ͷ��t�w��{��?��صkWB�Q^^�.Ԇ>��O�d 33��V�����6^����0#�D�͛M������EM�d��ݻ0��LU
~NS�����&P;[*{-..f���xE�$o`` ���l�V'u�%l�=w�(>��K4^������q⺺�����s�=�)5�󯱓���+��ݸq�_|}}=�m�����0�*rG�l�^_%+{�ԩ�G�ť��:���AA~���3N\��k\SEZgg'���.J[ʟ~�i���{��t��;�<�b�����Af�c������];p��z8q�K�B���W�;w�`���Q�ONN2i�������3g��U�'�|r�����ܹs�G���7rU�
���jm��Km�u������ᶰ���qR��q
�Qho��J�t�X�lzz�;���r�
wK"A����H�T�z�j�$�� ��2���=,
Q��;::y�NJ�F�V�褏q�D���vn�u���'�}�G�I౵���+/��|t�ڧا�Bh����C��������,�frA����ۂ�Dk<Ǣ�w?8�9S%O��=��O#�O�>��~̸UX���O<��5a�Cd��>���Z�6&��%����5�V[��i�h�X��6Ƭ_��,�7-�Q^�j4߻E9��F�͜�Л@A4�)F}�� A�&��AK���1�Y�B87�{��z��,$^�����g�6�7�F���Qđ�h�?\�ЪD���R띇���{�{A�}~�!n�Z��.)�Mz�JMMM-}��xx��M]�uY�;<i��#8�]0����}n���Ha����^Oy_k`"K����k+Q��5�jL�;���ȳAP�Ԫ-��>ì���ͨ�=M�R��E����K�s�:��1ק���_�_�K��v'��M��aZ]>������sK�S[������Ű͇�-��G�`PTa�%����/��UB����̕ �P�B�����;��w�a�ڍҺZ�qG�.F�b�T��*��&	�7�[��?y�)^�IRS���E������QԮo�-��Y1M	�2<,��R���@�+ ��^bа��uk�%��bѿ�hhh�~܁ ���a.JD�T&��R�ed(ĺ���7�\�ʥ��6T�7�����MqU{���)��z��E��� (	YPx��-�D`����}?� B�ر��c�F�	�w����M,�����uuu���-�=��8�<���I��4T2)�mjj�Ⱦ}��	�9~�Y�8��t�k7����>7�۷o�Y�^\�҈�{R2 �� ��ȣ`��[rS��������������&T���(az�&�\wɟ8r�0>9s_^��=�]!�+���<y�Y�5�QM����ɨeDBA	 z�Ź����ï^]��):��D��g�l���#��;�Y�X���^x������_�
�H#"Z����k�%m|�[���&��.&@��κDe���i�CoƯ���a��K��k�m�Di^�	�x���~��6eT�m�`cUE�Z�W�����?s)�'�
���(.\��o�PF�
���o����BA�sz��.�P��[��<ӧ�� �|����dŻ��CV�����,�c��������B��ݍ���و -�L��VW3�Ww����<~��/��"ϱQm�֭������ū����Q���W_�J�μMP���K�0�u~�,���Ew��Kn	��	�\��B�J���/an#.?����Z��a)��l+��|	��/q�h��E:��7��ŋ��?��+^2b"(�hmm�y�M�6E�3q�/pӾƺ}���^�2�SqÃţ������E���&8*^�"���|��Qx�{wD?f�_z���裏�ĐA&
Ղ� �4D�n�hB�#Ƶ�D��{�|5�ʾ��Mdg,ݸ���E�m��US%���Q�-�O	�(A7��r-YU2z�[�o��m�k�*�.�����$E^��&N#P:@��MY9\�j�J��,}�\��>���ٸK�6֞�H�W��dAmގt��4;� ��c��.%�qU+EI#qn��W�K�d�)'�8%�L�]%��Pa�g�wx����)A\�ѝ�|lp��l�I�B!_֢�{5S�4S'�m�:#����јn�Ȍ����K_E&=K�XVc��k���@5(�"έ��R�*�]n8�9") ��q�B
	|FԊ�$�v��^�LӀ����;�y.��Š�$�V�i5���`ˆu�i� �.'Tڇ7�,gA��K��+��@�eV�G"PD��v�P]Yym��ʼq��榨tF��b?jll��SE�Snw�������ƴ���U`R��mz4�4�R�
Ņ��먫`d��t�u�V�CF�B���ủ�����Ma�d�^J�L��,J�IeT<�m�\TyI�Ý���'!c͎���H��9�#"ɣw�{��t���d*�62�Բ���m�c��t��<8�����S`���d��ǚ�ɣ��H�A�ʴ�`�X�qo�-��5�hj���V5>d��X8v$��Fgf1�q��[���H����z"�v����A��S�h�	��b7N�H�������j9�]�[V���w�?��]�NO:-��d��`k_(z���q���%x�󘞑ײ��^n��A<��,Υ	pјH����mا7�łl��A��N&4�����B|=� 
e�9�9½8rn��4���r�h���m��N23��Y��|z�8�����A>��c�2**5���9z�� ��X��ڑ�ulj�&����󋔪0�ϩew��4W��K��K�K6$u2�j���X�\rt�Ϛi����ܻf(`���)E���u-�gv�=��������@dk�r�����D��8�=q��EJ���^�Cb�8cĸ������>_>-Q��\�.�H)PU����U���c�*�+��,�t3�����ŹcH�����1ܸ�Rk���aU�t��b��N����r �8��Kl���CWg�d�U�������,���	6n����9G��$�IÐ�4b�0�)�4�1k��� ��o�,���6U�	�e�`djnis^:�6����"c����8��ud8�g;�m��[�z=���i�8�H)�wt���a��kh��bz�W����F����8��Z54�}��������e�vI�#�c�0ݼ��w��]�/`��I�f�m�SUŢ��z/�8�4F7����T(&ΤW#Sz�U00"��9�7jO5]���t�ټ�<��/�ی �GV�܉|���P���H��}ߤװJ�
zv�:M��i~�r�g����v�A��ц�ϧ�t���I'N�ْ�K�v9���E3V��T5����� z����U���8�>F�O&uvO ������E����B����O+O)iè#�a�L��wz��)"N��wL�v���Hde�.,����y����isa'�&x*��v�yk�f������YT����9N���2��ĸc^_�t�A��1sr��6sxfgQ�{�䂴��]�B��I�"�s����|0H4�r��
�� �
�?x�Н�4�Z�>���/��'��$�S	<������%A��H���͚cV3��$����8�[X��4Zx��BD����A��Y�M-t���ӌ��~Q�ȡ�wo��q��0i��H�����I̗S�ǹ�ɧ؋`R�T�L���0S�N�=OSPH�0��K�Zq��"�ZbG���@7��:&y��\�x��(I$r9�E@-���T���O`*'z��*��A4���cW��F���G
�H_"�a�!-q䷽��7y	U�Ӧ3��o/E��ǩ���gJ'V�j~I�䀦ꔕ�Uj�WHAq��W��s�6+�kk��#d��B�*�_ʺy�.D����"�^X����ȐFQg
��i74��<T�{���A	�2!^�&��]����i�%2���$����߹'^}Y|��ǻ��1�x H\y~6L����J-IeH���_|����|��ڶ�a�Ȃ49������cAT�^ڷ�_nM*y|�AªRI�!�X�Ԕd����U0�(~y<��]Q���}yOm)��O���s�p[�y҂��M�a`��}b�;{�b��=��.�����
�h�)KL�5���,�������
�����O�r�h���$��38��lٗ�]�RH��r��e���Ժ�R�45����r ��Qc ��ˉ���q����n��8s����Y����a�U��f$�������v6�
���u���s�33���ޡB������H�]�����O�sEu�
�z����y��S�M�S�����"A�2M����b��'ǲ�EZ�sv7CǤ�W!�u���6d-�rS7�P���*�[�����з�8%�J!��oGFy9�ns�+ܹ�7>�MI�k�KXǭ&Tm݉t"��9zn���`jjZpVmm5&_<��ټ&o�3O�F���bQÂ��h���4Gڈ��u8{o���,�u|���غmώHu�5�.>�m9�\���fG��~��ws����;�455�X�t빴G�����Ô�xƖ�.9g��.��'�Uϥ���/�����V��̊784�k�ݳsؼ{�E~A�V�!+\����B� *�`����(�|�wП����i}�Y�����ѥ^n�<�!��ҭ��B���'K��R��<����O�"wz��L�-� -D���\�D#���y�i!.8M	f�����т�6dAڣш>x��jOx����	�~K��92���sC<�}����{O<�)���/g�Z�ދ޻J=��LW�#�r6~r����i��)'�;;��*��w��x;���R������{A���=�Ђ���70�|:ot>]nIJ�#�0�L���:'�._@u�֨N�T�TS#��r��ݽ�S����kU|-�!�ą�P��p�p�ˋ8���Z;f��B��̈��P���s��s)%.r��b�����Y�S��`O�N�Z[
�����khس��,�����ݏH�[���8�iD�o�:�������.^Bqa,f3,e�<�I�JF��e�Ӳj���1����E	�#�;�\ʈuz#A�q����u���ŕ��p��P/�m�MM��v��_�5��>�r�ĉI�?�2���!k�Ѩ��2�?��b5<�Y�@߹�۶���~:���'�ߌk7{R}:�֔'��h��$��6鱩o�b��~K&r�JE-+E2�zJ�4⺻���768ğwcԩ���P�� ����m�Z3K��{��=�o����3���
�bzɻ�s�j~�xJ�:766�ܝ�>0)��#?�}�S�.����"��3���t�Q�[��1#�<����GF�?39�I�.�4ó��ۿE�y��!-^��ǯ3w�{H&����x�ߣ�+�ɝHݚc���p�4bXD����z����~��_^Q!�>%H�8zt��ӑ%�ԕ�$�)N���+�)�
q
�B�B��+�)�
q
�B�B��I'�J������~_x�O�t�bu�I'���$��T�{���b�8�X!N!V�S��b�8�X!N!V�S��")ĥ2�I�=Ƅ����x�G/7����8���؏䓃�HeC��x�G+:N!�N��l��>�����\�������x��h�E꩜��F����{N*�T������9qb$<x���#��D"M��O���!�0���b7�ʼe?�:^$�8���/R(L����Dm�USY�bϥH���������j
"����_#���TGG�� ��cY^"���B��yT��"��B�?	D%��`�7,L��qY"3�r�5��="3��+VU!V�S��maS'��I�>SSS���|Rp��h�j������zoo/��"!�G5���ޗj*O�uuu	.I��S�S�#8���`�u���4$mtL$y$iDId����BM�Ȋ�w�C5߂G��EZ,���C�w�<4=����w�8$�=I�8
��[�֔�D@ӝB:��� a�jjj��;�|�$�,�dy�0<4�7~�&�Z�,$e����}���q������g���    IEND�B`�PK
     )u�[�W&��*  �*  /   images/ab942d8a-eab6-45a7-8f5a-30ef729b6f10.png�PNG

   IHDR   N   �   5�   gAMA  ���a   	pHYs  �  ��o�d  *#IDATx��}ip\ו��{7�Fc%v$����"�Z(J�,��%+��X�ؕrMy*I�&5����W*���5�Ԥj∶5�����D�Z(��. �  ������{.�`/�~�z%�SuQ�~���{�{�yZ��@L�!�(�ώỵ2�V���<Ո?]nE:��{Ct�4����ɴ����6��b(J�����Fa��#6ء4HZt�el�ȓ� qt����U�DXCM����3�&��'�Δ�`����DM�X��z	?���%�Kd�b��,�h@�����ޛ���H�~��"X�<��ƲM��8��Y\�˖�d���KZ�w��O�o��,m�V�F�/c�1����,_:u���8�2�J����M�^J�4�N++���3j��i��P��g{}~x|�_�`$aș�6.�V��V��������^�Q1qz2t������Ob`{jK�j0��aP�1=#�g`W�b����l���SD�A��"-=�_��������Pf�ä'-��O��ݓf��"
����˦���5�L�8�>��T��''N���U�>F-qI\�h|0 ���qk�6@5{�*;E��9��]D��ES0�T���T���r���[�u��O�V���/�9��j�d翂����1AZBJ���OĲ*"�͘�3*6I��b���9�rɣ�P�tj����Zt�._b��2���`V�,W��рnii�$��<ş�ȣ��:����ơb����Ec���b?�Ť��]GJV�p��o/Y<����.��3�+]�
� ]HVXIR��!���o.7��cL	E���%1Ar(���o2B*N��F3˖�������$� Y��>xf��D��A����B�Nh��B���k�����<���g��D��2Ub�8�H�8ZY�&��u�ˁ�PL�&37����re<PL�Zk�7��\�l�	��b�t9��iJ���=ޕ�o("��(M�o*�2��!K6qdTz�[�֑<
��!����:��,�8��~S�H �'1%ĭ +�)�
q
����{`t�B�A���_��W�	�>~�#3T�e���@�|'jT��(+AMY�l���a�����6F���֯�O�ǣ�e%.�1�Zg+�h+5�V+<�ˍ��8w�7U���
��X6∴m�V�ǟEi�tb0�q��n�V����x_;��0`9�,�i�Nlp��?��gc�������Oc��/q߰�˅e!�2ߏڀ�2�r���!�T*AR׬Y��vV���t�Vc��v���j��G]����|>?N��c<u�Bv������:n��z|���5����r �gչ�a��B���YKK+��Б����i���ذ�6���|[2`���aX�dCډ3�fQWj��j��k|�Y����.xl�%����q:�<<^a�^Q^�ڛ_a�i�u��a�7[`�A�`7��8�.�$�o����gv���}�����E�ǖ����:��Bډ�1���D?_����bA�~#_��i'N��@��!Q�u,���v��v��Z&qI N��.$�	�w��6U���[���Z2�jܹ	�u��A�~#[�Xq`"H;qY?��§���Ƈ׻p�]�ˏ����c���"ژp��}�$.@���ѱ1\�̓7ka1��\���
�c�ej}X.��V�E�jN�;�8�X<�����ܵ�����NI��+��6m܀��ȸsM �j։�&:&���qP���h$�9t� �l��������dU��G��d�yM�XP���ju�f�U�i#���n�84��d��Pn6Ð����!�)'������F�9������ǹ[��e�Z�BC�Ʉ�%%��kqϕ����,3�VVbr~���wz�+u1LLL�w�� 2�^�}p?z�9X,�S�l�c��ɐ�-k*��1���S��w'�Bʈ+g�bw���/JM�ũYFq}��݋��}0mm��8��Ӌm[��e.	�f�9��tH^J���(����%N�,�I�^�csy�{�C�j�K�'�ɺzN���$n�� UH:q�A��&?�Ȝ�S�ԬǕ;���3Gه���?+z<���p�L�>"�TJ^R�J�I����:��HVV~��g���U��uG�Aw_,��愉�[S���><���T�h�����0���SJؼI��i�V�u�B%/H
q4H���K�8���|iw$�4�oJ�΂+�'u�&U���I�N���P����T�?	OOy��ǐ�%�LzãE\�,�6�^:*0<)�χ���E��8o4�g�j����OS��nF��4����E^��Ք�Ĕ� ���0--m8wo-��|�J;�z�� h���͈�>��GnJ2E�đ��`1OpI�p��vx4zhsK�w;�37-� ��MUJS�IZ2EB�Q�N�C��8�h����[K;��\�	��t����9�-\��Kd((� ?3Q$D\h�#�d���т�4�[�a)�bG��Ousn��D��uى��F�ፄu~Zr��P]]�_r@δ}~�3| iKV��8R�d�F��d5)"H�8��� �doM'�AQ�?�_B���OrCc�S�Z{Pɨ��}�e@���\W�>7�&v����g���L���َ��͒�g��1;7�̜bY�HV�N1qd��1�c�X��)yLgg�|�*޻3���g���Xx��̲��&eG�Ur��<x�D��8�B�:Nc�����1���ۿ�?o��#���Y2Mx`�A<��jU��du�̪q�R�JgFrss���]�Y�֚g���{��Jx��%�� ���đu���8���[���ƍ�x~|���>^�&f���ū*���U�Ѵp�lS5^���P���C�öm��mQ�l�}|�9�Y�5$4�e5�G�]:����R+����h�/?��!ũ����>�B��o#*dR��Y!�%/�����%/[�U�J�����.?v�ՠ�@��1�h�i��S�B.Z�M	�#D�rr\���a6U�$�g����!�骸q�q����/I֒PF��,p4Mi�7�̄b r&�f��¤�I�Xzzzq�]�iS�;7�EOo/��l�I���0r�923��uH�绗�8(X��k"���>F�_��5Z��7�A3kw���``7�b�⋳���g^�$w�,$Dݹ`2S$iD��hv�EKX���Y����aq�1��<'���K~ga�ֿt�=��	�Gӳ<���I��B�h������_2�I0ge�g��@ww7�j���J.`HǙ�RI7�$o��ǰv]�>.�$	Gw�^��?T�BA���XU�ɈM����3�J�(��o:?ݰ�λKҗ�:��-Hi�R� TI�	�N+�S�n����7�?����0��_I�,�9�̎�~��vԸ��r@�Z��^�ϤT����ᨆzt#V��a�$�'TR��l�"؏�j��svr|���z���1j�07Ώ��m8�Ò�!�KӥL�������E�D�=�?I�jm��K�8��'D���Y��4�Q_Kk�=E@͓������z�gM�����jaL�l0m��@���M���T2��%D�i�u;PX��**q���fc�(��]f������ �-����؝6�k�W���w��5u����k�(GM�"ISg����t!��j�����Te�l:�\�6Â9g ��P����31���2ŕ��*�)Z^1\�M)!Oq$���ֈ,����+��WH<H%��ء��:~��b�01�e��=(*Z�{:^Һ��
�L3j�J0i����'D�6#'���qGj�H�DEnxF�J�3�j}�:��dY��$�5�36tCuL�<��a�9�Za�ܮX��M�0d֔����E%���䮩�"ˤ%Q�z�$.��o�E���v�?���(��Q<e��xw�^#�I���R�L	��RG���h�$���<,��% Oy4e�z��F�q]�w&B�1��n�+F���[$�x��۰�x`�L���LM�1�ٔ���vM)%��-ұ$�F.Y1��\�kVKU'�5k*�4����f����I4��躹�� %�3�M\d�a�6R�\��/�x&:����T"�>44�{����0'���~TTT`�����
�|Q�*��&���3�Q�y𦒥�;�ʎu#^�$.z�^#�9i��,L�wv����������믑�����Z�ݻW𸾾>~���<<�u뢭���?aN�К�]J+ј�ٔ��"%��=A��4�/t�L������R����5��!��
�X�l7q��}����{�=ޡ�ĉ1sn�W��/�Ӊ����K����Î��\���8�ٻp���R�3ª��㵻��#LŤ<���g���X�"����BgZܣ�QA3|�qt��m�eE�X���Ř��n�P��v���رc���H�h4�ȑ#��>�z�-����a�!� �gE�<�m�n��������v2C����s~9̲��ͱ��[mĀ#v_qCC�h��%��U��v�3�T����=o�H;t�V�����uff&�~�m��F���i1{����w�P�:Q|u����wаg�h	Fq�ͷ��t�w��{��?��صkWB�Q^^�.Ԇ>��O�d 33��V�����6^����0#�D�͛M������EM�d��ݻ0��LU
~NS�����&P;[*{-..f���xE�$o`` ���l�V'u�%l�=w�(>��K4^������q⺺�����s�=�)5�󯱓���+��ݸq�_|}}=�m�����0�*rG�l�^_%+{�ԩ�G�ť��:���AA~���3N\��k\SEZgg'���.J[ʟ~�i���{��t��;�<�b�����Af�c������];p��z8q�K�B���W�;w�`���Q�ONN2i�������3g��U�'�|r�����ܹs�G���7rU�
���jm��Km�u������ᶰ���qR��q
�Qho��J�t�X�lzz�;���r�
wK"A����H�T�z�j�$�� ��2���=,
Q��;::y�NJ�F�V�褏q�D���vn�u���'�}�G�I౵���+/��|t�ڧا�Bh����C��������,�frA����ۂ�Dk<Ǣ�w?8�9S%O��=��O#�O�>��~̸UX���O<��5a�Cd��>���Z�6&��%����5�V[��i�h�X��6Ƭ_��,�7-�Q^�j4߻E9��F�͜�Л@A4�)F}�� A�&��AK���1�Y�B87�{��z��,$^�����g�6�7�F���Qđ�h�?\�ЪD���R띇���{�{A�}~�!n�Z��.)�Mz�JMMM-}��xx��M]�uY�;<i��#8�]0����}n���Ha����^Oy_k`"K����k+Q��5�jL�;���ȳAP�Ԫ-��>ì���ͨ�=M�R��E����K�s�:��1ק���_�_�K��v'��M��aZ]>������sK�S[������Ű͇�-��G�`PTa�%����/��UB����̕ �P�B�����;��w�a�ڍҺZ�qG�.F�b�T��*��&	�7�[��?y�)^�IRS���E������QԮo�-��Y1M	�2<,��R���@�+ ��^bа��uk�%��bѿ�hhh�~܁ ���a.JD�T&��R�ed(ĺ���7�\�ʥ��6T�7�����MqU{���)��z��E��� (	YPx��-�D`����}?� B�ر��c�F�	�w����M,�����uuu���-�=��8�<���I��4T2)�mjj�Ⱦ}��	�9~�Y�8��t�k7����>7�۷o�Y�^\�҈�{R2 �� ��ȣ`��[rS��������������&T���(az�&�\wɟ8r�0>9s_^��=�]!�+���<y�Y�5�QM����ɨeDBA	 z�Ź����ï^]��):��D��g�l���#��;�Y�X���^x������_�
�H#"Z����k�%m|�[���&��.&@��κDe���i�CoƯ���a��K��k�m�Di^�	�x���~��6eT�m�`cUE�Z�W�����?s)�'�
���(.\��o�PF�
���o����BA�sz��.�P��[��<ӧ�� �|����dŻ��CV�����,�c��������B��ݍ���و -�L��VW3�Ww����<~��/��"ϱQm�֭������ū����Q���W_�J�μMP���K�0�u~�,���Ew��Kn	��	�\��B�J���/an#.?����Z��a)��l+��|	��/q�h��E:��7��ŋ��?��+^2b"(�hmm�y�M�6E�3q�/pӾƺ}���^�2�SqÃţ������E���&8*^�"���|��Qx�{wD?f�_z���裏�ĐA&
Ղ� �4D�n�hB�#Ƶ�D��{�|5�ʾ��Mdg,ݸ���E�m��US%���Q�-�O	�(A7��r-YU2z�[�o��m�k�*�.�����$E^��&N#P:@��MY9\�j�J��,}�\��>���ٸK�6֞�H�W��dAmގt��4;� ��c��.%�qU+EI#qn��W�K�d�)'�8%�L�]%��Pa�g�wx����)A\�ѝ�|lp��l�I�B!_֢�{5S�4S'�m�:#����јn�Ȍ����K_E&=K�XVc��k���@5(�"έ��R�*�]n8�9") ��q�B
	|FԊ�$�v��^�LӀ����;�y.��Š�$�V�i5���`ˆu�i� �.'Tڇ7�,gA��K��+��@�eV�G"PD��v�P]Yym��ʼq��榨tF��b?jll��SE�Snw�������ƴ���U`R��mz4�4�R�
Ņ��먫`d��t�u�V�CF�B���ủ�����Ma�d�^J�L��,J�IeT<�m�\TyI�Ý���'!c͎���H��9�#"ɣw�{��t���d*�62�Բ���m�c��t��<8�����S`���d��ǚ�ɣ��H�A�ʴ�`�X�qo�-��5�hj���V5>d��X8v$��Fgf1�q��[���H����z"�v����A��S�h�	��b7N�H�������j9�]�[V���w�?��]�NO:-��d��`k_(z���q���%x�󘞑ײ��^n��A<��,Υ	pјH����mا7�łl��A��N&4�����B|=� 
e�9�9½8rn��4���r�h���m��N23��Y��|z�8�����A>��c�2**5���9z�� ��X��ڑ�ulj�&����󋔪0�ϩew��4W��K��K�K6$u2�j���X�\rt�Ϛi����ܻf(`���)E���u-�gv�=��������@dk�r�����D��8�=q��EJ���^�Cb�8cĸ������>_>-Q��\�.�H)PU����U���c�*�+��,�t3�����ŹcH�����1ܸ�Rk���aU�t��b��N����r �8��Kl���CWg�d�U�������,���	6n����9G��$�IÐ�4b�0�)�4�1k��� ��o�,���6U�	�e�`djnis^:�6����"c����8��ud8�g;�m��[�z=���i�8�H)�wt���a��kh��bz�W����F����8��Z54�}��������e�vI�#�c�0ݼ��w��]�/`��I�f�m�SUŢ��z/�8�4F7����T(&ΤW#Sz�U00"��9�7jO5]���t�ټ�<��/�ی �GV�܉|���P���H��}ߤװJ�
zv�:M��i~�r�g����v�A��ц�ϧ�t���I'N�ْ�K�v9���E3V��T5����� z����U���8�>F�O&uvO ������E����B����O+O)iè#�a�L��wz��)"N��wL�v���Hde�.,����y����isa'�&x*��v�yk�f������YT����9N���2��ĸc^_�t�A��1sr��6sxfgQ�{�䂴��]�B��I�"�s����|0H4�r��
�� �
�?x�Н�4�Z�>���/��'��$�S	<������%A��H���͚cV3��$����8�[X��4Zx��BD����A��Y�M-t���ӌ��~Q�ȡ�wo��q��0i��H�����I̗S�ǹ�ɧ؋`R�T�L���0S�N�=OSPH�0��K�Zq��"�ZbG���@7��:&y��\�x��(I$r9�E@-���T���O`*'z��*��A4���cW��F���G
�H_"�a�!-q䷽��7y	U�Ӧ3��o/E��ǩ���gJ'V�j~I�䀦ꔕ�Uj�WHAq��W��s�6+�kk��#d��B�*�_ʺy�.D����"�^X����ȐFQg
��i74��<T�{���A	�2!^�&��]����i�%2���$����߹'^}Y|��ǻ��1�x H\y~6L����J-IeH���_|����|��ڶ�a�Ȃ49������cAT�^ڷ�_nM*y|�AªRI�!�X�Ԕd����U0�(~y<��]Q���}yOm)��O���s�p[�y҂��M�a`��}b�;{�b��=��.�����
�h�)KL�5���,�������
�����O�r�h���$��38��lٗ�]�RH��r��e���Ժ�R�45����r ��Qc ��ˉ���q����n��8s����Y����a�U��f$�������v6�
���u���s�33���ޡB������H�]�����O�sEu�
�z����y��S�M�S�����"A�2M����b��'ǲ�EZ�sv7CǤ�W!�u���6d-�rS7�P���*�[�����з�8%�J!��oGFy9�ns�+ܹ�7>�MI�k�KXǭ&Tm݉t"��9zn���`jjZpVmm5&_<��ټ&o�3O�F���bQÂ��h���4Gڈ��u8{o���,�u|���غmώHu�5�.>�m9�\���fG��~��ws����;�455�X�t빴G�����Ô�xƖ�.9g��.��'�Uϥ���/�����V��̊784�k�ݳsؼ{�E~A�V�!+\����B� *�`����(�|�wП����i}�Y�����ѥ^n�<�!��ҭ��B���'K��R��<����O�"wz��L�-� -D���\�D#���y�i!.8M	f�����т�6dAڣш>x��jOx����	�~K��92���sC<�}����{O<�)���/g�Z�ދ޻J=��LW�#�r6~r����i��)'�;;��*��w��x;���R������{A���=�Ђ���70�|:ot>]nIJ�#�0�L���:'�._@u�֨N�T�TS#��r��ݽ�S����kU|-�!�ą�P��p�p�ˋ8���Z;f��B��̈��P���s��s)%.r��b�����Y�S��`O�N�Z[
�����khس��,�����ݏH�[���8�iD�o�:�������.^Bqa,f3,e�<�I�JF��e�Ӳj���1����E	�#�;�\ʈuz#A�q����u���ŕ��p��P/�m�MM��v��_�5��>�r�ĉI�?�2���!k�Ѩ��2�?��b5<�Y�@߹�۶���~:���'�ߌk7{R}:�֔'��h��$��6鱩o�b��~K&r�JE-+E2�zJ�4⺻���768ğwcԩ���P�� ����m�Z3K��{��=�o����3���
�bzɻ�s�j~�xJ�:766�ܝ�>0)��#?�}�S�.����"��3���t�Q�[��1#�<����GF�?39�I�.�4ó��ۿE�y��!-^��ǯ3w�{H&����x�ߣ�+�ɝHݚc���p�4bXD����z����~��_^Q!�>%H�8zt��ӑ%�ԕ�$�)N���+�)�
q
�B�B��+�)�
q
�B�B��I'�J������~_x�O�t�bu�I'���$��T�{���b�8�X!N!V�S��b�8�X!N!V�S��")ĥ2�I�=Ƅ����x�G/7����8���؏䓃�HeC��x�G+:N!�N��l��>�����\�������x��h�E꩜��F����{N*�T������9qb$<x���#��D"M��O���!�0���b7�ʼe?�:^$�8���/R(L����Dm�USY�bϥH���������j
"����_#���TGG�� ��cY^"���B��yT��"��B�?	D%��`�7,L��qY"3�r�5��="3��+VU!V�S��maS'��I�>SSS���|Rp��h�j������zoo/��"!�G5���ޗj*O�uuu	.I��S�S�#8���`�u���4$mtL$y$iDId����BM�Ȋ�w�C5߂G��EZ,���C�w�<4=����w�8$�=I�8
��[�֔�D@ӝB:��� a�jjj��;�|�$�,�dy�0<4�7~�&�Z�,$e����}���q������g���    IEND�B`�PK
     )u�[��n GV GV /   images/5a738b76-89aa-4728-b8e5-f09c859dbb14.png�PNG

   IHDR  �  "   �?��   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  ��IDATx���|w���������j�dɲ,˽�v�$!q��;:� �H.wGr$��B�����s)$�@(C��;.�w˖l�����&�Ųg������gƊ�7kiFZ�|������LB                 d�]                 � �                ��@�                ��                rw                @N �                �	�                9��;                 'p                ��                ��@�                ��                rw                @N �                �	�                9��;                 'pϲ�Sgj�vړ�&���{�����4��oxL���E               ��s9l��n�ץ|�C�M���>'����"�Dc�h`$�a��	!�����"�^՗jz�PUE>�#���B��������7���aI.ۺ����_{���w($               `���/�kz�@5e���nE�/���8�?2�=8����ݎޑ��j�$��&�Mf�-5�j�-֜䲱�/��a�~v�����2��֖=�z�[;���               �Dg4�6��sj�S���ӊT�e_����0�����}ښ���h���T'���	2:�7V��tf��55;y�oWv��\Z�\��P$�W�Ն7�j����               �(�|��Ơ�5�k�2x�Y}=F��Y�E�q��7?ftvqg�6�qD��w+�A�� �~��:��Jo[P��"�r��a��Ը�]���~��~��ں�               �#ľ��\�ϩ���rٲ݅�/�,H��:u���"z~{{*�k�	�;��P���;���u�*��DU[V��i�fm;أ�lث�li�X8&                [�������u�P{�g���<�Cg/�I���~��~���T�j�y܏���]��A+�+e��gɟ0{ZQj|��yzr�A���]j뢫;               2'��҅�R����ݚL
}.]rrcjl�߭G^ح��R,��/���c?mN��&���&;�ۡ�'���e�S�!<��.m��%                ]j�
t��3���5rح�����Ƒ�=��.���}G��A��X-��R���E�J�4����+S�xB�_�ܦM{;               ���4_�9�IgͯI5��j�~�>~�<��Yz��z�]��ϊY���-�++�|B�+9U/�qD��|��t�               8^�]vv�޶`j��P�ש�٬w-��������{�'4�pO2:���y:if��-kjɌ2�j�A���f��               +�ݪ�V��{Ϙ%���*�w��w-Ѕ�g�'^�;:4UM���鲷�$��x�ϲZ,:{AM�����E�oث��~8               ��ȟ^w��z�?�h�}��W�����oT�����)p�_W�.\���A�c��v�,�����ˏ����               �����Gϙ�j���Y�\�Ee��u��g�P|
u��rw�Ӯ�ϛ�s�	�oNm������Γ[��s���              ��9}N�>q�x���q;m��s���\�{�%��T0��M��|�RUӵ�N�M;g��7U$O��               �.�æ��>G�h�1��D߾�,}���䦃��D��b�.Y٨��1Gv�E0���R�w�Y�����Ү#              ��3=X��w/Wu	ͨ��s;tӥK���L_{|��&�Ip�8�q�"�1�ZH�B�K������3;��_lU<�               ��U�uㅋ�vڄ�9gq�+���|A�#��&u��<���_���!��N�}�LU�鮇6h,<y�              �d�Xt�;��ғ�̘Q�׷>v�>���ڸ�S�ͤ�Ϫ.���[�@�KȬSfW��W�����9u�
               ���a�?\�Xg̭2�����?x����+�ū4�Lʀ��͕�ǵK�r0�A�ԗ꟯<]7��s�t@               �<�>��x��TSjd��f��_�D����ׯk��t�3�M�'/Y"��"dW���?_a�ܟ��{              ���(߭/~�Օ�e�H<�Y�<����M�'��&U���%u��ꅲZr?�>4I��;24���{b1�`4�*֙�[{��j���[��-�|��Z���k�y�������v��|�C���)��ߞՖ��              ��e4@��GNUE��\���50����	�ĎF��X<�O$�c�x_"a�U"^�t�J���mV[�Ӯ"��Y��9+�
�~�˪w��z٭V}��W'|�}�܍o�u�/P.f���Q�92���;��p�H�w]{����ښ����v���@��꒼y��y�ֽ����<E��g�              LPF���.?Me�e.:�=j���=0���ѱ_������GN��w?:��?3��:���s��`ae�י[�ݤs���f��?|I9�>)��XT�kϟ�S���]�c{����	=��}׌����Z���so�ۍ��|��*<��U���k���s�Ż�iӝ8Y7~�)�<�'               L%}�ç�T�}$M�~�g���������������|��&�{k�u�:{�՞��|���N�Q^Phɑ �;�h4��ߤ�j��O�S��,V.4-��7��ڲ����_������k��w�'��0N��k+��5O+��rز�U2:��'���<��G              ��W�s�:YU�y�~)�'��m�ݻ;�w`���Z�ӕ��кjU4���[C��?��$�w[Su��r�ש,�py��"1���-��&t�}nm�>yq�����z{�'�?�v(r׃�k��o�<_5���?8�wͫ/~oe�����w�V��{���1               w96����-+���	�_z�ȓG�F�.]�ڏW���\�=��͇/����2zi�5�]���ԙ��գ/��D3a�E>}��S'M�lo���v�����r���qw^��HrqY�uW:7��ܚ��낅�l���߫;޿R��)���              @�1��7^�Hsj�������v�����|���wk�֏_���������O�-��������;_}�|��s��k"���|�C����*�R�-��;^?��mW�~P�[]�oimM|zcՏn]�P������L���J�n�t�n���H      &0z�x�	y�q��	���.krݦ�H���O}�1+����vKBV�  8nƵ�p���蛿n�K�B�aU8&�Ƭ���,�u��"�Ԕ�      �M>k�Κ?-+���m�u�?��?�z��!M0w\s�S�ł�o>�����;Kggg���q?���^w�o���_ń��؛�_�⼌ﻳ4����w�r��VMp���;��������+=�zZK�{�.{FϚ��z����      �ƪ�
�	�b*�Ǖ���Hȗ\7�5{3] 0nF�}4j�pĢ!c�����V����&��     �-+�+���ge|��xB/�hߴ�;|�;��&�֏_�Br�r�=�����냅��ܿ�i���[��~��	k"�p��٬�f�gt��x\vtlڹ��_����jy����o����8�6�Ȣ��zK��`���ơ>���!      �>�5�wLW\~gL���#� �4ޜ}$�R�b���F,�[���7����B�      H���<}�%�p�q�?:8�򮎫?}�E��$s�G/�Akk��u?��)�+/��82v�+���Sk���{fB̨8��g��g4et�:G��Кۯ�������%�%���#7��Ss{�ϙ�����o� ��O�k`L      SY�=�2OTE��J=��2&�� ��+�|�1���Q�z�6��sԦ��z,.      ��鰩�=��se.f�ƴn�����׭��I{�筿�U7}���Λ^��9�%�L���a�թ3�_O�T��0�|�C7�Y�
Dg�˻��ٴ�{�WoXۣ)����u��xlac����L�����k����<�xb<     `�cm�7�
cxbrڸ6 �_�'Te����f�=���sԪ��'���]<"     pܮ8�EӃ�_��h����W�z���q׵�lomMT�}���V�q�2����ok�ƽ]z�`nG�'L���ՋTV��ȾFB�ĺ����_p�����[�-yҔ�y��Us����C��Jt��3��3o     `��Z��'�
�Wzc*t�  N�͒Py���1*����wa��Q�B1��      ����fŌ��o���/�?���׼w������_t�}�����U�)-�8ҽO�բ�/]�������V�������9U�WG�p���G�q�ի�i
{�9���~�w,���㴧���eok�;:t�sP      ��E	���ɋhzAT.뤝U ���'�PI�D�7qרU���7��aw     �?����/Z��EV<�Я7|���w���ۮ\��#_����/Ϭ
ҽ��"�.;�E�x|�rU��}.}��y�����#�nm[jt0Rn�|�]�{9�΅5�+�:�:���nM�`\����m�     �Detj7����EU��i�Z  ِz��K�E%!���t`ȡ�a:�     ��+�1W%��'��|�>t��Bʗ�]����jFñm�LK��V�T��lnӖ���E9p��y*�:Ӿ���z{_��?����~�g?��?��x�����O�޴N�<�H$O�G_�-     ����WCA89�r��� @.�*�*o45�	���ƀS#F��     `j�=�H�-�K�~��Q��}��rŚ�
����C��>0#�5z������ܗ�b��^�HW��+E��wO+���t漴?��M{��v�u6ߑ<0�?�k.~*q�#�N�]�|uI^Z�1�=0�
�	      �٬R�7�Ƃ�ʽ���׭�n������~v�M��^O~�� ��y5�����n�XF����y��Z�͋��pԪ}�v��w��     ��բ�]�(zN���p◯��ȧ?zѿ
ԃ�k�J-���'�>}N�)��WMi�.Z1C?xz�rM�܍i�?~�ܴ�g{[oϮ��-��n�K�z�ƛ����3L�T�O_[}�ˮ��6[_y�U     �<G\�
ê/��iͽP�Vw�\�x<�3�n9���p8�a�[,D� '��G"��cccM�����rddD�P�5����j	����mخ�}.�	     `�8Y���
Һ�p4�'_;x��csͻ�9��~����%����Θ�'7P���rI��ߵ�^��i��ގ��W�zg�y����u�%�w?�γW=�������%uz|�^�<�'     �\R슩�V]^$դ!ی�yyy���W�ϧ��2?�g�;��� �{l6[j���?�D"tJ�Ac98����Tg�l2~���ES�g̪��N�t(�\&     `��8�U�Һ�h<�������+�|S8f��>�eǯw,�Q6#]�����Y���G_Q.�ɀ��i��jN�>����zx�>���0.�]�z�힇���%���<��rUט��#oo�?|�Y     d�q�&/���Z�e�u����B��#� ��d L Ƭ!>�/5����>�������7G��z/rǵ�=�E�T����"q��     `�y�iM*���V߸�����+�|F��VK��{<�����<��4]�y��Z=��.�;�;��s2�~�I��d�����/|b��|����r�#��W4|ޚ�)���jnm�6��     @v$T�iAј���N����U\T$�ߟ��n�� L>�;�^UU��X,S����z{��ӣ��0>�I^GB�JB�����t     �GQ�[.oH�>~����7]v��q���G
���9�}_]Y�'�0r�F�۾��rE��=N�֞:3m�㉄�m9𩻮�d�pBn�j����w�>�zU��atq���O	      ����/
�ȕ� �ѡ=�����D%�ũn�  LU��Ţ@ 5���Sݾ��ݭ�.���f�ûӖм����°vt     �ĻO�)�Ö����t��qι�	���]t�{�c�z�u��rQ괖jͨة]�}�9p_��A�^g��?���3�\��.�]�oo�=2�:P���skK4��D��u	      ��Q-(	)��L���p���Le��*M�=�.� ��.���_�h��W$QWW��vv�ȑ#�F�i����3#�����~��	     L8�<�޵tz��w��6�m?�VK�ȝ�n�z�:����[:��t�7&~�M���F��[�[�:�����/��8[0M�Uћ����A�gs �mM�>.=���;     H�GL�KC��{���n�A�'GQQQ*�  ��xH���"5b�:;�q�HF��n[\KJ�4� �M=.�r     `"��9�Խ=O���_w�5�S0�'/�����~�����g���)�+UU��C�Cʶ�
��9�Z�����$^|���~xL0�]׭�����.\���t܌]�T���|�     �ٜF'�@HM��,J_V�՚
�WUV�:�j �<��~�#n�ݻ�t���T���s�8�:�|T3G#z�˭�PZz     ��i���e������CO�z���L�vp��꒡���<��V�E�h��ߤl˩��%'7���s�ۿ���Y��^��������JM��g��5���<��      �bUB́��BrX�l���Ju���s�r  ���PYYYYj�B!�wt�P[��ҶϠ'�s�iπC�t��t     ���5*���R��k0�y0�ZH�����}���n�,�}3͔�Y\���j�G#ʦ����RS���´��tp����j�������\v�Ϙ3�U�'^�H(�S�    �ɯ����2� �h�^W���< ��p�\���M���~8xP�JKWw��HCADվ�6v��ƀ㭏     ��է�n"��K��n��F�����ߚ�ȯnX<�l�ٵ]��6�F���[ٔ3��g��x�dyew���iu��\���������]��댹���K�     p��ք�B���"��|>��֦:�ӭ ��RXX���1��Qm�i���3}?.[B'���.?�;=���     䎙�~5&G:���s�-�_�U!�v�=7�}�Q�u��a��tpO��:cNUZj���c�W��!#��=���ʁ���
<f�>oIw     pܪ�ZZ2*���`{iI����U\\,  �ی������L+G�h���4}?AOL�N��^���8��;     ��jH=�&v�PȈ�?z���=��w,�}�ٵ��<�H��Q��D��Ԗ�TK{��#1�=2�>!c�N����ue�6����"Ք��@���    ���&��$��s'��X,*+-UCC����t:  �c�ZUYQ�]��ڹs����L݇͒Ђ�1��E�L�[}a��     +�բ��Ԑz���uw��E[��Y�w�C�_R�9̮}��i��u�����;�^�QȨ[�Xݺ�W��X[��3��i�c�?�m     ��(q�trpT���i5�`{Ey�f̘���< �����X%+V���v�RO��7��ΘΙ6�W�]��g�o��;     ȼ%�A�{���	E���.2�hJ}R�O�_���ڧ�T�?٤��#����=-j(3�n4W[��Ǆ��r��[�e�7�]��9��    �_dUBs���w���577+??_  `�Iݓ���رC�����6��/)S�7��z4%�     2봖�4�~e���_�v�^!�v��?���ݥ�S3�E�nͭ+զ��ʆ��W6W�n��^w�Ν�W^������?y���k���\f֝,PuI�ں�     ��8�:58��˼��~�_���TTT$  0�!��+��ѡ;wjddĴ�ިΫ�sn���:     0Eج�Tf�l�hL����⾫����?z���K̮}jK���/k�^3�Hh�ၿ�f�ZK����W�>�q�p     L�/���Q9��tm��|�5k��e��@  r��bQEE����<�7v�R86���ת�Qm�uhc�K	��     ���i���8L����[��K^��`��U����=NS;��#�}��p�Z��3̿9������/���UG�oG?�q�M�*�$y�����     �o%4�(�yEF�����6�U���jhh��j��  `�0���֪��2r߿��҉K�%V�;��;<��     �ϲ��	+����U_�amO�COn>�)8�̺U�y�,��pϰ2-����� N��������u_��=]syrϒ�3�.�^*�æp$&      ���*��s����>{�ly<  �7�á��ͪ����m����kJݠ'�s������l     H��i��}�{(�ُ��!�u|U
~���f���2ߔ:����KL�i��;�?%䄃�C�,����5]��*�ڼ�[     `j+v�tz���������2{�JJ̿f  &����X�\Ԏ;�DN��/�^��U�Z�����
     S���PC�������Z�	����-��*>S;�ϫ+�z���b�k�~����׼w��⍅��50�����-G�&O�     Lm��:�lD6�	��MKud���
  ����!j�֭���8�zV���lTgL/w�u��     �i���Ե3�	����3v����2�;�̚sk��z���-�7O�<:�_B�h]�*z��x�����̺-5�;     `��kqɘN�Z���ռ�sUTĵ  0~N�S�.T{{��nۦp8|�5��9^{\��*     �	KGC���w]s�z!gt�ޞ\�p/�w�"�S{�2)k���<xM킟z�{$�-!�t��(�05��\�Mg     �"��Ȓ�1�,<��]� �Y***T\\lZ7����|�a��ݫѨ���     ��3�:`z�C]/9�k.~�̧�G��^��u��M��{Cy��5v�|�ڵ{��2*�}�x�6�Մ���R�s������1    ���nM��QUz�'T��vk��*
�1  L]��ͽ��-��=��P�bWL�֯y51�     �zґ���<(�}��{���&3k�'��_�vP����{}:��C[��s���,��3����f֭/��k�Ļ�     ���&��bD�����4w�<9�6�   ����j��q�N����ۍ��a�zC��    ��z�*�w�Zs,U<�!�t��>�\�p/P�e-�>=h�_���'BNj���P^x��5��Ћ;	�    0�����FR]L���bь�566
   �|>�V�X��;vh߾}'T�mK��a�;�U�M      㑎��{�t�^�vH�9�C�{���ƽ1�L��%Y�W�Z/���X��m!'�FO.L�W�|    ����S�v�3~�5�^�.X����_|  S��j���f�~m޲E�h��k����o;�j!�     �ݴ�|�k���*��^{��S�Z�x�f�,-���)9����#k���gj�����;�����##�6�fy�+     0y�9�:�jD>��ۋ-\�P.�K   �PQQ�������>�:vkB�*���G���v�     L0�4d-��"/9�k`��"�0���>���@�2%+W�y.���v���r���^�lJ�6��<(���     �>{Bo;�p��i��2{v�{*  @6��|Z�b�^ݸQ]]]�]�jI���=��U!w     pґ��<#䬁����´���"yM�������Ccto�a�����Ӟ�)�7�Q�2�WV�E�DB     `�p��:�rDy�n7�F���  �
�á�K�h�Νڽg�qױZ�S�G��ݫ�sJ    ��'X�1�^,���J�Y��m��r3k�3)+w���)����;���=8�US�_cV=��"�ۡ�Ѱ     ����uvը
��n7�cK/V   @��X,jjj���Ֆ�[�8�&>6KB�ʇ���^��;     �ӊ�ݦ�����^�vH�Y�c����̬��3?���d�W��az͑Pl����G�{���B���;     ��Ӛ�Y�#�nw�\Z�t����  �ˌ�f<�^y�UE���a�JgT���C^u���     ��<���ݞ�P����:�kx�ʤ��������~!�E"�n�k�Nӫ    �LKu!�Q�����F�}�%r���B  �.%%%:i�2mx�%������a< X5������
     ��۬�������Bnk�1f4f4K:��NV�y�;�+�.!�E�	ӟ�1��"     �yƥ����*uǎk��߯�K����:  �X
�r�
��a�FFF���1Ϊ���ͫ�!w     �?|.�L�8����㻈��i]�*z�+n�ʹ�~Z��FV��!fKX�BNK(nz��ag�M     &��%c�ɋ׶eeeZ�p��V�\  `b�z�Z�|�^X�^����U#�ת�Q��ͫh���     `�r:��X��㻀��EL�;���攕��#���G����z̮�s�    ����֬�8�� �d�r�R!��/�������ө��m�W�      Ғ׍��CB�E�Fw)�Y�2ݐ:;w�CɉDB;��v
9-�v�]�I�    �	�6/�E%cǵ-�v  0�8�N��l�	�ܫ�Q-)ӋG�     ��!�����
�L�g��\V��ۦ�hBѢK�
9-;����&�    `b�;cZQ6z\�������y�� �I��/?�$��a�������̂�zǬzc����     `��X�OY&d�	9/��ͬ��c���J�=3�k&k�6�{�$�zT�Y���욑sl    0Ѹl	�^1*�u����Z0~�/�  d����ҥK�~����侴,���MGG3;u4     �-1s3�)6�
���v�f֋D3�\CV�ј�'��/��f�)w�%     �>F,}epT��������X, �  &=�áeK������踷�*�S�#z�ͧ�(��     0U���g,�6K���\���h���������i)r��j�]3�O�     �3�8�*ot��j�E�Z	h ����r�e���/(
�{{�=���G��C^�<     �T�����n#�>x�vSo���a�?'+����ob�%q��T�iv�������     H�i���������j��Ų۳r)   k��AF'�֯W$��%�����-     0����z�_b�Y�BNkmMX��ͦv<e6������#㿑��8�r!�9l��F�?�     �����V��&�����\����RK  ��(???5���_T"1��R�&X�cv��      S��u;��尙V�e����	>^a�ԙZs`d�3��,���K���BN��8�̮�74&     �ی�+�F崍/�e��Ra.����  `j+**�ܹs��k���+JG��P�F"�6�     �є���cZ=��H�i6K�4�k�d�!uV���K�������L�O$4���3     ��Z!�{c���b��B\~�_   ����448�={��{[�-����z�ͣ��    0���L��^w�u��U��BN�l+̮�?�G�GM�Y�uLrZ�ߛgf���1��㟊     dN�;�y�����بʊ
  �̚5K���:r�踷��j	����%     0ut����Ҽ�BN�Mz�Yr�9!'�sͮy�oD����{W�����V�:D�zB��Խ�o(�:Mm	��;,     ���քN	�ʪ�=�^YY���z  ���?�^X�^���x�}Į�M     `jHG��fM�.�9���nv͎�)p7�nI��"�i5K�ߍֻ�k�z퐐s���f����     �gAQH���������ܹse����<  ��a�۵x�"=�쳊D"���x�pEpL?=���    05t���v�˵T�Y��R�kf�)uV��=C��mV�������9'�k��5���    �\U⎩�?����Z�p�lV�   �y<͛7O�����%��ΘZ�!m�u	     L~����Z�9��{VQY��Ys`$������;QY���ВASk�;/��TU����{:�     r�ՒЊ�QY4��U��٩�   �˂ee���վ}�ƽ�ܢ����	     Ln{�����V��&�����M勴�XCW�Mn&���n���8a�~�"!�|��_�u�����=2      �{��U���̚�UUU	   �nVS����ԛ�a�H+����6��     L^G�GRݷ���jx��h��$WrJi��<�kN������l����'��x�sW��3��?�q�M�::�����i3     ��	8c��k����nn   ��j�j�z�g��o��wLM����9     &�D�ͦ�sk��S\��_�sNU����{�f�!u����'K(��a�ԇ�d-�#rYr��B�()�\bv͝�{O�o�s     �~K�B�����n���ϛ�Z  `�<nw�a�M��6�m���Ю���     ��v���p�(�rʧ�y���4�cv]��ɴ�ܣ����:sO���C"��S����Cl�.    ��R�Q��6������   �_UU��vv���}\�9�	-(������     9d�]r��5gV��o���i_��BN�{=�X-Sk��� 2-kw���ݦ�[j�[Z��ӂ����|?|������5%�?�%y�     ��a�$��$4�m~��O   N\������Q(4��d���w�;dެ�      �l�o~Sa�æ
��3��˄��P^x��5��V��'o6MV��R��8-������O
YWQ���f�4N�m{     r��@X>{��?�f�j������E  `�r:���Ң�_ye\��Ɩ���gm޷�     &�ޡ�u��8�Ժ�kD�='����S�
ͮ�y��G���7�9�p4.��jj��҂���{ֵ�[gov�-2����     ��#�f��:�655���
   �	��������qmW�iz^D{��     ��K���p�Q^���o<|��\���U%�����X�7�(�p7���vjic�Ժ��*[�����+/�)d�}���/+1}>�Y:Y     ���hL�q�/���Wmm�   `���fuvu)_����!�v(���;     �ы;�h�I���4��E�O'W����5am�^��u��C��ޯl�j����GL�;lV���O��.dMS��o�Qw�.�     �BgLu��O͙3G��    ��r���Q۶m�vƬ<3"��Ow     &��{�*��aGעc��>x��_y��7����U��;��f�5R�	eC���l;���3Of��\�Pv�w?:�+W_xPȸ��{�YՁ"��v��C}     �aAQH㹬SSS���/   �O]m�>�����S�[֮��tq    `�����#Z�Taj�B��Z]�wOru��sj��IG�g_oW�d=�~�oD��z�<��,��e�����&W�2�����t����CY{     ��bWL��b���N�C3  ��k�=[�=��㸯����hk/]�    ��~����wâ���Z�~ ���CBF}��Gn��̮;�j��)p7�fK��w���w������7��KȘ[�}�Җ��`:j���&     �����=��TӬYr:	K  dBaa����t�m|�VZ�T�P�.�     L6Ͼ~X�h\N��Ժ%����Zr�2!��Ԕܘ���ooO+ْw�+�U�'����
�NkMy���w	�\U�5������{���P�     @���c��F���}>_*`  �̙9s���+Ǭ;ք�
�z��%     0�]�_�Ѯ�Z̿g�xF��Z����ׯ�2���������t���k�mH��΁Qmx�C'�,7��ɳ+�k��ѕ�W^���v��2����od�/��8f�     i4'��7Ϛ�t<  �?��ri���ڵk׸���k[�S���     �l�xi_ZGI�����*!�Z�~ oYc����=8��ugSN�?ٰ/-w�æ�?H�N����<P����5�c�~��    ��+p�U�;���EEE*++   2�~�t<xP�б?�htq�Q��~�     ���Ү�:�7���kz핳*��������/���VŁ��*޴\�1�0r�ٔ3wcʃ��Q�xL�=�����o?��[/_}��6��Oण����     d_�?�c��itmojj   ��n����A۶m�v́�v8gv]     &�x"�'^ާ�5����Ms���_r�TH�۾���+�+�LG�����>e[�܍��c���#g�������[������k{�Oܬ�Y~Z��?�����     ���U�9��7:��~   {j�MӾ}�422r����qMK���?���F      �߰W�9�IN���ڳk�J�����r��� �ESM��v�w��^oWG�_CJ��	�~�����&y�濬��1�6�lr�Y0U��~Z����H:~�v�զ��     �7�0,���?FC�   �]V�UӧO�֭[ǵݜ@X���v�:     �z�B����$ga��TU��yf�vWie!��tD�!�lc����}��w��x�À�H��L0>��AY"!$��rZI�����U�uuO�TW�U�V������SM����ݳ�����y���ޏ7���)�������憛��+�i(��?���F���7��,Z��
��%����}xӅ�1>_z�ة����>��?z��@ƺ1�W���;�����Uk�a!�B!�B�:V���>�����!����B!��<�6n�޽{�J����17p,ٜ�#B!�B!��V6�u�m��4���]��r���o�s�c{��r�!|��o���]�ڬ���$�?�V���V����ۆp(@X ^}֖�&����x�[R7���?{�i�w7������!�B!�BV�-�YDTS��;v�B!�����[��SOz܎�,�B!�BHr��<~��!\�{cS��Xo�ቅ�����G�����O�Z$�<��_~�$Z����N�����+.<�)�k��v��������WN���Ǯ��+/?c�����'���9!�B!�B�ǎތ���}}��!�Bi6oތ��?�LF��nKW���"�7�͍B!�B!+�W�.ݵ�)-����O~�����ǿ��={Lu�������4�5�80�{�=�V���_��Sxݹ[mҧ6u�/<e��w����y��}I���S/9cӏ:�����/���!�B!�BV������!}����A!�BZMӰu�<��ҏQۺ�xj�i�)!�B!�BV�bN�^qFsZ�E�k������w�/����Ajb��[�:s����OZ�K�=�V�%�s)�t�^���On�k��y`d!�}l���={yw��#�ݲ�=4� ���8���B!�BH+pro6�U��靝�!�Bi=�����a��c;{2xj:��ŝB!�Bi7����q����My~����gm�6��7���\yH ���?���]�/h�k<��8z~�DK�-�v�Sx�ٛ1�k�k��st{&wۯ�×�H���n�8sS��-#��|�ʯ�>B!�B!��<�b⤞���Vh�B!��&�Hc��8|Dއ��8�l�ݗ	!�B!��r�\���~�wi�J���a���m��r����o�D����͟�|�Ʒ4�5���A�Ѳ�d&W����7���׹��u���~�����=�'V���뻞>}��P3_G��i��~B!�B!��;s��r�횪b� �B!�˖-[�-N��2�N!�B!��)_���x�Y�1��Rꡞ���]n�?�p����'@<�䗾��ל������;�}���x��,Z���[���~���m8}�@S_�glz�5߼������u�:H��M#/����i����Z߹{/�o�?,�B!�B�Zek�|{����A!�BZ���~���bffF�1�:��W�Z�!�B!��^,���¿?�?�yM}��C]�W���a�s�zͧ?��A�|��?��Ugn~��67�>��ƿ��I�"-p7L���|�W"R��Z/ߵ�������_w�K���I����u��~�I#m��n�k�N�+?�s!�B!��V!��X�)��e�fB!���gs����G�>?��X��P���EB!�B!���m��+�܄�w�6�u��;�o8�O#�~����o�7�
��_t�8s㛚��nq��l"�V�����s��O�_qZ�_��#'E��w����Co?��y�����-?]��Y�����=�d&B!�B!��VS����t������韏'�B!`���x�q�!�����B!�B!��?|�!|��F,�5�u�:����;�ڵ������s س�T���ދN]w�r��=���9�VeU(P_��i\|�zl�m�k��28��>�^���~��o��0����>|��G�[��ȏx�={�B!�Bi�t�}Æ �B!��P(���Q>rD�1~�B7�� F!�B!�����T���(>��g5��:�!�?^��:���W�?��+��Q�?��f���M'���;O۴nx9^o.�-R�2�"������õ�{"��g�7�D�����C_��������Xc�sϗc�2v��wm�l9nq`qxr���# �B!�BH�QM�������@!�BV�������9�_�B!�B!����y��Ņ��k�k�4�={��<6��C�|�=��k��_{ӻ.ݵ��=�e�t���a|&�VfU�-���u�X�
9sY^/֔ן�������k{n�e���7��ϯ��������z��5u��'�uiyÜB!�B!�gCG��g߇����@!�BV�5\4E:��~��.�wB!�B!��1M�o�� ����@��x?�����w<���������:���1վ�?��36�)�6����-���9�Vg��-�w�^��u��޸l�y�6u���M��ػ���Ц�����g�l��y;���#Z��JZ\x��$!��V��YLwT��vɏ;�*4�D<\�p�,zw�)D��;#�J~��B�z~/��Rƨ�H���J���
���T~�0̧��q"k"�3A!��6t���_B!���P�p�}��I?fCg��DE�B!�Bi_f|������D��^�z�7^����n}��ǒ��7x�a�)����{ֶ_]����|��������Up�>�Ė�l]��q��u�����������ؾ�o�����m�_\��w�����z;����O�|���@!�ԋL�pzwDAGȺ#���j ��)4E�f�����0��>��f����T�@)\���+ӥ��Y瓕W�R}�4����gߕ��fB����
�k��f,>G8����P!��B�Aՠ����o��5dMYCA*��uV@>mb6�ͤudx3B!��P�W5�;�.TU���(!�B��c��u��Q��@L�DJ!�BH;�)
zb
b!a� +� �Z�f� +�X��eW��g@-�^�뭔����gК3ET-q�j�P��3U~�0����P�-�l~�[�2Yʳ���n(Hdd�ߚU�5�2���x"!���<��8�t�c�ϯٽl���߃/>m�٧oJ���9����=��6��|wө��/8uݙ���]�H�s��7�Ar��VU�����Z?��s9:c�{���[Gw�������ѭ����g���Ǳ����ι;7u�#�,������} �B����J_\�`\A_�j&:4QE�j�Fz�L
�\�T� �(�%�_����f�5���tyV
����Z��i,/����� �(Ў����k-KJq�t�W��mk��\����f��������3��o.>W؄2��H!,�E�0�H!�15$ti]�t
�H���A7����B!��P�@D�3�
�:��B!�����G4E:��~̆��Bi)�2��}q�!a�k��������/�Ӻer.�_z.�l��2��`)���7"Y|��Oh)f����A0]��y+5z�&
6�U�ee�#f�T�0�P�P�e9���"gj�ME&��TNE"�gML%ML&�	B�Z盿|�n�%�/�|��b������F�֏^���|⪷܈U�;�|9v���/:u�]}�Qˌu������9�V��h��?q�}��;^V���r����37�fvg��o���}'����\�V{��݋���?���3#��g����~�TF�V�B�M11��o
�"@WHGT�A320s��z:��aŐz��������Ei�ƪ�����=��1.�܎�Uӂ9ט�C��ޝ�v�q�}�q���o����X~�o��m�jB�U�E�D�����2f9�'�7���A!��V6tȷ7����B!��^���q��A��;�<2!�BH3��������S�1�X1EG9(��z�t�t
��%_1��Z*���j���*K�*�n����|y(�k�p�$
��sn�Y�y=��L*Yy�Y슏���ͣ-?p�,d��,ܽ1��B�
�`���-op.�ê7���7H!��v��o݇��/-ݗ�S7��o���;&a��y�[���=�������go~�X_Gd�����1����&Ve����g����>x�9+��=���/K�s{�~��w:>��O��O�����7�~���:���!u�? R&������&�A!�=�*��c5���3�bj!33���I"�J��SjQ\RX�P��uk�D��t���qI(�;�����\y�q\>�8���w� �`��8�;+� �^5���t2��2�(?�
Z��b��n�X�_�B�!��0�u�I�Ь��d��E�Bi;�u�ܭ��	!�BV5���cVa����r~!�BV7a�q��x'���3d��a�*�JCϦ�XX(��+P�-Y��;7g�
1���
���Y����qŜ`M�B,ۚ�o�Q�U�o���\�l�2o�5:�uX�`���c&"=D���ݢu-V§�׌�i��M�ӑ�=H!�+�i_���1�ױ"��b���]����O�����˛�-̇>s������9g���c+z���b����j��}��o���:�!�]/Νf<��柏�=2�oG&�?�>�Sh>z��F;��r�H�[G{zW����о������B�������jAp�	�Ur����$���ֺ�Y����%��P��s��֪�ν[���<��׸�h�b�c��`�m�)\��c�\�����¼�h%r7���������x��Z%�kC�D�+�H�j8��ł��������!!��DTQ����tw#��B!��^���
͜�e�����p'�B����`c���.�/b n��s:�T*U8OɪPf�����~"�c�2,�W(
��=��.�
�ʔb��nEYw}v-�r�ߝk�ݢ���ߙ�q(��!���=@4G$ڑ�MFN� i�0��pl������ҢL̥��ޅ�/��;^��������_v�=�ؾ�><�����+�`����8{պ�����ypg̺ Za�Y,_��ꀻ�o{�
������a5���uh8��>���S~�����N���o?��������M'G��{7�t��i�ևC+��2F�b�o�}?�z�0!���a'��� �CYD���M!��G:���Q��T�V�-�^��6g��j^6��f�lmw	���cѱ�\ðO�)��X4v���Ea��̱m�j�c�$06���`��^2�!��5_��p,�bߌ��\��B!�1�!{���vB!��Տ�i�����c�c9�_�V#!�B���l��R1ҥ` j�S�6��&��X���Ղ�f�E~�t)�WI�_��/��c�oh�w���Ex�����7t�Wy�h�o(����YR������[�i`g��X<�XgW�>m�0�a"�60�a��BV�����_��杗r�+�XGx������_v�3{�L�<=�������>޹�˱m���h_��N�v�?x�Pkv�������_��W#m�:]��� 	��قV�+V^�s�t�ħ�9�������{hb6}�����?~�l#_��|w�P\������8�}ڦ������]Xװ�t����o�BH�a�O[��Fv}V��������\!Įd�TzYPR-����z��]78�kp;v���u��v�)H��-��Ƞ�3��5�p�{߅��c�@�mξ�ލEa�~O%aZ�������X�@�3R��p'�`<�bߴ���	!��F0�I�k�!�B��gp` X�=N�BY+��	as03G��B&�D*�(�s���R칠�X~�!<J��ʰ||� �X���ߚ,n��hͯKt����c	��*�B�w(�&�f�����Jw��7�#뀡ő4#8��p`���9^�B�r��I|�_�§�y	"��������s]oo~{G��������g_�I�6����'�z�Í|���!r�X�-����_��y�����x$�Z�],���V���"�n]���w(�[%�^�jO_��sy��r�4�����dO̦����s��Sɔ�h��)9�X�B���O�緎X����n�Vԑp8<�ARUm[wG�̮h����躑�x�@W�e>�!�
�]�����{_ !���%���>��N]�,¹$��y$�I@W��C��E��b/m�av�M���ã��)<�hw����cѱ�\-�Xx�Sn�E+T�S�9�@�h���O�����^��Җ�Zߍ9(��P~m0d :/�����S���a6�:?�J!��#�a%5����B!���	��E��5���-��B!�Fƺ5l�Q07Сd��)��g�Ng�.�@BAjџ�t�*/Q�3���R,�P:�� ��k��\?�ЎlIV-�a��X�w�0;$�C7�P7��w�M��k�s�C��;�F:�DS�̘84k@7�BH����?��_���Hk�W�{���vr~hmW���s��ɹ�љD�d:�H:�}.��'̜q"m�Љ��#_��ԟ~��C�Hh$�P6�5e �����l���uD�\p+c�ۭ��DZ�Ъi����ՠ���<��To�hZ+8���o��Ck;Wt��?�(�����}�A���} ���tGU�P1�Y��L�3�@ƀ�U�Q�-
��.8��.��k��#��l�{����kα̱�|��;��	�;�A�,�h�J P��9�81?��OCˏG��CQ�����H��X��ϰɁB��/o�r�V�ݺ~$�B!�����B!�rr�C1Gmc7B!k��'�����) �@ra.�CM�P�
�6O�d�W��~�X���h!�'z���A���q;����z����Z�� �wi߰�M���Kw�N&a&߰'|�1*�:eFp<�s�:����͖BZ�����t������Z�����ߺO�����o����oi�̮����}���-�Jq���>��G������
��d�:>y�����@!����Ul�+�ٻ��������T��U��H$�`��PNAJp\d�m^����~c�9���8�X�6'��WCCа{#��}-c/+ж(J	��ǆ# �����'���0�]0�]��E�xa�-�B�n�$3� �B!큥m���c||\�1��B!-��ʾ�?�>�!�̒����L��;;[����
��ʰD��L9V#|D��לh�7�5�9�?4%<*/��y�h���Q~�W��7\�����x0?71�Y*ǚ΅px����\�ޝ�B����)�ٗ�ħ��b�wEAV���<��}ý��n;Ж�ӗ~�O.�_qB*/<V��d��ƣ�&@!��Xa�S�4�F���H-X�LAM��0{rQD*��W�݂�vAJ2Ю
�-dB�ݽ�d���E�ns�&h��~,+X5#�$��6_��yA��jl?�1�N��\�C4�=��2B��z�'�<;i��\{\�B!�����p'�Bi+�0	�Ũ�B!�D)�>�!j$���A:��:��P�av���(��vg����Z�e���ߜ�Xt�7�܂��n/�z�A|C�p��7���B��r,s�%�p�j{�f9!����Ӹ�ڟ�Sx���?��E����n���V[�-nyp&�R���}):ca�����<>�ջp(�'�R�bb[�қ���Zfr�Ш��)�.����X,^`�
���U�vQ�]-Vy�#N�"P5"��*J'lk�Y��'@�0�;S�V5o�1������d�)�\=�w{K{�p��O����3�����x��R���d�7��򶅄Bڗ��\Hɺ����!�Bi��@�G��B!+�h���*�#���X�����0��.5��b1�B,�2,������9�2�N�	����փ���k���m��G��7t�c�ܯ����P'���xvR����	!�ɱ����_`��_��NY>�<��?~߾�9�mp����cxߵ?���~!��!�¯�>�O�x�YB	��U!f�c~z�n@�ѐ��P� �_��)H�lo�8�'P5F�*|��[Zp��ƕ_���Ae�����).��5gؽ�xI���ī� !�ZĪz+_�E�r������}���`L`(?���DGg�xf���Qx�BB!m�l�������B!��=��]�/TU"��i&R:uB!���U��!��@R0Rs����:�!����߿C�����w�=��z<D���eB(uY[Zw�����*��[a��cY~��Z-��Ҿ�`���aw�oXC)Vi���͟?����9!��r��ځC!<9�C*BY�X����+w�^��w�� �g6��_�p��ڑ��[<1��_{;>��sq�� ������;��o}�pH!D��!l�3Ы$���F*��VhUА(QjQh��{�=�)��%VY4C�*�����$���Ħ��űR��l�9kns���a#L<�Z�2�sf����̥y����岗�jia�Z���֜B�0�.���[6���:��ޠ�ԡ���XP:�oN�S�Y��BY�����ވ\Qoo/!�BH{��*:::��� ������ɶ�	!��eeK�{��P
Jf��@F�2�")�ó�OT�%Q�%p���7t�#Z��+|��;ז\��R�X��+�2�:#�U%Y���X���p,(�rY��+t���~���"��^�U�oX*�͏Ǻ���>��.Le#xvJ��&�	!k�0q��?��L�CW��X�EI�������_��T�ʚP�����7��=goƟ����C�`��$����o^!�o6�j8u�D��Bva�D
ꔊ�b(=��"�@��0����#<5��=P��x��/�
�b]fw�P��zU�]�IKU�AEH]�KM���y�LM���e�tQ��ۃ�n�w�9���iz�a��5�\3Zj�K�T�}�|�X�:�o��)���F]��v��}Hk�8��c9d�cBYt�h�ܹ=�� �B!�GoOO��{�wB!�^,q�@�}UKC/x��;</�w�H��;��C�����_�ݹf?.�����[���K�*�����EEY�	;uW�;b�",ۼ�,{�+� �;�P�+�j�w(��b���+�y�s��ǻ��B�{?���U��x�4!d-��Gb�|�m�c��>��a�e~��{�ٜ\i�jeM�M�>�O�������o���B�DSLl�^�J��	d3Yh�V�]+�H�XLf����#N���P\p��u�r�(�s�y�u��5{�])����|�u׹��ŧ�Ƭ�">G�n.-���Ax����ι��{�~I��U	Y�q=A�~P���ǂ�{�897�?��P~���^�H���1ު�BHk�ѥ����!�Bi?���G�H��5A!�y4E����!�g'��d�N��@���9�٥�C�^���z��^/����v���/>��_��/�U�<��}-e��|F�c��8�.�z�a�k���B���/��E>a�k��l�o'G��CR���!<5�C�y��Ҏ���U����T��?�Z�>!�15��gnz �<sk�5p���м������N��_~
�!�Z2R��B����� �����0N���e�ca���mZ��*p)��l���R2A�z�,*�C�Ő�G�� P�C�g-�����B����&?9.�����#�k�9��!�5�6�7����5W��e�|�
�/>�,b-�ŮF�1x�=� !��c���N�Ø�-�/�����
�`�\O�@gk!���/"��`]?1�N!�Ҟt����!IB!d-b�b�:��]f��	d
�Xb���=B�A|��5�[�z�c�B,�",_ѧ0��R,�1��Eٵ�ؽ=��Zʱ����{e��7�n�	]�l~a��z<CO�P�7��m������I��Bx츎���;!�����'�������`�0�\�{��õ�<����)�^sw��n��?4�x��􊳱k� �k�
!��1ءb׈��P
����$0a5��д�a�*��)L9ũ �� A��*{ �z�,49��kp�+��z�}���5�q�׼��������qNuнJԪ8�<_|w��ͪ���U%j���P�[��|������k�42ip�
�/�Ǝ��H�rΥ������ul��XON���D�B�J�%p�F��k�0!�BH����l����	!��Z�ܫ���bC{bz��eR��/��������n�bE^��G���>�Ǹ�3��W{��u�|C[Hݻ��x�9���P�	z�y{�e߯xP9��/N��Aw���
��л�Oq��������+4%���ݠ�0�xu�Wh5�?~���&�����{>�3���O��]v
B* e9<�����C�	�5�d��ľ�������ڀ���K0���γ��q�S�ˆB�*��;���6ųP3Ә���:c�]`�U`w�KRA��T^�v�|Yh�X�Mh���"��x��J��s��c����W�U� 8^���V�9���A�KbW�\Y|*	Q�/�9��*�+��� �h+=�Q�hd4��%\U�6�D�������9��\�50��QL!dy�
ɽ�ttPC!�BiW"�4U�n�]FT��e�ӄB�.*v�J�&�L$�Ni�R,U����=DE�����
������%�rNX�e�+��j�����Bqٕ3�.w\9W9_�&>�6�����
�� Ǖk���⋉}B�\E���:K��J��B�~�w����X˰ܼ���Fb���x��^!!�m�du|��O�����j.۽ĝt���o�|߸�idrk�}`M�-�����g��헝��\�Ѱ�ĉ�$�������_��"�����C!�ܫ#n�bnjX�_D$�"R�%�^�ك�"��C���dE*�P;��$C�KBՒ�T����}�k�^t���׸�c���s�GD+� �����|I4�r�
��E�ҾB���_�D����{U��?�^�`U�pe�D"�s���\٩���u\5�52�\�/΅�رt��1!������w'�B!m���utvbnnN�1�!��5B!k��
�2�����R,)U[,Ŋ�U��l����7��s+����v��l>�T!�(��]�%���z��Kߓ�� �Nm�X����q����U����p���R,Q��'t��Ω�����%zy���d%���Ӱ�B]#�0"}8��c9dX�NY�<1����{�ғ��������%����<| _��1��Ma-���%��w�/��8n�ճ��ғ���@���ff!��|7��ܚ�!dmb������vf��sЭ[jZ��H*��f�%�^�HU!N���Łw��Q�&
�/���Seؽx�x��<�s�sn�n������Տ3�.��jw�,q��z�+ /ދD��^�w���w�<6cQd�	��d��^�Uզ�Us��<��Y���6��Ąى��I�BH#�1M.�g��B!�����$�n}Pr*B!���ҧ��!]�,�'af�&5V)V4Z� 5M�˯K&�^O9V��Q���5T̋����?(�Ek��Z����)�p1VsB�2�X~Y�X�`՜�V�%��
�aw/�P�����	��2t��GCW� �n<vB����	!��{�9���=�Kw�ǻ^����������y����'�ܑiܫ�Idp��?��޽o�d'^w�VtD�֏i|6���z߿�y�2LB��*�U0�. 1}zRG:�n�+lX��$��JcUN�r���<Ghw�{�ճ��778ϩ^�>��w#��n؛j=�9_ٞP��fV�S9�
�{�Tr�����K��xe��o����F����RM�.BVb�"�1\1�5<�t�ON���D�BH�X��^����	!�Bښx<���0��!��V����rK���40�!���B�$�B%��������p{ �j�sNT�%������j����2�~��>�������潎k�y��by����/(S���\
��۳��X�oX�u��)(�N7u���j� �'��͑��4'��"����!���a���M�򒓱m�5�����;�?�o��4��Ybm%�`��?��G�՟=��>�x�v��V֧>n��s��#�3��u��Z�1���~��榧�N�A����T�]��D��F5�WRj��f�|D)���6.��T�0�S����v��Z��=W�f��������߽,��.f�"R�߽�~�l�]J�4��5��]���C�K��QY��t�B��˿ot��[#!�BY��@c'�Bڄ���������G&�.����q�7��^�P����;��}=CQ�]^�	�׶�����m.��r��)��+}��W�5�`�h�~�����=C�B,�&.�*yx��XA��A�n���;�e�0&��_;�;ABV'V��և�㶇���x��;q�����n�YHeq˃���ñ�H5��0��M��_>��|g�4\�_|�z������H��'�rxp�qBH;V��ׅ�)�@f�2�4�I)u񶁚V)Jل(-�H4�.'J	��a�B����E*g(�)L��J㒈�?W�&�w�����YrN��݃��e�dB��q���h�t��D,	���Ʌ�����+��%
��r�����>}#8�w��:2�B�&����b �B!�K<��^\��@!d���Wîa]��&��(H�E/0s	��q��F�ܫ�C�2,A����h��ʗ`y���(ƪ���y���y!�8Y_0����݂���{�Y��d��
C��z��B7�0�_�V��8g�	:j�NЄ�Չ�W�}�+l��37��݊���)^z��4~p����#���@�a�]�B�
�[�`w��ސ�6b���U�)�l���p?� �~�(��BښH����6w���9��BɤVhi�B9%Jl��Tv����Cx�;o��T�t��m��I�W�L�c�9�9��ZƵ�:��F!#f��ڝǵ�+*��{�л��%��HUja���D,�<o�ۛnw[��Z�EA���5=��(.� �7c�����̦i:B�&�ʷnZ%�B!�K$��^�wB!�E1�k$���Y��H&�	IMC$���P����B�OP�K�K���b=�X�>�!��(f_�p{=~bа{#B�~�bP�Pf/xt�op���b�*��:6�������wQ	�K�]�͕��=|Ɔ.��A<3��v'��>�&��/?{_��)��s��׵ʩ;��/��|�?z��ٵ�D������Kᦻ����8.>m=���:k�0b���B�?{�<s�<}i��	!�K,��v���EHN���#�ZlY��
�va����.ѼPk���ցN1�~�ڃꮡv�M��&H��굼�n�ZE�Z�%�n�OȒ�d����㠂�нz�v��W����ұ|нV���X�]E+]tl'f&5�񲘁��$"���0��[�B)�T�B�Њ]B!���!�:?�R_ ���h��3�4l�B�'
��t���bq�",��k�ӳ�]���-����b-��⠻��Y�b��
��6*��H�,H�=h�=�_�<�u,�����B����y�~�X�A���v/o�*�������tF�6��v�Ơ���(9�� ��!d��������G[�{*��1�����v�a��������80�{�)~���	�u2>��w����C*vo�[��{� N�4�xde~�V���}xt�	<��	<wd�p!E!�J<��uj!Ԟ�<c�(�,X�O8�nZp��۽B��!w[��j��&Q�]u����X�Z�*[��B�[��*H��Ya�Z��+���c	 �N�=侜��hι&'\Ʌ��,�ycQ��WF�q���.b�,GkC��z	ZU��v�%�^�怹��ѵ�v蘂�s:!��]��ܕ��	!�Bڟp8��(�	!�� �b⌱0�u���G*�F:]y�g��������9���"��j��ay{�~>��S���m܌@����M�e��A�B�|3��Z��Aw�?(�����r,g��t_Zw����g��j��
�-;q#��7��ƑL�=�C��]%��0ٜ���:R�,6uᬓ��{s1��R�w+���)<���x?�%���b��y����f�����y��F{�}]_a�~�c}�0|#H���Z��sx��la�>�qxr���tET�t��e�'�YB�Z(�HIp���{�۽�)�US��.Fم(�XdW=Z��T��TK�]r��]�w,s\�+.���J�p{�d���������A�P|���f�Es�8�^)f�D,�he~{#�Sв�9T�5�R�{���oC�Gнj\�l�&���g�:.�2��P?8�`|�awBYk�49�"0�D!�BV���Ȇ�bZQoqQ�!��e�j��G&�F**x�V���;��A��@ޡ_)� ��ӳ�����z��Av� {-�ߜ�8�Zй���IhY�����?��fz�A�B��{�r,Q�������s�a--�n�a���ŽU"�m�x�`�R�������BZ�'�����P8�a�X/N�oV^���Zy���Ɣ7Y��'f�8<1��[��<���N#��'��M���\
��쑃�y�w�;���8z:��?<t���G���R���h�,�Kf
�LV�\*�م4fL��Ǧ�1!��%,Q���al�/6�O����HYd*�QU��8e��ك
U"TU��.<�ϭ��	O� ��ze��W��"�>�Z-c�qa�� �=�V��pCZ��E�r�G.��+X���_<�tY3������U�w��X�����97{˻g�]$^��*E���g�]6��K.�Cї���B���P��4��B�Z@�u3�wB!������"�������U��BȊ`��箏`sləcГ:ҙP�g����ޡ�Xk!V�R,a��Q����^[1��g�,�o�����m��V<^T��b�]���kz.�x_�����;�ޘr,�gh���6��ݱVtX���:�n=�������8>�?הӏ	!d%��K���=V1��0�ׁ��z:"�툢+F<Z�PwD��Lgr��F��`>��L"S���&��Mb|&Y�������o}���!�����A~ƘVhZ��Cv!�d�x�@�d��L�P�W��k*TI��]D)�0�� UZ�Zs�������mέm�w^�V���F@��{��%p��=�ͪ)����Jv/���W�w7��&b�ir�γ�W�M����SsЌi\���ً����Bڙ����6OB!���X�}�w��ƀ;!���eǠ�����Ez>�D���b�@�X��w([���.��]K��a��yR>����oݯK����	�{�؋�U��^�Ң���z�9�{�������������
»y����B/O�o�o�+�9�?ق,�]�EEY%�*�����@�9���+���zh���(��so�"�;��x�h6��-�aB� ����㳅���HBiY,Q��~��1$���
���
U�*�2�^��`�\�\�,����
�����(���9�X��{��[���B,r���y	\vAH0/z.�����լ����K��W!`���M�}�F�@[����0;��^ӧ"�?Z�-�d�S�"���BU�4U����B!kK��VP�x�H!��la�@Zb���'��v�?��;t�E�`M�v��t��+Ū�+x�=Hx���{��8)7�5�&��s~�2jG������J����)Ò���A<C�sd�����s��dU������b�*�0X�]f=P9�c��8�����c1(��xx"��r �B��BZ�����I����r�!�(%���{	UKk�bT�%�;ŨF��D)�F	R5ڋ�c��TS��-��p_\��d�[!�����ye)�M�����B���p��"��9�V�W4�L�*	J� ���aq���
�;[ݭ�u[®\o�C���<=N�B�U��G	t"�B!���w�LB!AY׭�Q��)�MO�C�T�%��[���!�B�Qx�+����<���X��s����K'+������^>���c|���as�kz>��'�?��ceʰ�ޠ�M�kI��^k�
���2����X
�W��;A��>�X΂�z��@~��>��?f� N6r8k}7�C�暴c�:!��F;!��'�7�pc��,f'�C�P�)����@�� Uoc�S�*�-1Gu�+�[
���T�[�����%H��~Ⓦ UK���@�St	N"��)z�͋ϭ�V�v�"����y�g{�Z"1Kz�[~�w���~���
Y�Zjog��+���K{�hUo�]Z�ͅ���HO�V=��ū���H�^��Z�$/�4�	!�B�A��4u�il�BZ�Ψ��֫�3�0;=LhHi��x�=J��Qޡ�oh��˱ľa3J�*���{��Z�Uw�����e�+��LY��9N��k������f�Esr�aP�Х$�����c-�_((�ҍ0��4��~�����6�	���&�Y���B�wB!+Ʈ�N�M#3}���(�
)QȽѡ�ʦ�@{EÂH�rIբT��
V�-j�)D��Pu��+�6��$�rZE��KdQʿ6��$��� K�xQ0�3��<�	�;���,���}��Jf,�� ތ��E�kȽ ^�x��~�m��wWUs�������!3{q��rԮ!dU!۸�ɓB!��N7�C�z�B���O�I!9yƔ��J��Y�;���EX���7���C�2ޡA�E�Y2k��A��~��<���9)���C�-ê�c���0뼴�`�e�J�dʰDs�����ߧϾ��XA���EX�aw�b,{�=h���gX����Uw���FD��+zT��G�b��濏���BY)p'�����T�t=Н=���Y�&�����ea�qJV�Z�J"�(��#R	D���vQ3�E�P{�w�qq��x�%@9%/�IF|�<%���3���&�M�*=����K�x�s+E��H#�;C�N��X(f	ּ�+���w���л�^!8�����"�3�^KSC�s�x^bv
�	�a8�{O���d�BZM2��0�N!��&zݧ1�N!�Fƺ5�7�#�p�DɩP�ۋD"�eXn>b�@����+PS{�R�꠻ES����.ǁ
��u?�P6�n���3��F��~�[_�=XQ���Y����Uޠ���A�t��g��Xr��`A� a��V���-��K��Ɖ����pź.�Cxp\���BHp'��t4����������Q(S*ҋ�v��v{Ƚ$>9(/A�O���D*qۂ]���WTn���U�
ԮP<p�&��Ϛ����4",=L�Y�Z	x��s����b���ʊ^�w����,vy�.������Dw7˹oD��y,v�U���W5��45�v݅c����<�����ԇ�� ~u��B�f7!��*��9��!�BY��0K�$�Bd����ׇ�>\��I9��?�
�{b�|���K���:�����9����W��Ƌǵ�k�m/U:
pn�*dh�W����~�l��z����}+�r����cA�}��cy���=�V�*��t�~�g���+�
��B�@�m��p�)vcB��wB!McK��s����Cv!�D�jZ���+�)�`{��5,D�%1�[���d���E3�����`,j�M"��Kp�
��E!E�Z�����J��Ur�v��T�O��	Ż�S���b��Jl�
���i��6J�jdؽR�2<����%�Z�rXU��R[C#�e��zy!�L@���e�
:6��Ssx�X�BZ���h?���	!�BH����i'�"ÎA/��!7s��,��?\�`���U���;~��/��}��ڽB����縟+��y����}�{z�~�wн��ޡLA��?�r��.7*�^�7�˫�=�.��Z���tw��3��xU��h�������	!��À;!������1y�z���>{�(ғE�)j�-8)Q��!Hɶ���U� ��(U�*Ũ�}��$
���-�p/��s��*��� ���,��x�9���V����7��ڊ��U)B��Ĭ�k�V!�6����pwWT^!�+W
X>�U��/��K�r�V��P(T�&�bC~��B��]������
��2 S�i0�N!��&z�g0�N!ąΨ�K6(�L�ca~��P�۳�څ�v�b�Z�����^�%�!z��[�K2��^j/?s��������~^XU����eY2���<:��,�f`�PQ|��`>aб�_������VwY��t��V~�3��;����#ؤ�p��>L���&�Y�΄B*a��BHC��p�:��1�����h4Z�dC�v�I&�.��C�Ά��H����dw��6��Ū�|\�/ι�P�S�Av?A�/�.+5>�n��~��H���D���J?/w�M,���.�|��c}�����`,�7�s�$�.+X��J⑟��r/W�-�.hk(�[ZdCg��!^Y����.�V��c31<=��B�JbH�]�|E!�B�pיG!��`�@gd��>}*��B4��{�ڝ��A<Ċ5E�������;<;<�z��V���;����<(7_�-��`������]��ׇd'`�<O� ��tԋ=��\鑐��ʌ�����C�>~aɇ�)Ʋ���	�;ׄ�"�Pv/̇�J&�����u�	!�T��;!���Q����&���T����m�@�W�H������r�}�i�l��}��XtA�p{�gԘ�{a_<�
�{�M�(�,'<y�N�b�L������g�������[X�o��d�Y�\�������)rn�V����A�u����/`���e��)`�ޥ�*A����](^-�4l�sص����~�~)jW����������wB!�����o�@�>��BH{	naT����r[{4�*�
z�g��vg���7��ٽ��ܘb,�F�K���t�]�#V���U̕G.�kb�I&�����Z�e<?ْ,�c-ޡ[����U���w�7X���.w��pWUk_�_�����rн��|����
��tq-D��B��	!��/���Lt��#�0�D*�H$�f�im�	�ˉS���8�liث������W��!��av7�?�4�^k�}����$h��� 'A~���k�BU�yq�J�r
W�9W�'�^��p��w668E,���]��hxw�ݗ����{�!w{��+�^��Vwun����_���G�&��N!�v�� �	!�B�F@�L7V��F!��l���,����L�-��J�d�����|C�B,�b,wqJ�dC�>~bc}�ʵ�^��kʲ���V�������0|��skg��;tΕ~�}B,O9V#
���� �a��ݯ˴a��	Z�'|h�_��0B=���x�~!!��Qp'�"ͩ�!��I`~��)Gۂ�0�Ӹ\�r�P��
B�b��0U�(T���B�W��O���{�O�
�7ShZK"V#~��� B� ��P������A���fq�K�r�J{��{i_o�]�� ��\���{i�5��U���л]�
��-���8:^�m�3}��p&�kh�:!�T�K���ks!�B����}��N!kMQp�z�p���G��,���X��/t�e<C��h���m�b�P.�^z���b�b�+����y���%Z,��׎c�ʲd6b0x ^�#,�U��nw����"�z�����z����*��z=C�b,��
�!w���.�"�0=y��^�m��~ܵ?��W!d���;!�O,a��M�kS���@bJC8^�B���v7�JV��;C��R��`Ws�P��],JY42��/��E�T�|�������yy��]�r�H��Ĥ��~%:y����	�~�Z��	Z�߃k�C��}Ѐ�ۚ��%���W��+��.�� -�^��-�[rv
��q\����QܾHf�\BH3�%/	ҙ!�BH��	x�g��:!��֠'���M
"s��^H#��J���J�Dޠl��������ڽ}Cg���ؖ(�jH����{�^�E�<�V�W�Z�[�%�Z~�_�c��;\���	������?εJP�����R�%*�r��aw�B,/�01;�}���߄�ᎃ*�S�	!��a��B��NK�ڠ�3u��$��@�x����R2��^b�(��lmwګ��m�BTu���M���Jc�x<؎j��[p�MA�4Bj�����f|����e����z���{#Rq��x1�n�<��X<�tN-���w���p�lg0�D�JQʴ	V�	W^awQ��K�*�4d-S=�"^ѫ ڿ�>��Y6BH#��;�M��B!m���n��=i�wBiw��p�`ɉ���	]��˔b����fw��v�v��>{o�V���!����j;.IΉ�ۋFy]+�����ѥY+Q�����]|��kP9�^�U�K�K�z��=Cw����S�U�ݟ����^lu�'������t{OdA!�=a��BH�{5�;�Cf� �)YK���7&�nkd(�P�x�J��	����)�@�ŉ�����
Q�"���P�h�h�g5H�NПaPA��f��i��l�T���:�,�Ɔ�~��Z�+籼xe���X�r���~��2�Uy��\���a�D�q�a<���o�0�N!� �˽�gp'�Bi{��`!���@g�"!��-g�aG|s�Ǒ����9�w�G���J��C�2���$ˢV?ѾV�Ń&{�K�ιz����w���֊�؈_g�!�Fd�[�U�O�<��8X9V����q�й.�	�<Cw�P�˫���@{����#ؑߟ�m��~�u �����[Bi'p'�R� Lu�c��Q�'�BS8$L�����.X{�&:��^"�P����nXO��|^qЀ`{�k���r��k>V[��Z�,���(QJ��j�=�%������/�Q,jW��]��ڣZ�
"\��5�	W^��"�J,bم+�`��p
���Sˍc��^L����}:�4�	!�fd7�����!�Bi?��t��u^BH�)�x����1$��Ȅ�D�
�/�`)~�a0�P��"��X�+Z��Z�ܝ�J)V+z}����K��khdAV�ʱd�K&��5WU�UK�=�W(�s[��	��CgA�o9�O1V-���f�������	\����QܾH�0$����wBYÄU��-��Ǳ07W�*n#(�B�����[\�م��]��R�	��V�y�~���fo���V�Z�ZF���<��8%�J����!��_���aq�+f��n���ܗD��vww��?��'^�-2�v_�$X9���|&�@$�<^?A�s=n?,���!�%����=#�!�BH{��]�Ò�BZ��.��0fB�֑����54���>>�"nk�mm��-��S+^�UK�}%K�����F�Y�s=��Fd5�����y��� ���2��2Aw���Wh˄�E>ae�U���Fc���z���G�/�=*��q��0��1�N!��	!d�Q���
"s���J#�����b��@Z\�%��u;A�G������	��	V���@��
�W�_��_���;̾��+!,�F1KD�d��d����{��{Q�Z
��ķ;�ޥE����	�{�ޅ���@�@��VÂ{.�i����>\�	�6o�]G#8:��B�� ��T:̀;!�BH�J���wBY��:��y�OEn�n�~�X2�v��v7�P����u�g�Zi\�+�1�.p�d�K�X��:�٭DA�j,�*=u=��Z��^kK^a����+�����X��a1���8��B&.޾O����BBY�0�N!k����7���x��b�bh�'��lnw�j��o#轷Q��9�^�p��
���'o!j9���
E��(`-_c���ts{���_�h����m
{{��K�j|�=�he�t��e@�+E,?�JZ�r��C�!w�}�4��8��4];�၉�0�!�o���L&���!�BiO��{A`��BV/g�aG|s�Ǒ���D����vY�P����n��o��b,���Zq�R�:���h��Z)Q���Y��ˍ���3�n���+%j��Q�dz���qgq��m�_�5]⿪��E_�=���.}Ӟ�N���b7q;v��E��$J	�  ���3�w�ޙ;��|���w@B0x�����x�}��p�
����u���w�=�KU�e����Aw�kKs�`��3WO���靻� `�@�  � ���S۴�x�����^�B�B�h P�	�+ũB�+0�����ٝ�!bQ���i�Vq�&q�a}|�Z�EL~N�Ǐ��%N�	��BV�<c�Ƕ�͏)����ʦ��Y�]&`���>�J�lo/��uZ�����*��]"^9���=�Ӥg����G����  @E���kx     ���Ɔ��Zw  &
�}�B��P��W���]l�;>a�P7�^�x�A����]��^�{�}G�#����;J�Ϊ�w^ܹi�sTH�$�FA��r��y6˱��^�{��.�����W����0�f1�q�����ame��4����ct��_ߪ��g|� ����;  �0=P�'��h}�.mV��QQ��"�B�
����xT��@�	�A��e(H�P~1�}<H|�܍;6���sl�Թ���-jP^���63�|�:���Z7��=_o�(b��v����c�'`��������V1�t��:�TA�����umu��7�ӣ�;�կft  ?�u����     #M�Z5or-	  `p�
9z�b��n�Qm�J[�"�۷��;�l/��}C��!�S���
ǈd��y�}Pb�9q�%u��?�-l�e�>�
���U�.�

���B��eeX]ϰ3Y�������+@�n��mA��n�KtB��w�Y���:j,�_�;D˥����&�w  @FA�  F�''��pw)An\(��%�L�
�z��^�]ּ o[��l�-��t)1���ڶ�U�*��$�eߛM�I����{�#L�OK�
%��;��K�_	�{�js��U���A���UAw1�n;��R� �J��pU]���%��ţ4G'�׷Z�2��  i­�;�w�<��.��    `��6��7
   �,����D��Y�Zڢ�bg�g�;�B�wh^�lW��lhO��ݽ�=�Οݿ����@�(b��a�?��ų�U��c�r,��s�����>�J�B�����V�(�6���|C�,x�ۛ������S�i����M�$�  s �  #�g&�4��V+�=K	��)�(ſ�jW�=bT�(�p�	Rq�)�jW6�+�)�Ͼ��c��)ہvS�b��I�L� b%�=�	����ΕD+C��x"V?�8�}��]lfh��;�����y��{��agG������}�R���R�f[�����p%��=o��N����si�t�~9��� {��;��9:X
�!�    0�l��Tom&T�L  Y��x��?�CͥjVv}���p7-���ll�)Ʋ���Gt���V��B�l<�HR�Y�?�0de���8�+t��
��,�.���q3�p�������+��,�b,��
dpw�� -�c�_�h�>�T��GDG��+w��$   � w  ����}�<b�N��$Ԯ���BC�+P��RњLE*&H����P{2:���40�{�$�ϙMQJ�|Q�)ռ�Ĭ8�w�u���kOؽ���лJ������PO�r�)7���k	WRъ�gv�!wӀ�+\5D�J"Z:�������h���;  �;��q����:    F���u��6�u$  �����/�ݡ��m/�8!�����o�K��b��G��IR؍|D������!�R��b���h�g���rAV�>a�83������{��.�<Ü���<C��s����,KA��b,~�i�y�Z��b�r,a%�F�&}i��Ν���.��&� `� �  C�l[�ե�l�6.��S|?A��
S}��8N7�.����1�n��bwǑ�C���~���Yl`Ⱥp5��J���lSa��YI��b�L��!��,E[C_�]|����֠�����6=�U���������įEA�E��?�.�����\E�  ��|����~m_[[��G�     -VWW���9��gh  ��`��5Y[-Ri��܃B�E���b��,��<Ġ�{X�]�Cdb�����
��B)
��0�m�{QH�{TAVZ>�jlt����~W��� ��	�߀v�=�3�����,����
�?�.�e�Xn��q1�`C�w(	�oVnї�s4vAw  4� �l��}�~qJ�u�'L��Rg\�$F����ıLX�J�R����C�s/@��7,"О��$��a��&�sE8KR�
�o*h���6�/�Un3�j���A%\Q��՝k(^�	W�vwؽ���=�*�mj���f@�]�����;┧�]����n���g�Sm����5�[ ��und��]]E�    `Y3����  `�����e��v��r`���]/�./���,�����2�I>ԎR,s�8GÔ���8A��d�
���M�B=+AG��ߣ{_�������7�r�������лS�%�|�����/��[zk�6=w�h��Yzu�D�U�  �6� ����ǖh�l[<�T�r�z���=H����D�(B�
Q}�f�=\�JW�t�=�8�:O�3.6�l�Ra�~�)h�mZ�2N��%��vw����$\��X�����n�Q���Ղ�/��C�`o�B�,X5i��w�Vw퀻0�#`����;ݨ�)�q��sAw ��byK?��b|     Á�u��V�   ������M�Z���b��>�����C���a�3Tb�<Ĩ�Xq������XL�3Ho�X{��*kY�V����y�6���vUa�n�>��*t�_P���wz��a1V�k�����B�����fe���G4v���e�����
  �� ���](����2m��e�TX[�l)�>q�n�SrA*<�֬����Ѹ�F�=�@{RB� ��������MB��=o��-A+����qQ�v����b�]G�����L�R���;����~�muϻ���"^�P�����b�]lg(�o���wό�Jy�~y�ul���  �K���U�    F�L���n4giw  H1ؾ�ۋ]_PY��hm��kb��bp�ݼ�]+��ON�}Reyuy����3��Q)��K�X��1��V���0긨^a��Ӽ/�+V�]�o��v}��r,y!V�#l�o*=�N�{��|��fw�Pluw���G�Aw  H�  �|�t�ۿD�K�,��UAv�8%�Kĩ>a*X�R�R�!w�O����v�P�y˂���AV�c�̉3/�s��`C|R��(v�4[L�'x������&��A|,_�]%bQ�x%�u+w[z�U�x��:"UG�r�+���ٗntW��VY�]�׷��\���=@�3���z��L��%  �Z#O[��¯8���    ��`�u�ǟ�M0Y  @<���:m-�h�U�v��vo�]]�^���y�q�CYѕ�Ku_r����c=ԎR,���:���H� K��Q<Bռ$|B��$�����m�m���{��>a�z!Q�_���/K�da�v�V�����\��Y:��x��+A���MY�}�hl�<��N��6�4  $�  �A<^�����Ze�j�Bp�]jkj�������(F���U�������(��R&����Qm`�!%)2���e��B���
S:�+N�d�=��%����M���c�"U.@���u�^SC�/��ks���
��l��v[޻��Fw�pp�w����{k��ڢ��}��Q�n��7��	  F������ǯ���~��     �����x��,���  Is����]ܡ�e��X	����(��x�����աv��vm�Ђ����cj�Z�=�0�^-�&��fEYq�I�c��m�QO%��>~�_(����2�0(�.�Uc��ݒ��*��G��W��5��A���[���9;w�^�U��-� �6� @�8{�H_<�IՅi�-�\.�E)� l
����L�*x�{�)aJ&>	U���P��A��m�M���%Zŝ������_��T�9l�S&��ld�#`������9��+�64�
V���������/`��{��v;�O�r�"t�uĪ�L�R��1��:�/ыW�k��9� ���V�N��[�Tp    !���Ưn�Z��	  @B�
9z�R���ߡz�������a���j�P��n\�m��Hw~Rb���}�=Zw�bٛcs~���"q�(�4
�P�|\���0�.)����ð2,=��-Ē����^QV��]��+�W�n��M��d>�t����4�ߢ�.����m5��k  $�  �����g���봱��ry�`��h]�k\(�ۃB�wF*N�UM�J�e!�����(��I�Yx����!aJ���V\1+�U��(a��e$^���)(����V�:��kto�m���U[��os���*���sE�B��'�VW�\�B�]y���~��8�x  Y��p �*    �Q�?�/6���?   �S���K:�5K[K��[,��ؘ�7T4�������C�2,U1�Vȝ���w�h�a�P{Z�XIy��X��%�/��%�����b� +��Xi��g�J ����J�r�}�]�:�_(�{�BwL_��t��7�CW~�d5+3��cT������z7���  �@�  ȁ��p�uy�,'�K�RIj�5-D	�w��6�{*'
N*�*L����a N�>���G9Ԟ��{�96�y�Q#�sd*��=FR�j���{����zawy�O�2��U�}=�*���e{"�(\y���f�^����.���{a_���ͽ�	�_nT��W���4��$  V���"@���     `��V����e4g~w  �I.�K�_*��wis�F�B;��������?���ڃ��@��j�&�X^?д����s���B�&�kc����>�����hz�
��Z��;6ʸ$ʳ��{�a�4jtw�������c�}�p/��4�;�@����ms�	���X���� ��hP~�}��Z(��Wo�[�/�s  �
�  0 Ɗ9�ƥ֝�[����,N��A��_��)�@���֮/L��R�v����~��a��վ0���,d��.�%J�϶8��c[��9_�U��{?A�U�{1����9Ab�L���z�J�����BC���=ls��\K��.�ݫ���'�9���y�ŝ-m`�v �𱺝��f��¯X�_[[�Ç     n*������  `�g��Ra��˫Tw��E*��mm�{��~���ҳ��$�Τ�"ԞU�tl�96�&y����sg� k��c%���vW��x��{.�K�/������r,�ս�6�^������
�
��}y{k�ƫS������Iz�N�   ���;  ��ۺpls��7��r����S��v�h�i^��Q���aJK�j?���)��� C�iVI��3�����9lD}��nf�)N��7�l�IG��.��D��}� �/L��*��\��73��+��R�).C��-G��M���T��b�,��aϭ�Y��x�9:w�~:���^�  �D�i�p��5z�RA�    `Xl]י�����6�  ��O��EZ[Z��R�il���~�|�R�V��.�2.��'C�*�D";�!�#̚?8��Xix{�_�[�e� k�ʱ�'F)�
:v�y��>���zz����W�v��c�W�V����X|�������F�g�Q����2�x���v�>Z@�  L@�  R��%zd��//S��XN0D�
���z�#H	+X)���X��.FyC�Ο��*���!M���ci�c2�tl��q�%}�ax\�
P~L~V��β8%?�U�񠰻)�����U�h�
��,�x%of�	W�x�w����6����h��F�{|�U�šѠFe���D������O7� �n���߿��^�B     `x����w�f�ɮ|  �g�P��tz��Ӵ�,Ҿ}�����=�=D_V��,Ԯ
�{���X���ۃ
�\F�?�9&�q�ؘ���F�(Ϗ���Y.���	Uc�P�/쾫�/'�/��>��:~��/��ʱ�ޡw�f�+�Ӥ�|��S���ͦ�g(��*ϰ�p��k��t��@O\=C�U��&  w  H�����ܩ�-�t�)�u!��u�]���_JP�q����	k^�Ѷ��(��*�qQ�G�cs~���
6~���f�T�y����2�nS�ҝ$^��'����zc���,YK�(Z�3���m���� kgؕ�V��{-�Aw�ͽ����ѽ�t�Y�pj��}W/0
  ���&KF[Zc���h�^�r�D     `8�k�zݬM��&��  
�9�����X�A�9*����b1V�՞������d�C�՞�Y��8�;�d���(��γ}�,?^�*��}.���:�H�˶���Wv�^1�*�����%�9��k���b��ap9֮�G����KZݻ�Y|,�
��0�3l4
T]��O���&/����Suk�_k   Ip ��8�?O_;פ���T[�S�����He#���� ۽-���q!Rk;?	*q�dm���ڇ[��;7���$��ɖ����n�=������DmZ��%�J<O�����D+OP='oi��X�&Y�=�c*�����V��v7���,Ch������xI#C��~���N�����S�z�͠� �a�Z�m;�z}˯�tvb�     �p2w����M،  `B!���^����mj,֩P(z}C��XZ�={V}�y�F�=�=D�kk�Z�=p��X(����,Ȋ~O�'���x��7��vw}@�����G�e�a�׽r,�{�O�b7����cyW�nݛ��Q�F��w�*��/n-ޢ�-�Ɓs��7Z�4  H��  �)�^���}k�[�M*�K�0�J�r/f�E*Y�BP�]���\��%N�!	���T�T�%o�5Q*�@{RBԠ����I�J�{������63�|�16L|��%�*�ٿyK�R9�h����d�Tp�]�����+7��ig�6�Wn��7�p��
�����"=�_�g:G?�]��� �c���~o�H���V��?7��;    �3??o4����y4� �6Ϝ+���}�X^��b��ڮ�[�ի={}�0�0Jk;��u
���C���5�P��1I��;'μ��3l���vq���h� +j�=���F��?n�Y����@����u7��0ms��cy}����+@{��n��^����<C�ݽr��t��w� �͟��nah  ���;  X�+��@c�6�6i�X���1�p��P�6*�S=�J-D�B���s�hI��+L���ݯ��D�#P��-@��v�M�'�R�1}�L�$�)��q�)��6�'�1��T���m
Xz�7���N�{N�����	Y&��NWp��"�.S���x�5}��v�����fw^�p�2K�,R��9z��5v  2�ݪA�}~���     ����5�V�Fs�m�W�  ̃'J���eZ[���b����IWyWz�	���P]�%��ʱ��ʱ�	�nw���Ϣ��q�c�g����:� ��sE��ldE��,�������{L����E���\S{�G�zC�U�U+@˂�U�U�a7̮���momё�5z�����1�xAw  pA�  ,p�x��9�LkKTwĩ1O��/P�.��܋eU�=�u���E�\�8r����$�N:�T���a�C� ���FU�r�0�%J��+J�=lޠ�]�
:&{-�'�hi�U758"��L��W��|~�	���W�6����(\�{o�#ri53���Vw7��y?�{n�}�L���7�!Z ���Z�s��X~���S�N     .�ݻg<�N#  q�@��zf�����R��U�a�K����D�����;4^�|~��3�P�p�z�=k��$��(�
f���(�|��P��'4�T���x^�l���}r�WH��2�0(�������\_н}�ݛ�~a�b,�g��1�����ڬ�����eZ��7�  �  ��`9Ozq��뭋ͼ#N�[ڃ���KJ��`%��u�)�@ej�-L��-D��(X�=��L�ƙccn��</6E)���le�1>�F�$�4�+W�j�X���1ꦆ�h�+okjenhP�ܽA�f�ɽ�iro:��w:"Tgi��p����/��U���w�շ��H��x��V9L�Wt ��z�V[�ᒞ�>;;��;    �2{����*,F  �Q�}�j���7����b%��m�OX����J�0�?���j��U~a��H4�����c�u|�9I�c��K��_��|���b9V�^���_��7Z���x���@�{���;{�;J�p�skR���y��W(~�hhc�.}i�5�����ֹv��e  �P�   ��.�p�H����ؠR�$�dK�D)پn�F�=L���S��vY���s�?�����/F%���*��(��γ}�ax̸�lp�����T��gY�
;�䱰��������
L��$�T*�*H�
oh�od���K��+'��iuw���~�{l�r����'���Uk�����H�.T������m5��5	 0Zpp���m��sss���     ����2U�U�9+�y�6�  ��g��Rn�6*Uʳ78���.�Uav{�a��h����p;���kkO�#���2О��wn�eL��,de�'�g���$�%ƙ#�����$~!u����bI�B��u<��{�Q��9i�]������r�G����ϰ��
�-�L�_�?H����u ��G  0�ON����Z[Z��R�ʝ�1�n�����"U�`�q�]7�N*a*,��&�԰�ړ����:���A�7���y������
Z&b�^����Α헷4���Wъ�_�bqjW��.ޏto73t*W��������~���ze��}j?-�'�i�� ǝZ�����������s     ���;w���`/ ��ġ}����O�v�䴶���y�bs���n!خ�!��/���ů�$�Ο��{��a���y<���a2�tl��Q�$q�,>VZ�(��}^�(Ȋb�;6ʸ$ʳlx�6<�x~����G���x�<������{��A��_�#c9^a�7T�bɼC�R,޷��A��8+@�j�0ͮ�3 �-�@ �&G���O/ԩ6�j�BwIA����*W���{�T�68ОD�=�0�� ��=��{�sm�1g:6����:ϰ>>cC��c�s�<~a*h��*��%-P�O��A�_�\�X�\{�+RyD+�pUp���V��<���7;�UG�������p���t�W�m{{��kS������1�Z�h H��Z�����rA�avvw    �!�?�޽w�x���   *r��+9�/MSm)Gc�����m���a_����c
+>Sp�]ԇ���x���H���1�m�1g:6�s�<�����K�=V�aМ8�⠼°�s��e����D��w�#����������0�нt�z���_X��&�f'����,�������A������S�
=3y�~<M�� �G@�  B(�.l�z9O�o�f�A�r9r�=�y���B�^a�_��lW.%nwft�o����6��2Ԟ�`���8s�8G���~��Ay�Ǐ#L��7�d��MbL����9���{����{W`���|�U<�Jv��3������ �J����/����zhg��|�<�d�Hխ�y] d��+)ݬ���z-�J�677i߾}     ��������&��9Z��  �u��X���YڪlR^����~�Prw�A����w�P��o��u���[�O���ˠ�ä���9&�qQ�ǝ��y���Q�Y���s�U�e+�n3Ȯgc���4���M�}�<>�W�������:�.z��q�*Ў7�ms��݃ݍ��+@�+L�k��r �>� @ O�)҃������z�,yZ�*�J#���������.'(��ۥ���B�,�ޙB$]>О05*�TZ���8ӱQ�ۚ�乒$�H�$&ϟ���gN[�2�E�*�M!Jg�nK�?Ԟ�6���{~���ū�>�=�h��ۼ���{W�j�V����:A��"�ݬܡ����9ze�  =��S7�ί�333���     �67[�m�\_/S�/� �hs�X��=�Jk������<ĠP{��(6���u
��Z+>���!���&�����6�$=6����:gV���F�/�S��Q<B�<�X��M�OL��*�1>��/l����X�~��R�+��*�Ck���?t��V���ݝ�i�ѽ�]���t}{��4�ыWO�k����r�  `TA�  $���/6�6?M[�"���)�t��%���b��`$L��������(�+L���IZ�ګ�U㢎�:'�s�����}�	��|�q�)�s����G��&P��M��A�_|?�2�v$Z�[�h���V�foN^&Z9�M�/���	Vݠ����	�V��<v|s�^�z�^���+� �g�V�Z#G�E�뗙[�hrr�y�     ٤V�9��¿�  {�}E��w�h{�:�V�4&x���P�7+�r��!eXւ��v"��:����_��='α4��1g:6����>�0}q|�0t��!n >J�=�Oh2v^a��$�%�z���^<~�?�������{�g��	ۛ�
�'���7�;+C�aX1V�
���{me�>�_��&/�On���k"  �w  ��K
�ؾC��m*����Z��
T�օ��v����ۉT�Tz��dǙ��2���4�7��>G��X\a*���)��I�v�!^����Gb=�Q�xt�V2�J*Z���f'�����۝��f&gS��{D�B����@��
 �0�
3S-ѣG�Zܷ���޽{t��Y     �dzz�X3Z����~� ��xz�H���hs���K��b,�r,���5�����������̘6��I�?L�#L#�>H1���sl�Թ����5,��=�;�G���T�=-�P6��x������sN�VNr'
�y�����'���]������7��cicI�AO�S�ը��wN�۹��Ɲ: �(��;  t�x�@�?�BkKj��K
bT��������v_�n{�J��la*k�����(c���:'�sd�&�%��|��t�a*j��lއ]�����3�d��Oнs�v×"����OW�R��{E�fG�b�jG*\�awU�]��lk��T���_�=@���{hs $��5���3��M�    2
�}��i�� �'�����p��Ţ�;+��.��>�t�g�p�l������(�'��������o����9&�qq�ę�����ϝ�vn�a�96���qQ=G�s�=����_�<��'�3�.z�;;�^��
;�v{;{��^�W���W�չ��ɶ��D}{�h\��ON��f��bm�  `@� ��)剾~�uA�4M��\�8�h`��˖�S*aJr��d���p��?�`� �����G�ccn��6�>Q��q���sD�l��mއY��3�/39�i���rbC�VKC�P����[��{��7;�j�+Q�jݻf�D���ؤ��=49A/��G˛�  ���,��v����^c���iee��9B      [ܙ�u>�����Vp �r�]z�r�VoSm�A�������՞��MJ��}����s�����1I��Y��8nsL�cm̳5?+�����":ϕ�c����E���f�+;�T��̶_���������n�]r�ݕ��M�B�
�j��=G�K(��f�D+�
*�r�k�s�܁<m��@?��t<T  fp �i��(҃�9ڨT)/��K6�|�T�����ڷ���r�{=��*�qQ�ǝ��y��qu�+B����&�t�4ĩ��Q��Q�����_O��of����0�����w�7�s�}g'/���uG��,A(��ogP	V�h���%Z�8G?��$  �͵�2}�Ħ���7n�g�z�     @v�Ͻ�����fkE�6�  �ΕcE�ܑeZ]�Юo�gU1�y�=x�gY1VP�=�`��g��fq�cIε=�d���8sl�M�\�H���ԏ��͏�-����&x79����U�}��tw���D�Aw�Wt����ao�gO9�b�g�b,Y9V��=.ޠ��x��^;NS�X 0� � ؓ�_�?=�M����-[R0��ݸyA��^��t�T�T�@E�P�T��g����S!V16��4��Y��?�q�c�̱9?��f��?_����cfE����+d�-P�O+��?f{��w�� չ�tW	U����������u�n�{�#`���M-�JK�r� l�-/]��_>N�[9F7� Z �1�V���o�^w��߻w�֫U:x�     �lp��]����L�_v �Qf_���/�+ש��o{�
�P��=ĶW������v�R,�@{r�v�R,��A����8�;&�qQ�ǝg�Y|����ʰ���+�G6�v�]w��8����q��(s��e�)d5hw���{P9V�_���՟���>����h����ʱ6�W顝%���Ezi:G۰ C� �=�W.���-ڬ4�\.K�%!�.��6/t�TS���V�ݽO��~A*���x�L�Fw^��C߇-�I���`�}�8e2vU�q��������L���`Et������ɖl6s]!Klgh��bU�+^��Un�])Z��,Z���c�%z���������k' `��n���TKt�P]k<�f^�~�>��     _�]��2����ѝ� ����E:Ӝ���&�d������r��J����3�{��X:�a�`�^s�K�|�4�øs��dL�c���=?�sQ�(�d�c�3�G��g�+��m{��1I{�6��/�?�[���۞a/��{����O�d5]����궹oVnѷO��͝3��]�� �� �=������-L�N�D山^�=D�
�K����v�0�,0�.�ڥ"?v��Y��$X�8ns�ɸ��α9P�N
��s������{n��T�<�Av�qY������NQ�'t��	U�6��������.���Tb��ʠ�İ;�o,N�__<Bo�=�% V��N݀;3;;K�>H���     ������ϛZ+�Eӕ   ����vn��秩Q*yW|ho�/��-���p{X�]�?�`{V��$C�i��Mƙ��2>�3,�DT�O���h�A�����)��
�Ρ{~�c��#��B�O(�$����w�_�:��7����W}�ns�׷��Tc��v��ϭ2�m�  � �_�\�#�[T]l��ؾ�P�I��^����=�}Ad�m]�X�=������x:�m�1g:6�x[s�<�^����%L��f�=� �\�U��$�(�9&��j�AwjU�	�{����wX��_��	U͐Fw_�]�a�X�'Z	b�����6�����z|�"��u�:4+ @�6
��]�#��x~�q�=���     �����sZ�|铕 ���%:�}�6��`{�/,x�a��'���
�=�|���	���^)��H�P{�`�0�����8�l�9�d���8sl�O������%$��:�~7�����
Î�y,K>�lp�]~Wݩ?���ʱ�<�|~����|�X�����.msWc�x�^8Z���E��-�"  � F����:�-�'�A����Z�����8%�%N!���l�9&�6�ٚ���4Q�([�Tй��G��ƚ�O:c!`%9�fx]��Aw���n#�6~��d�UO�R�34���P�#V����B�����'V��Uo��Wf�g҇[���y�� ���r��pJ/���ܺEW�\A�;    � �w����ϛY/R��'  ���ӟ�ߦ�b�gE1V����՞mc)�C�`�M/p��C�c�u���I��I|?q�>L�o��'jx=h~o�f�]5����iK�/T��k-辻���c�x��'�����������kc����׍z��}B/>x�^���4c �� ���im��Pme�/�^*�7/����@�Rk;��T���ܳl�05�U�uǘ�3g���i�o�򜘊da��D�]5/n�]66�U�qSQ)�����s���"�x,�����KE�]uC�i;�Y�{�O�R53���f���%ݷ77�rs���H�u#O�&^; �\_-�Ƿ�@Q����?���z�     @�8�c�|i��e �Q��ã�ڨ4W|.u���u������b,R��͂�=?�I����f�#̊?��7���hc���o����u����u��Q�ŨAv��$�D[~`ǲ���[�S�C�{�A�X�_h��V|�hs-ƒ��|��4O�*��������  �w ��q�`��rj�����r��Pa�f�v_�}��$���߹7�`�����*X%1.����l�#��e�8B��-Q*�|I�m�u�R����%D��?��;u�
AwͰ�_�R����z��f�fG�
hs���V*�J<.63x� ���Y�Eߝ8H�O�{sX� `F�Ռ>^��<��=��{tee��9B      ]xE���u�y�6���Y   vN�����h�2G�A+>_�����&����!��T��s��ilf�p=�Ax��c���57�s�:�ϕ�5�6?)��d� �°�I�_��o:6�ߚ�C�y
��!���{��Ϣ���V�����g��9^_P��S���=��B�ց�)z�����w�i��6w @�@� 02�r����"\���ݶ8l/4/�	��Ĩ��8�T�°���FU�Jb���8sl�M�Y'��%�Xq����&��l|\!k�*�����kt���t����`�mso
�U���/���Ukk�բ�W��2�����~��	=4y�^���6�  |�R�ǏmQ9�=��G�>�y     ����]�i�Kho ?Nk{�Ֆ��+>b��>����J���Ty�}�����^Ϣh�I��:>�$Α��Q�@��F�1�����A�z�q�@���i��ǒ�U���u���x=D�^g2�H��{�����{�&m���a.��Z��X�����U�����@�,�ʩ��4C @v@� 0L*ЗO���R�i^(�K�p�/�Դ ]RP&P��c���@�+N�.Ȃ�D�Ez2��,	S�"J��l��26����:ϰ<������-aJ5?)q�d�	TA���w�Yн;��B��Q�����n؝H�aX��me��W��@���:�ج��<KJ���}���;g�[��y�V  =�׮��=vt[{���"����ɓ'	     �Í7hkk�x��V�fkho /g�����w��;��*خn���{�^�P�!�����ڳlϚO�5�P��1&�L�Fokn�v�<��d�cD�����mޣx���H�/��h��t��	��P��1��sꕟ�-�'���6��v�{�^�0'������r(�����6�_�;@��& ��A� 0�|�R��nRmu�ۼ���=�
�5/x��~AJ��nE��T�u�tnG!�E,�`���8slηu����fw�r�����l���T�׻m�|+3
y���e�������v~��q��ྦ�X��o�>g�q<�Ƕ_o��ƨ!�$�������� ��(Tⱸ�����W��t��%�w�vQJzw���uA�D�_�r�\�`%�7�FO[�����k�՝�N����Z���v� 0�|�\���ԩ�ӿ���'ND�     ���u�ƍHs�[����  �e���pu��+;��vU1VXV��Ϯ�(��c�o��C�/�"
���٠}&c����۞v,��6�$=��<������������>^T�0hn>�j���3&k^b�~�j�iP=���~���f�]��� ��۾�,���~��3t�c�m�__��.ҫ3(� � C˱�y���Z[�I��.�ۃ�)�8Ծ k^�	TV�)�@E$���.���Y� X�3.�8󢜇C�Z����hyyٹϦ�򶾾N�j����֜muu�9��y���t?��r�����?�9r�y���� ��C������[�>���ǝ1�;v��x��{L]�SA�M��6��q�.P����l���Αl�].d���9�N�-��ngP�Y2�*H��uD+1�rw�)�*q|�r�������q�YA3  �Z#O�����5��^�z�     @�|���/Y���]��� ��!z��R�����+>����
/Qj�c���J��H�?0�/؞�'8J�a�sm�1g:6�sm���A�gdo�7���,�u��X��9~x�Z!�6s��������5�=?>��5�~��{~|���q�x?o&D	Ǉ=�Iy��yI�ޓ
��O�K�9ǆ��/4kt繒����B�~0�Cnr�����{�TM�~��љV����N��'��On���� � @� 0�<{�Dg�����߼�ڮng�I��jkl�
��\�"
n]@�=[��a��-Z���?�q(j~~���t�������h�c�J���b��I�j���l[��|a���k��O�<I<��x�ۣG���Ç�[�?~�Μ9����Iq�)��&��l|\!+m�*��cqC�I��M���wG�L��i-C(��BU�~�p%�r���&��z��5B�+�ڣ 	������5z��J�^�L�s!w @0��9y�N���u�'׮��Ąc�    �d`�lnn.�ܷ+c4X  �i{����X�x�~�н���A�=��:�v�j����
��be1�n��tx=Ip�=�(���3=��������'�X�",��7q�f߳�b,?��s~�,���㍿f=�-�r�𼟏�/Ȟ!�[=�$o�#�g;Ȯ;�tL��z��4��c6�B�s�����=��z�F��{���H����/krov
���
�P,�<CeI�F1o��{���e��;Oo��	  �w �P������˻�Y�F;��q�]-VS�`�\��.h7/P�0.J��T̰�^�j�}����(����>n?���ݻw��u6�x���ܹC�o�v�t��
��ysŹ������Z�b֩S��ĉt��9�k�8 �x��&b�ߓ�L�B�
;�V�]gNRb���t���[�`E�̠
����knmq��2�*ߚ���['���U�e�w�������������Յ#toAw ���f���R�O�"]�5��ߧ�=�     �4[�!�z+
��ݩ  ����<}��6�n�NQ���a�������Cu�����څ-�lwoU���ۓ�	��?�{�$Ǚ��3Gg>kK\ru��}gs��n����~|�o]_���x����0 >_����£� /k�w��~�R,wc?�����<�cϐ=B�UAx� |�P5��WL;��o��%��m��6��݃猪��"4�����c�՟E߰�*���&��V�ů����'/�K�y�n  �� ���S���pq�6kT*��"T_�=��]���Z��
T���ym��T�
���FI�ʒ`e��1&㢎W��d��:��YT���u��u떳���
^�n[|Pc<��r��N ��ٳ��,p�>�d�I�SA�GM�29�t��t��{w�lBU�Gw����+q_�~�h%ib�u6�5���]���V������x����  r>X*��G��l���4�޿O�[�     �.�>��666"���v��B  ��wȅ7*����|Cي�E�+�_�Y�+�7�y�ʍ��~/�~�=Ͱ� �☍�cLƙ��2>l���ݻ����Oq`����
5|�oYO��h~.9υc����~�;}����-�ŕ�����k��aߋ�8>�jl�qA���9�z�6|D��%���&��=J����y���W������W��w����0����=CI1o[�w�;g��[���H� �w @�)找u��^�F��R�@Լ.P�� QJּ`n���i]t�=���A	V6ǘ�3���͛7���&�y}ff�	�Cp-����xs��@�-,lq�������;}������-qJ6�f�=��v����qC�Q�S��}ϥ�����%��D+�k�h%��>��|�$T���s��󸃫����g�'��hmk�  @d��:���=u|�h�{�Gǟ^it     sVVW���t��sE��� �}�;���D;��i�Y�;�uJ��0�d�goQ��K��s�p;�t?��::�2��k�Y�#�nv���qQǫ氷��u��Cd���|;ݺ��¬�����N�7��;� ��/^tJ���;���{͊|O*��+���h�X�}Ĥ���T�;$�� ����r�w�P��W��Eo��)�6�g�����2�p{s��6���K���.5w��� �d�J �4W���ZY�Ri���.	���T�@%���`�b�i^0
��\���S���+�>(a
�U8qE+^��C�lf��߸q�����M�,NT�U{�7�M�����c��}��%�z��s��Z���Ç�E�8�j�iP]gL�*�x�@�Μ8���I&c�	����"U ��'�$Z��uD���{���`���}��<m������4M���hf  x�p�L����`I��`�z���ߧ��z�     @|�s�;��ܚ���JoΏ  d���3]��3��!����o�g�K���W{v��ڃVy�n��߆�˲}�����9&�qAs��daa��9���E�#�}��<��j5�~����_�i���~��𻸱G�-�&�����8�wcl��I��h3�n:?hLп��"�
�Dҍ��������]�Ք����y�g����!~a���ze����Q���1���$  H
� ��O/h��ڨ�hll,P��o�*g�Y�]'ܮ/R�O,J�}���{��='α4��1'��8����wC켱 �K�n�v횳��)��փ>贼s����rn��\$��{*�ɱ(������ݻGq*���]J%T�[�u��^r�+Zy��v7��mm�\gS53�VA�_���Ls��r�2�4��f @��K�U�G_9S3�7{�.�>s�&Z     ��?��)���'�%Z�.  d��w�@���Q�K�COQ��7�~��.[�9�?���7�����]�f�S�o{N�c6��cc,}��}�7d?����Od����/ߡ����G�&¯ytg�71�~��	��{�P56	?��� ��cI��Q����a�t�t���w�+@�eY2�P|W��εD�x>���m�����Xk��da��|�~6��;  p d�c9�օ-Z[�Ky�T�!U�}Ik{Q*N�/+n�݀��(ۓ����"X���E��=���O>��i�d�D� *�o�����¯����裏:��'''��s�P�8Av�q�,PKb�������E+7�޾���$�_+�VA-��}ϵH>��Ag���%���v3�M���������5�V �63�E�[+�ĸ��_k?v�	'     �h,.-���t��[�ϖ�Tp- �.�����gk�V����w���l�n����S�U�j��������q\w��8����m����|�>�d�������$x{�W�}�k#���X\�u����-���$z�Wv���A��QǦ��}/&���]���
�=oP�t���}��7Ty�&�X|�F�N���������U��>  �� �L���"=R�K���n�B�#T�(P�S������rq�+L�8a*P�"��G��+NeM�ʚ05��U�q�a�C�~��#>qC;�����*D(�)�����
��������#/a����#�<�Z������v�=��x,��eHW�Ϻp��Ztw��=\���+]�*L���$����(R����o}���zf�U�^�_ߪ  0o.�o_�R���%�}���駟}�     ���?�����?,�9!w  �"O�.�d�U����CU�=,��kn/����E[�Y�!�z�n���ݒd���m�xix�Y�m�#�8n�f���\J��?��>��g��� -\/�������_��{�СC��9���X�'B���sd�+��19>�~��9�������o{?��o�s$h��5�N�=�7l6��1�0��u|����]7��)�ꌩ.�џ/���s�ν �-p d�\n��������N��cc}��[�`{Ѹ�=8خӺ�#R�n���ĩ���m�������cq�&9���b�@;���y�ZXX�,�����Y\����l�v<x�>��O;"/Y�B[�Z�#,�6��,����e26�}j�ʹG��ΐ�h���xz�n��+J)����J�
Z�����k�������}�Q��	 {���<}�R�G�l͛��Y�����     �x���$
|���J�   kr���y%�kT/��v�g��y�����`{���������C�:x��Q�'��h�x�q��.{�b��-����$ ����Z�O��\��� �r9���,ǲ�T�]g�m�0�Yۧ�7B+@wW��c��e�a{���.��=�X�m�Awɭ�#�-���۹A�&/�O5��  ₀; `��<P�N��Z�"oj�50�7�X�k^nmW�.�ǂD��%�"����)BJ�JS�JC�2�6D����w�	���`T������_���ǯ�.\�'�x�{�1G���,p��TQ���H3�WԲ)h��'j������T�D+U�]&X�m��}�zD��
�����9�hU[��o�>H��N��"� ����2F�i��g��|Ժn=r�;v�     ��K�w�܉4���^����ٔ   S�<����^���"�Je�gh���}�@uV|nߏ��}DF�CtI��`���zV=�$<D����������o�M�����x ����_��Սxc�5��ɓN{��rQ��Ą��5��g�+;��|R~���A��|d�tw���u�A�#7ݐ;_s���*߰���X^��N�*��X|NW�LӋW��/���udS  �@� 0P�9W�s�[T]mP�\V�S%�@���_��_ZP-N��v�p�,��1*q�w�Ɩ85,��A��GE��߈�e9���G�k���Q�j�
A
�Y����̌����K��0�۹��g��Gy�>����ѣG�sl��ecvOJԲ!heI��2/L�ᱲ`�J�
�\�J��]lr��=��h����s9�h��Y�G�=������^f��z������	�Q~�{����/?����     ë5~��G���\��� �,���"=�y�j+M��Ͼ�,c�P����������C4/��R�=K>a��a�s��a��]�yjj��z�-����� �;g����_w6�_[yh.�b����w�B~�pI�+;���8(�P�?��A��ecڷ�/�;�]�Y�7l��e�X�1o�{^����Y�U]Y�/\�;G�ӛwP� �� ��Pl]�}�*���5j�>$pxAG�
j`��ڋ���`q�+T�
T:Bӻ%�>�8eS8ڋ��Q����9��R����hii�  ���#��#.Y��C�T�O>�Y�>���=ֆ�eS��r,��g\1�dl����<��{�p�RT^�tB�m�J\~P��.6��r����U���U}��x��|� -m ��^�v�H7�Kt�`�h�Ӱ���٧�6z]    �k�篷�~�h0�V����  �B�H��+M�X�I��Rh1�?Ю�zC�E��vY�]�;T����]�9K!�a�	m��Q�i�_'p��]��׿���!�����_�_������C��SO=�ln������s��
Îۘk3���8(o0ʾ�1��n�]~��d+@�J��0�����o�X�m�9o��p�t�q���x�ɭ)�����^/R��^  ~p ��ġ=w|���O��O����eb��l`W��t�T��&�_�bT"Uĩ���6�4ħ����b/���o�;�C��.mllh�Z �`��������~���v||�;޶@v<!���m�Qq�'j��q�V�Vw��{��=��+Z��D+���J����{�t�./����Ã��<� ث�v~��ߠ}��U^"�ͥ��I     r����V3[1G�7�����_( d�+ǋ����QY�R���U�X���xޡx_�z�wt�0����3I{��ld�}�tǈ��/d�������۴�� M��
����+�8Áw^������}��s�z��16��6Ι��dlZ�L�������C�O�l�v�5tV�*���M����7�
�B,�/��;�W��k����r�  �� ���D��7o��z����zbTH�=�}A��.n*QJ���j�YV�	��D����~[cm�:'�9M��-/��r����^�J�B �����=������g�q������-P��hיg�����|[�vq��hŻ5��h��T|�F
�J|<qs��p՞���p���`�]�0���>U��_��／�]ٹN�'/�_C�; {���k�����3��s?�v�i���      �壏>r~)0*�WK4[�E �_�T���7h���ry��3������E���;4)ƒ�7��0�Ŗ/8ja�4���q�iyu�7�|�	������!��=��������1\�Łw�	��C��~��I�L�XV�B��Y
��橂��Vd����5��%��ۥXM�o�b��=�0�R��'��	�K��[�
е�}��N�.^�_͠ ��+ @*�r���s�X�F;Ţ|Y���es{�0�me���┩@����Vf�]�:�>�}Y�?�c�㋋������ij��o~��!F0x���������'N8aw��_����w����ε9'�~A+������}��V�k��n�VwY�=��]&\�Ʒ���҃��w!�����w�h%�U|�W�/ܠ''�G3cT��{ {��e��ޠ��Dk~��û�:� =z�     @�۷o��7"ϯ6r���> �AS�}��.m,\�|���cI��cx���v��E����[^�0x���۞��q�eϐWyf����_w<E @z��I�������6{�����f��}�st���@o(	?�Ʊ�}Ĩ~��ؤ�����
Y���	�-,��{\y�{{�[��in����]�P��ʱ�V�n��txm������S�� �� ��9�?O_?�F�J/�.6��,+(�D!���L�T5/�*y�]�xA�ʊ0�Q�D�����v�_��W�ҁ� �v ��������^z��������/~�Nk�X�~�"�nS���?�A�������J��w�6�!��kg�q���N^����b�ΐ�tﷶ��}���]��XD3 {����ӷ��i�dv�˿��ޢ��%��     {���%z���#�竱����N�  `�L*�s����괶����+���l���|D-�0g��s�� |���n��0����4�s9�� �����������˗�r��|�3N9��Ç�ー���IK�G4	�g1�n�C���A���|�S���
���{�a�����A�>��/�$��f���ţ���1�[o  ��;  Q?U��
w���E�1G��5����m]A�ؿ��Z��k^�ol��S�J�b�D�Q� X���fA�������,� 1����?v���t��!�җ�DO?�4=��s411�kK��������N��q�+bV�B��J)X�uʮy��J�r�,�`��.Ch"X���`��A���K�.�/n"��^b��������s�֧$��^^E�C�l
xV    �=
k�|]'����ݫ  �3�Jt�1C�M�(��M��D1-�P,y��'��D����O�1��9lωsL<η�����\�š���M d��{��g��輿�Oȁw.�z���r%��.i����U�����Mƴoy��;�!���6w�TY�9����6w��Ϯ_蹶�byW�z��6w�_ع_[[�Ϗ��쑋��x�  5� �ϯ橸|�;��@�X^P��=P��1aJո��]����)ه��ĩ,�س"LeQ�⥃9���;��+���.  F���������c�=�S���x�`��?�����ZI�mݳj���V�[�h�\��s>�6��҃�K��UO��r��UN4�$M��z���L��N����Q�z���^an�@�/��SǶ�箬����|�Y)%��;    � ����F�z�o�R�,�*e �A���ҷ�Qc��J�U�����a�������ü� �Pk�gwe�;�9/�F�o{N�1�8���Ρv�>��й �����������իN�;�\��V�v���4�B��6�%9�F�"R��ܥmR~gGZ�Em���^�н���]��t�y��a�X������)���K��T���� ���; �:�r��󛴾x���r�eA�ܮ#P� ����(N�"��q�T�
�*H�b��g)Ğ%aj�v��6g�x���B� {�`�+6��O��Ot��ez��睶��~�����f�=��i�)dE���Pq���ݑ�:��ab���� l�if�������y����w����[<Fwװ�  {�?,�љ�:�����B�Bx�]z��'	    `/���~��T�V��c�W�����#  ����g��h����l�lnW�����=C3�PԹt�C&kޡ�y&���?��q���+��o���y��/~AKKK mfff��������������}��_�'N8c���G4	�:��<՘0��G�dw7YA�x^�����=��)��o���,]�Y���s=���c�ze����	z��AZڈ�b `4A� `��
�ľ9�.mP�<������۽K�T��vUk����S�~�	��]�J3؞��d#����:������4==������ ����wy���t��G��;����äh���ߦp5�}��b��˾���Ű�x$�s���*�.�w+Yؽ��J�ۿN����  {��������OߺX�r~�L���m�����    ���no��&����8K�^��O��X	 0��(���;T[�SylL��cu|R�D�C�Ȅ��M��$�؜g�/�Q�۞�?v��z��W�@;{���nm��r n�u�W�~�嗝�����B,.���W�BgϞ�E�P���bV<��-�i߲7�+��[��O�
}��&m�=�p��/��cuW�_�_C�
����3\Y��[�?:Gܯ  � � ��/���i�n}w��T���=\�R�f������SY
�gI�JJ�����z�~���:������ �˽{��?����p��qG�z��gk||�cC��#j��oK��j�]ܗ�hE�%�^��_���;�]a�#^u�)��W�`�����x	^^~�;��m� 0ڬ7��ʽq�����+��u3���>o>��C    0��縷�{Z�����R�n�� �oN�*S�,�P�j���W���ڶw(jZ:�!pg�x|{)�>(�0���͛7�P�3n�  loo�k���l��OO>�$}��_v�|�;.�@��~�j��$�z���]��+��u�܃�����r�^)V�z�BUΪ/�.��s�6��v�.�L���W��c�g @(Z ��Z�yp��+�(W,�>�+Z�c
T��3�*(����/V�Mq*�`{�ι�B�w����g?sD����#� ��~���o��lG�q�ݟ{�9'�>66�KR���?�j�l��m�V<�=�c\QJ%VqSu�iTb����to��*��!/�U��&�6w�`%�V����3��7˴�2w F�{���8FOߌ4��kלא��I    E�p;�qp��*� ҧ\$��KuZ_��z�2�0�?W{�}T���w(���+>��C&-�0+~b��m�;�o?��cz����7���S�%�  q������{��y{�ᇻ��zQ��#*��8b���d���ή^���;����t�A�0�Py��ks�b���������?n���D��� �X�ѷ��h�2O�R��v}��]>0L�R],�m^�^T�ɒ85������8��+J���?����t��]�� ����B����lǎ������hיc;�v���&ъ���w��E�J&V�53�!��@�W��k��EcP��Ks��3��'��2� u�[,ѱr�.����ǟ|�Ρ�    �_�p�}nn.�y��<�:7�����   ��8���V����w�J�t���������۳��I��Ohc����s�����_v6�� ���|���������裏�/��x�:a���B�~[~���$C��8ct���� �~�f�{P�]'��^��"�j�g�5VP����]�ޅ#����4_�/���A� �+ǋ���UW6����*G�*���*�p��8%knW7/�E*&-1*+BԠE�4���n߾�R?�я�
�  M�������ߝ�ĉ�o|���~�i�=��z��Eݟ�p��P��/+��qE)�X�ii �Vv�  ��IDAT�'��A'��煦v�A�����[U�Ly�&�]�7�D� ���6�����t�M��&w~]{�G    `��ro����lno�����i��p;  ]��(��۴Qkt�C�K�:R�](�����a�ޡ��ݽl�=+a����:G�9����*ϯ��
���� ���/~���q؝�P.��ַ�E�ϟw�������uΑ�����h�Cl��Dާ��뷹������ð�{^�N2X���-��o���nЍ����9x� �Up D��tb�&mmR/�..%hԾ���Tr��w,H����$�a��j�v����g�(��o:�> ��g�L��(�{�5���	 �'>|����(��SA��G�����9�P$@Y������d���쓙��{f��_uWwUuUuuwUWu��y���j��!�]}����imm�C=��~3gΔ��g�}6����v�WN�Q��[�1/�V�뎴H���L�J�msM����|�lAw���!w��9N7�7���q8�bbo=Ο7OփR��_�^�W��g�Q��n�h�`ȝB!%�n�݂��������h���B�əs�v6a��Wc��ڮ��Y�!�������;tr;�+���Wnkoo�ڵk��/�7ޠH):�ۑ��w�u>��Haw�N�0Aڧ��r��~a�s8y�ۡv+��#_h�A=��ܕM�F>a�����/Pk˱��R���m��%�b�P�̙����K�H�wBHN�@��u~�5�����d[�]ZAe��,8����H����E*����^���0%�`͚5RS���D@!^D�n�ڵK�.��wߍ�?g�u�v;v�����\ǝ��sB �C��ҳ!v�wY�R�U�&w���rL)L%<�ĵPF;CR�ʧ�!��L��._�E�v��yS�ĎJ�|%�x��A?���W��"���o]L�-^���?�B!����������V��i�®����
��pN=�{��H��9�b�ǳ�bi}B����������[�ͼC�1/y�v������
=__֭['c�������g�7�|SZn��v�x�8��Sq�i����Z��K~�Ѹ�Aw����b{�F�����{:�.y��8�*���"�����1�R��O�_}M����u�k�h��z��͛�U�AD��R�P�"�X��sg������q�r�n&E)�H�mZA�p�^�ݯ���LE����y\�c���l\�&��[���ó�>���BH)!^�6m�$-��v�$^�q��x%ޓ��H���C���0����z$-R����(�ܵM�JqJy-��������u3q��E+����q��Qx�k"�t����r�m ���q���k@~�عS�0�/}�K|^$�B)D��[o��C�|�;+�Qg!�XL���ûn�DeeeF)��G4�[+�Jl7���;tr��ٱo!����ￏիW�g�AWW!�����J�K�妛n��e�/��^(�n��h�ioPw�Wt�C�v�g��^���/YP\�������E	�I�PO�K�+z�2�s�5����}?��WZơ%̔;!#�	!��1.�ϏnA�#��V0ש�vՔ��Tb[B��o^�
TzA�l�T�H�/L���mq�k"T������矗D�>� �R(ū3f��sϕ�$�����[�r�E��g_/R�1;E�|E,���9 y��)������ٚ�E�!�v��z������p����)3��@���dO8����¤���q ~�?�a>��Ϣ"�E/B!�/���#��E;l���	ack%!�X̟�Q���=Iy��J��}D�p{01n��۳�����u���k̎}߿��>��hhh0ܟB���RΊ+���#���B�N�6M��_h4^���H��=C9���˾��K�ŵO,]�������g�cY��f�ֽFS����n��>��F��a�tl9Hϐ�� �?%�ٱ����;�.o�nO/ZqJ-T�R�q�0e2��@_���y��Av/�Zv��9�)�D��$��;{����%K����]j�=��p�9砦�FڞK��h�T�+'�s����O�H����+��63��W_3iŪt;C6a*�%c��hӢ�0g^jb�;!�J}W�C8n|$�sttvJ�����gQ]UB!����ny��w���#�����`�R,N�DEg�w��f+�2��ޢ�Y���C�z�N��>^�c_+��/\�f^x��]�V�!	!�\ؾ}���u�]8�䓥��)��"�w�������R�՞�>�d��XT~a� K.ǒϧ��c"̞��!wq�<�Ae�ݤK�W�n���s���AB��	!��2;�Q=M��3��Z��,�^X��xZA���D)�"�aa�v�Qn�S�"B�+L8p@jj_�l��$����x-ܴi���~��8��3�`�w�q�v+�s��R���;-Z��k�;�IY� %�*E��$V)���T
V�qy�AI�RW��V�\E,�*�ш�G���� ��!�ͦ�J���c�zuww�7��g>�i�7�B!^c���x�������h��5�턐"��pA�0�Z2��u|�|�����:�vm��o�?,�whe�b���<�Xcv�ke��?��ڟ{�9����B��Z�E�L�<Y��>�l̟?_�^�_h4^�n�y�C�z��U��[�
��wU�{� K��jW���69ܞ����^w�p�Px�Շq���x�abfkBHy;!D�/�u񋂶F��T��ve��,ܮ/N�:���I�Ȑ��o^pJ�*���S�g�І���W_}UZ���Dmm-� -�\��(�����i�o�������k�;p7����/�h?��7��9��s���{�߽���駟��c�9F�D���ژo �h܋�U�������z⧾H%#�U�v�f$���V��,m�f�I낕��u/ϝ�'wՠ/�!�o�T�?�G��?�>00��o���=3f� !�B����mۆ��F[��1���j��Oq�ʠя����J���ۥP{.����XZ�0�;4���7��x�}�V���/K�����S����Ŀoq�nyW��ǭ�v����/nݿ[�]~}t���}������wn��)����#�<�G}�{�t3A�3t.��sxe�Kb.��|�6w�����BEA���n���K�����mۉ��&�U�g�;!e	$�jv=mt��Z��4ܮ����3��J�J�0���*�(��ҋx���b�On
X�8W1�W�<xPjk_�r%v�ܩ�_�[	��p�����Ŀq���n��倷S=�[���������bq7����\uu5z{{]�!@	�ެ��ߖ�;�C
�_x�8�裥m��rٷء�\��C�*D�R�k��3"[3�hqO��SXv�*����t+��u|�B��}��i�;Zp�Qx�s"�w�xH�>lh�B��)���:N���������ı��f^B!�D�ܻ�6���Ֆ������Z��	!Ea�� �c\+��=��v=��4�nnϥ��?����&����� ��B�v��F㍍�����-�Ο,qK���N�����n�	�~�n޿|�n����w����׻��>�m|���,]�_��q�H%Y���l��ʘ�=D���XMl�I�vQr����BEA����,(�����%�Ik�B���Z9��E�z.�ނ��+���%�b,B��	!*��&�!�ѝ)P�uY��n���)N)E*��9O+(���Lҭ���܉u���w�b�˩��q����{R���'�p-PJ!�����N��E�p��K��VD'�q/��>�n��.KG��wY��^_�V�Vs�*S���'���7�j"������ ���u鍃���o�]����ݻ����O}��v!�22����;7ڦ]vGEs{-�n'�8�ѓ�8&�/��*bc�=�f�˞�<����2�C=�{��Nzy�l�����,ϫV��o��Q#�-��7��[�L��Э�������oír&���Xܺ��ſy�f~v�o^~�s����wss��>���8餓p��J�wYK����e_/�ڕcv��Ny��u��D�=�#J>���mj�䰻�_6�0�B��n���}a���_���)�oc1!����'B{�o�QC�J��̈́)u�]_�Jl7��ە��l�
j/hF�BP��S�w/W��E���?��c�裏�A!$;�5tÆx뭷0m�4,^�Xju?�ä�N�Q��[,A��qN�V��XZ�)!PI[ �����Vy
B�9�D����"2�L/�P��ʢ	�+aF̉5b�̹X��!wBʍ�+#^?X%�|�U��xk[^[����'1i�DB!���{�b˖-�)��%���բ��vBH�Ҭ F�w`0�s(�H���ci�C=��)���>n�K-�ng����R�],���!��_��^���ӧ����1u�Ti{�~_.�s�n�ѩ�z>��3�
�_�hqG,]�%����_#�Ψ��,����k6��z�a�������~�;_d"����/�ab�F�5�n$NIc򔂚p�R�?z"U���B�L�����Eq�+�����'��چ[ZZ@!�>�k�0�o��6�u�]8묳p�E��c����)F岯ۡ�B�qC�R^%�䰻|;-`Ɂu�Vm�]&S�J�_B��o�5/doeP���!�q=��`�l��!�����=P��$`���BH|��n�\u�Q�K�B!v"�A�l�jk���ߏ��``��1��9g�hk@ ��s
��gx���{��b,m�ݨ���C����8'���W���b�
�K�dB)�.Y���sN>�d|�k_�g?�Yi[�~_.�k̮0|�=�\�C_�����м��ωE��5K.�X��aΩ�����A��	!�@k��/d,P�"U���`%�����b��0��RP-L�7/���d��8��0%��[�⩧��O<a�T��B������+W�s�����p�gH��v�Q�_H�]9�h冈�����!ټ ��}x8-^%�k"�л:�'XAլ _n���U�N\4o:V5�fEHY!��׷T!�c��§�mhlDGg'>u�񨪪!�B��tuu��M�l�1��xy"�B&��Do�^�B��Z�P�?��B�o(�ە�X����R�2��:���
�g�H$��_~�?�8�y��}	!�������O}J���ϖ�3K5���q���]W{���ͱ���/�z���!���ʠ�O�J�6��U�a{=CB��	�|1,�Bo�ެ�
Zm_P��+��f"�6�nl�N5���n�BS2� F1��Z�^}�U)`���S�"���o��&6l؀�K�b��Ÿ��P[[+m/DP*��\��fc^�����ar+���XFSʘG�p�|;�8Y��.\!C�R/}��p��xf�tP�"���ack%�)�>��&���v���8v�����B!�"L����uz_Η��p�`��vB������)]�m�DEEeN��LQ��]��R���!Z��B����u'�)�X�}�ϫV���C�0L!�8lڴIZ��n�/<���1~�xi[���BƼ�!�)沮��^��M�,����{�/�Τ�+���2f~V��H�����r,��U���;�<���̾��	)ap'd�R��_0�=m�����Ys{N��S�M+�c��B�2��70�nwB�rr/��f#!J=��صk!���x�&���I�Z�`.��L�2Eڞ���˾�KvWLѪPQ����Ou�]��'��A1�,65ԢR洃CC���J��o�.Xi���9y��O@Kx���bkG�Ըr¤!�t.��&�U��ۇ;�8T�?B!��KOO6�����n'M�!�k��V!�8ʌ�A�0� z��JcUh�J���?4���v�3>�5�gx�b��X��>�бl���ק���}�B�;��-�܂%K���3�ĥ�^�#�<R�Vo��1'��vx�Ny��!T���^H��b��p"쎄_9�	�y��k/m�=3������ϰ�_�4�u]�����!!�@D��W�t"�ѕnn7jp�&Pi�T���i�]n��(��v�8�Ǵ�� >9%`�y��c���X�l{�1�Q�H�"��.mmm���{���㬳��7���b�B�]����dv�B���x���*!@�1u�=��!v�d�d�]y>=�*-<i���6�w3���~SK�����?�D�^�44��R^l�@w4�/M�E�������x��������̙3A!���ScS�o�nkk��t��#�w��%<B��3)�#�{��B�F��ٌωu���d�]n�6�Q��p���P]�0Ҽ�|���\�����aThѯ�?��;$�� >��8�S�}'�p���KAw'�󚇘�zbL��^!�Q�P��:M�F��2�.�N�T0=��I�azh����[�������G���!z���"�2����h_�P�S:B��@��T��n�Bf{���v]q�`jA����
�{E��ul�Νx��ǥ?�p�BJ���~�\�O=��$\���O��ҶB���Ɗ!d�-Z�+b9�.�zj�,9�nu�A=�JtO�.T��:��<ON���h4�c�0f�,����!���� ��S�/O�Cm�� �x�x����b�1Ǡ��
�B!�m�[��]��z��뛫��!�8�	�C8|`��`�;4��9�7�˱�c������v�{�nc�q����b&Hh���q�FB�.�5���^5kp���c�8�����^�C��1����Ct"o�g�����z��XI�P���2�ҷ�o�K��u|�t94��ar������i��q_��ҁwBFGM���D��^�BrL+J
T�i����a��H���'�&���T��v�� ���� �����[��_���~�iD"B)M��/J��I'���.�H
�k��*�c^�����ldP"�Q�􃪰��\�E)`)+e���P2�:t�ԏ�D�R�+r��߈Sg���;r'�������:���^���hin�ܹsQWW'}>%�B�">kl����;̾���a^�W�����!�s�Tv5����|Ck3>����d�]Y��m�g��v�o���q�5&�w�Ԑd��\������x�������>K!�9�k��M��y�f�J�-��ŋ�2m��X���9y�Ӟ���ɞab�gy���e�p89�s,vGRK7���-��{���z��k:���j����}�8e��Bϐ����!#��MaR�}�T�B���L*�i�D*+�٧��8Ԯ�X����S�8}\>co�������_O��!��>�p��oH_��Wq�gJ� n���R����e�J-V�S�`�P��)��T�)*Aw���>aʗnf�*V%O�^�Tj��us�LC�-τo�7����jp��~�eO��P�uN���ߏc���ĉA!�"���ۇ?�ȑΈ��Aw�_�#�8�9��5mM	/0�V�ܳ��,{����nm7.Ʋ�ڮ�U�a�7�ԟ�ޡ2��-o�M��+~�<��ݍ'�x�<�����`;!��0�5���7�t�q�s�9��׿�ѣG%�^��Ӟ���i=Cm�]l�%���ɰ��Ǭ�]q6U�]Y����Ҟ���R�]�J�DPs���;O��3$�`����is��l�_پ���njOߖ��Z�*-T�C��"�f7�ZPG��
TJaJ�0��b�M^��l���{�n�:
S�R��Aw��p�����K/��+���jW�3�nv'֍�VP���b�[�5Aw����h�ܓ���zPޞ��K73����Ī��1(�Gښ���XY��C)+�}x�@5�	��I��ϐ��7c�[oa�ԩ8���PSSB!��\:::�`{gg�#������*�چB�$��aa����6�[����o(ƅfTh1��7T������=�S���>v�m����>���﵄Bʋ���q���htA�q��Iۜ��<�����5��P9��3���٢��.{���U3?�!��w�IԞar�h[͛�"�����x�	)s��!kSjo�
T��v=�J�r�ũ���B���^w�;�3�ƍ����kײ��BF�=࣏>¯�k�N"�p�B�ڢ�Aw���v㶈e�xc�F�Y�}+�úR�2"q?���5�,2%S�F�c��2���sM.}�{��n
V4U":Đ;!���C��SzQ��o|���8x� �O����<��� �B��A|�m���8p��#���Snn��֎
B��T�����֌
m�]��}�g+�>�cYmmW��V�C�Bz���c�q�1l_�b|�AǾ<F!�;����%K���c����7��ɓ'K����<������(y�g��q��(�cP�"��2ʠ{�3����B<C�7T������s'c��j�3$ī0�NH���/����m/B��a�"d>�`�H%R�����d&P�S����t*��R��<N˫��*	S������BF.MMM�����c�IA�s�=W2ќ�{I�*�����K:�.�Ti�JZK�R�r�	�ʟ|���ޒntW62 }��H%�M�S�U���	�K�K�� .�5���FO��Rn4��ԮZ|iJ�����Z���{�n)�>{�,���I��	!�R����c{}=����H�]3�Ԡ5~C!N3�ʏ�L�D��+nO��z�XٽCm�];볱g�-�n��g~�ȼ�]��Wnޡ���˗cٲehnn!���šC���O<!�b}����.m�b�]9榇X�u�ϗFlO�) ���Y�&��F�a��U�=�{S������ �тf�ó���� C�x:q��!A?�hN=m���4lm�2���4��`��@e���hzA���4)2��9n�On�Q�
�oذ��?֭[��C!�4پ};~������D+'�����cgh��9�����C��^P�v��Aw�p5��F���L��K	U>y0-bA����)D/��!�]�8{J/��G{/C�~����v� ��/~lcpp��سw/�Ν�Y�f!�e�
B!��җ�w����l���A�o�����+�b���~|aL3z�����:���w(���g}�c���skn���ڠ�@ֱ���R��u�|���\��=��n����ւB��E�E�D��q�%���/�)�n��h��Xщu+���3�%���>C�jʱ�H�w�3L��H=������g�pO�D�7�=ԅ3&ⵎ�h	;�B�wBʌ����A��--Pi�̦L�Sr��f�JG���g���� h廏ǭ]����?��;�B1cǎR����>*��?�|���K���}�Z�{���'�ԍ	�J=���F9设�3Z�t�Hn���r��@����RjX��p�<ak��p���!��p��js{%������}Sa�YD���?DCC���~�GH��	!�R�����)�YU���d�}(~Y�n{>� !��Yc�L�D�R>a�A�ݒw���YU��1��j�BM!V�w�?�`�{�N��<(��)t���B!J����t�R�}B�b]v�e�Aw;<�\Ε�>N�����ʞ�hlW�JQ��9�jʱ��X��7Ty�r�^3���3����@__Ż����Iϐ/��;!eĘJΚډpg�Z�ʳ�=%N)��	�Jhϯ�={�=S��~��NAȋ���)�}6oތ%K�`�����}I!�����K��<����
�y�������r�-�ʍ�|.��b����ˈ}���Sr�A�h���O��.߇/pGJ�ʼF�^/*N�neH�����I��cchvv�R~����Z���|b\���G"l����0��1{��esB!��"l��؈}��K�m�D\��~��"��R�Oa�o���b,y�F~az,fן���b,S�P�!3�T�ޡ[��w�\�Z[[�f�e˖I��B�"���`�ʕ�袋p��c���ڕcNy�^����!whf|V!��=CM9,� �<�fN?�g���f���o��3��(>U���3��!�0�NH�0�6�S&����G��]!V���n4��_h�G�Jl�Ƽ�]�%ʋW���zܶm�p�}���g�u�ՈBH����������K�v�Jp�%H�c^������%_�%G�hgPW��(�jdPݡ�g~�1[��Zp�E�T�]�x����/� R�G�*��z�L|D����d(���vk����}�
������A�K["'�D���q�@!�����&��8p��Ҏ������+���R�i�B���Oa���12��Y��c��l�ܮ�e�p1	��}�p�t+��iuV������l_[�b��ntvv�B�t���{�/H-^�W]uƌck��b�=E�B�ꂩL��'ƒ�v�c)=C#����ܳx�)��Z�]���#����Ĩ)��� ����RL��G@_�?մ`�ڞ5�����H��E(m�]+Z���:�V�R�ڭ
Tv
F^��&N��;v��C=$	T��B��>���J��?�y|�[��	'� m+� ee�|'�sc��+�� }$�-�FM�]���ވ�lrԁw_J"S�2h�Q�=��!ZE#�ۉ�)��� �m)Wv��8�s>9~ G������x�ۿ���;�f�����s�͂B!N"��&ާ��+"�WZ�x���lm'���f�pXo#|� B��v�+����`��l�Y����:AwA.ޡ�a�R�
������ᩧ������c�BH!:tH
�?���R1�%�\���*GC�ʱbz�v{���y���I�B�3�Y!�2H�lrO�z��r,�P��v������F1cp*������	q�	)q���o�{t���L�ʵ��,�.S0loO`��䤸eǺS�仏<v��A<��cR�]U�B�S���ذa���/��k�����q�)+�"0��X�v��c�@{b�ئ�����>ԭ�6w��Sb=)V)��uE+�f�J�J��&T�8������r%2�hs����1&��LT]]]x?�l۾3�O���F�!�B���L��с={�J��b�D)�;�k��ǝ!��j!��s�� �5����WhWs{�7L��[(Ʋ��5��x�Z�����R�#�^x�,]�MMM �B줹���r������&.\(]�8��c������g��G�Ɣ�r�]��Jݳa�3L]'����}��P�T�6��g8��'Ϛ�Ww�3$�Mp'��9����vb0K�٭TF�z���p{��y��^�����⒗,yLLu�����.Z�!�"ރ֮]+���;�<��}ƌ�6�)+��+0��Éu;.�c�����p����ԃZ�Ji`-ɓ@ne�АR��6�'���@�'^!y��x��7Q�"d����;kp�aQ?~ �95���/hhl��ѣGcڴi�?_R'�B�s���c߾}سg��pQ�{ooo6W�w��턐�r�\?�3>�cYmnW{��cY�b�c���Xwc1��s�=�{������B!v�{�n�x�X�l���J�y�O�9��>v�ԋ����h�3�:�.��1�=Cy��_��ͼBs�0���|e�\<�T�/�B2a������B��!�����*k��Ԙq�L�2��:-�y
Tv�ӽ���1��#B^+W��ZD{;!����hŊx���)���
�;֒ؤ+d�BB�F�(��]/TВ�ݒG���XZ��1m���he��u��~�ޗʸ�����Oq��ٓ�U͡�9w.�k�`EH93����Q��� >3��k��b������m۶a�I�2e
&O�,}N'�BH�Y'��)��;������Nk%���~#������M�,�C�����;Tb��۵��c���~�_����sz������n�:��oÖ-[l'�RT>��#�p�R���W_�N8A�'����Ct�+ۺݡ����Ҙ}�a:ܮ�'�f���|FAw=�Pڧ�	��;��A)>T�)A�03$M��0�n&R�n�M:B�Yk�=�"\�	�	T�$Hy=�.�5k���;�����A!�xѸ'�V�^����
�-�<�W���i��m�PAKO�I�	)ޞlk�L���[m3L�U�kE��ӂ�<(�82�1*Ɣ�&�>�фs���
V��;�"~��W�)5CR���
��"^K67K�x7n�N��)����*B!�:���hniI��;;]	�E�}x��ۺ*�@!EE����uO��]'�n)�����F�X����>g������������w(<D�	!����o�--g�u���N�%�.��O1<E/e��[L�P�/LݿOn�J��~�ǩ���ޣb<�ڄ��ƪzB�'��p���Z����70��Զ/�E���JY�*��iqJ�	.Y�/��2�)B!���������˗���/�9眓�����v�}
	�[=g!��v݉лr��X��!Mz�L�R�G���׍��>�^��L�*�T����H[Ο7OR�"dDp�7��w�b��>=1��@q��"^S;::��>���'N��	��~��>!�22D[{;�Z[�`�����f[gH
���;!�n_\7�޶}R�]p�cYnn��+ƒ��,����@�ޮ�r���J�;��y�%�~{�}���C$!���}�Y)�r��[��&M�d��S���!�qL1֋Q���&Zܡ�p�Pymh6t�ZP�����,����a�m9˷S�'��0�NH	q����4J��(e RY�������)��*�(7�\�ٽ{7|�A),�FA!�x��%��������xu�5��㎓�e���c�1^Y/D಺�Xb1Y�Q62���Z�J�v��Ku���6ܮ����}�~�ί�˷#�;��@�B�5vW`w8�O����"�����yV,����_#�O��	�e��ц_�!�Bʕ��!tuu���M
�w�o�]�!Zڛ�Cx��=Q�ۄw����Ds���gh�ޮ;۳%�P��=�Y�Sޡ�oX�wX��u���屾�>�\�w�u���A!�x���<��#x�p饗��_�:jjj,���C�3��g���{�"؎<C��'� {��kH��)�к�.=��H����{pѼiX��B���a������ATjHNaJ+RY�ZP�����*U�ݧ�2o�f���d�8���H��M!���l�ڵx��7�x�b\y啘2e�'D+7֋�Ġ�&��#�+����S��<�,ZeG�ϐB�J,CCzb����=��m���ۢm;�p�l�dȝ�Ct�'�>��Qc��?n��Aw�P�5R4�E ^+G���;cǌ�رc1j�(B!�'�]Gg�l��pqfVɆ�����Jb���"n�;�����B,�`{^�a2��K1�a{��o(֡l��*��ipz��;��>��e�=��lojj!�R
������oǪU���o�w�#3@�b7;G�x�z���S�0���ɭ�x���I{��V�t�=��Y�T�]�˔ڟ�;�����.����!e	�B
�wBJ�S���K��CYE����S���օL�*o�J'�nE�*��� �A�h��Y���z+v��B!����<���R;�W��U)�^YY�x���rib�g���xZ��i	E�{2����Ҥ^ =q��(�S_��B��\{jϭZ��*��i���X��84O)?D�}kG���C~�Dk��)�d����Q�0j�h�gm|?�@!�xd���AOw����� �F������Q�C�	!���-�A��`�7̘�9��ڬϙ�a K1�ٌ��|��v�L�ʱ�;,�w(ظq�ܼy��q�B����_���җ����j|򓟔Ƴy}V�)$�nt�z�V�5���3�}}�=C#�0��/��#M����<�wʵp�>,�7��+r'�ap'��|Y��5"J��h`�>�`����˜V�	��+��ħBαm�6����k��Fq�BHY!f#���;�������SO��R])6/d[/�(e�ob,&	S��	�J�"��)e�J�bג:���U�X��*�J�|��a�V��zp79˷3�B�Hc`ȇ�����uc�8f\�Ao4Ɋp�XZ��T�"�.�⭮�BUu���Z��/r�����BH��W�Ed���ߏ޾>�ŗ��O�.�{������a���vB����sD��9~M_a:복p��w���V�enW��3��)��ɰ���|�)�8p ��s�/_��/�B!���[oI_�:묳p�5�uh�=E7B�����������J0�������ˬҧ�~�����X�X�AoX��%��aΜ@��	��~k{���jZA�Ԃ�)��
i_(u��Iqˎ�B�S�>�����?�)�K�BH9"������ӟ���~:���:̙3�v��.��f7C�`�)���u�p|!R�53���LO=�^���
V��2���[��yӰ�! �q����ht���Ǘi��8�L�����&�(�Yg������!������Pb�o�|�VW.�>�Jߠ�UH���a�B�A(�Å�{�h�hm�m�gec�v�g�R,+3>붶k
�|I�F�Z����Q����������$!�Rz�Ϧ+V������*\r�%	�3�h7=E'C�vy��mNz���H{�iIZ|>�b�\��d��g_:]4wV4V!ʐ;!���;!�̹~)ܞ���ۍ2�4�Z�xzA�p{	
TnNn	Z�iᩧ�½�ދ�;w�B)���X�n���
\v�e����Ip�Ǌݼ�m��M�u���)��آ�R�:�9Zt��P����C�]�ʅ޶}��n�7�8� !#�7���UC8z\3k㟉K�5A|V�h�%�B��}~l;T�]���g�	!�A����EOgk�3�!ܮnn�ll������b�5��9ﰜ��Ny�bٰan��6|�� �Bʙ��6�|��x���?��ϫ
�����}��;�^�л]��2�;i�0�ص� �(�p{.�3	+�r'�	p'ă�57��ܱCՠf$R�O/�hoW�TÀ{b���<*P���U�9��}�����͛Q%���/n V4:������s��_��_YY������n���wYXw7����/�[���7p�o^���^��뭛�]6Դ�߅�������o�s�Q�V�C�V��d3C1E)���z�	�im�r=�\z��*��0�}P��>���}XĐ;!$Ns ��Q�a��(�����n�%�BF��}gO��B�@!^�*,�ٍ���W�-��^��p7�吻�Y����*��"C�)�8ҽCyl׮]��?��g�y�_x&�2b�"?��}��v~��`֬Y���͎qc�X�w�=C���Xz���oh�/Ly��s��c��;e�w���#&bծ�3$�Np'�c�3ϏXkSFS��p��@�
��M-�k�B�;xU9	Rv	Z������;���)��O����ߐ�o��n>w��C��u��uĭ�����_{ܺ7����/�/F�߼�Ϳy�z+���{(n�׈�{����o~��Y�����1{��4/����(�z�E�l�I�#�|�F��ɠ�I���he% ���D�R�d�B�D�}�~�BZ&Ta�بx�wB!�x������� �wW`_O�m��R�c��C���0�s�k�Y���C�Y�M}C���^�{q�h���~�����?����ɭ� ���M�߆����ߞ��!����n޿���w��s��r1���.^o�,gr�o^~�+h*#�o���v���R���K/�%�\�����>�c�Z/ďtr_'<C�|��Mg�2���*����Ý��`���Uː;!6;!�̹�ڶ��@����&P��N-��Yim/o�ʫb�v],"���?�	{��Um�
��"�(�틍���p7\:���.~�n�]��w'�n���Y�y��@��ߝ�_�p�k������n����_ĺu�p����+�,X��[�r2_Q�l[�x���&!b�CFm�z(�7�
V�F ��X4�A���! =~B������JL�ƬQQ�3�J?�(%�B�"���}~���t(��a�f\$�+����gd���b�Bʦ��r,#�0[1VF�]tOl�¸K���-�ϫ^�޺��r�-ضm��.�������pص��߭��Þ�Hn������^�(rӻs빋�b����^��x�q+���߼��+�d�#�o>��x\����SO�G?����/J��}f�pb�EY����5�2�|=�Kم�պ���y�;�p��V�EĽ�B�
�	�g�"�ј��	����f�
Zi`�/ 2��S��g��xY�r;�n����؈[o�����kafB!�"�%K��oHm�����Ri^Ю"p�)J�G�-1&72H[��]ĺ��KL9�mf��(e.,)�W�c��'r_|�,���	!*D���? -ۀi5��UŌ�AT���Bq�����A��	aO8��!^�BJ�P���z���+C����À{��Xf�v�w�Y��_)�ם�<�;�C
�U�B!�x���z)�~����.?���B��X)x�V�U���>����%�Վ���X�T�(�n)�	� ��	"d1�n��@��,O-�g���*;�b�O��ŷ}�-[�;���� �B�5�lق뮻N����ZL�<�s��u����d�*-ɂUb�4�`r�Rm3�פ�!��Q61Jo�\X7��ݙf��}��/u"X'��3�rSj�0�:��5����wB!�z���ā� ��F�j'��"�~�lno-0ܮ�j��j1����澡y!V�ޡS^9z���z�����_����fB!��G�X�B*����q�EI�>�������d >�3To��Z�3�B��̛�=r�&������X����R��2'DeW������A�)e!J��M+������/RNPv���書�����B!�#�V�=U43,X�@%�h�y�\������ے{@V���É��m��h��`%o7�ޏ����m/9˷��AI�W�����l�@e �)ՃR�}R� �V��B!��	�����d�]�BH���p�~��[S!�\���`��+�#,c����7t+�N�P=������o�믿B!�X�������W^yE���c�)(�.�y�#�z�Av�mj�0� K`���8��+T��S�d�m_V]4g�7U1�NH0�N���:;�����p{�Ԃ*aJ)Z��T���X�B)Rv�O������׿�U
�`!�B
c�����o~#�V?��1{�lǛr]��(e�o>���<�_B�J�++�E��`�Ijj�*X�#"����Z�\0oVՃB,30��Ξ��*�1L�a��R=�	�C�c �BF:�+`~���P{k���ka���@���EnoI�bn���cۭ��Fޡ/��;���z���p8���_Z���@!���X�n�}�]\z���w�����C�'<A�z!�3�nt;<Ch�ܕ����7L\������ʽ�6�h��9S���C1ݽ!Y`����Ҭ �5"h$PY
��/�n7�Z�����N^�
Y���o��w�!�B�e͚5ذa���*\q��u�SM��{5�^�6��2������lj�$X�MTc�w�e?X�x�Ѷ�8�l<ɐ;!$O"�>��V,25��Tc\��WI-�����8!���oȏ�:#tE�#b�?�b�Bʏt��9=�M��Pr�g3��,��=BS�P�g�`��v1�����:��~�z�t�Mhll!�B
�����s�4#�(�:餓��|���1;����b{�v��9y�����=&�A��3�e���a��=���h�T��>��3��	q�/�aTw�$*�M�zU����������1]a�R���������tHK�,�c�=B!�8�h;3����O�Su�Q7-�^jM�nK��=��_�`���`��~�k4hדc�Vr?O�3xJ���A_|	�@o 5&��C1��Q�/��z�vM�g�?���B����P"����3�O-�h�gԇ�0�_B��@�R.�BO�A�7�z��<��!�h��a���S��a�]�z+�^�av�zgg��c.[��3>B!�m�6)�~����Ø1c<S��]/f��u��3@a��*u�(�Q���h­�pѼi���Rd>7=������4�R��n�ҋ�4ܮ]��)Sz�}�X���X^z�%�r�-ػw/!��<������·��m�����/Gee��"�v�Q��<�l3���	r���Ա|ꛚ�1��PmQ�i݁����S�4	!�0����V[#��*@����z�c�m��g����U�B
g0��4�4k#C�1Ѹ>0_��?�K��uB��I��C��K��k�Ê��!��7�l7���0ܮ��Y`�y�,5�P�ꫯ��#g|&�BF|���G�|���G�җ���KY���^/V��}�0a��y��� m�y��g��:���/�7˶@���OOab_#�`fk�B�2�����J?�S������R�������m�݆g�}�4XE!�gm���_�6w!Z͟?_��	�)ۺ�T�籲My��`S��a&V��V��i~F�v�̹s�\�!��}���sB!�B��n���&�a�����XJѺo�_�%p��+��S�b�g��Z�
�B)MMM��O~��~�����1~���ci��#���~�P��{�1��sG��!//���Z�bѼX^�iW	�
��OLaZt�xMR�@��n0�H�K�=-V��� UB�v/
TN�SbY�z5n��V477�B!�"Z�����K/�D���*GE'���b�RV�ɂUz�A�
�6���,d�~a����۱�F�2���!�B!�B��º�nW5�+�C�ٞs�g܍��f�a"�.}�������_|�E�;ܳg!�R|D��#�<��k��?�!�8�U�*0�z1��J�3�b|Xnp�x�>��Ɏ/�Vk瑯��G*�Be9V�n\0���g�)!V`���"P7>����Č(���)u��3E�@���Xe%ܞ
�g��<��	*ۺhmS
�Y�&34E!������=�܃w�}?���t��ˡ�!����n�Jy_Z�Y�J��vYf(X�o�����s�~C�B!�B�H��y��q��Vh�B�vP^�%ܮ_���!ʺ���v��@��׳����`�ҥx���B!`�޽��/���>�_=&N��I��ʹJ�3��"��T=�P���5���ؖ��=fҊe��,�_�uέ;O7𚎐l0�N��L�ǿU��`t8����^�H�R�ۃ9���1��v�He%��T���*;�|����?��o����B��ٴi���.�/��r隭�����l�[��1����u��^�)��{$�	}M���s���(!�B!�229k���M�R,=�Ь +�p��;4���v��(o(�C��� �~��ޡ@���b��B!�A�W�^���~����NS]#y�#�;��x�����ɞa�i]�"�3����s,��=�0N�}'N;b.^��b,B�`���P�ǉc�1��)����@f�=hw��0����/Rv�Y�zGG��<��� �B�������ߎ�����?�9���<��`��U��N+���1�s?1�O�Q`���O��[(XB!�B!#�/���ѐlOy���(�L۝	��c	2�C��K!�n����)y����B!�E���p����O~�1c�x�#�zl����l�v?�v�3��Vy�:!w��1�M��Ġ�3�~t6��Yuxu=CB�`���]�ǩ���ۯj`40�/�-��@rQ�18n�n�G_~�v��ٍ�mذ����� B!������ޒ�ܯ��:,^�X�heE�Ү{A�2ڷ�m�VYZ��*kX���%�J!ZE"�߅����N��B!�B)|nz�5"Taɞa��K��S�	?0�G1V��v��(�ǯs��J���!!�R���U�V������~�3�x�Ҹ��v���� ��y���@zfA��+����ZL��tn��%�.���i�N��{9�3!z0�N�T���Ξډ��1�`R�2�V0cIݝ�'�ţ�n�C\*'�*�c��0��n�w�}!�BJѦ��?�7n�~�L�:�VQ��w�ڭ��H�R��c�[�@yU�j��R?����H�W������w�!wB!�B!��9~J����t��v�0q;��ݩp�<^.�v/{�����^�u�]x��08H݈B)5�����W^y%��?�555յ�������m�z4�&<�t�=f0�]!w5�׃�XƸt�Dpxd�;�l9Ȑ;!Zp'�fB������쒚��۳TF!��U�p�|�PH��\*;)���-[����MB!���<�6oތ믿��~��*�I�^��U� {�����{��V=25����t��t���M�} k�&�%<B!�B!��'GO
b��.�|~�`���=�GLy�����z�a>�v�~��v�ns�X�uz��BHy �����c�����/~��;.o�P�^�л�����Tz�Z�Pr���Y�f׊�q�pnl�&�BC+C�(a��	��=/�ۏp{k�(�jo׈U����L�=d/�p{�)+��YѺ�d�����B!�������_�_|1����a��ўlb�����ؔ��!X�"���K�,��|n����-����)ڱz�0���#�B!�BHi2�� >�߃��Xf)����u}À�?�y��k~���a4�#�<�;�}}} �BHy�u�V\{�������/�\��s�#�;֋���6������ܕ�+0��2Wl>à{bc�0r?.�c�cOg�!D�wBl�º(z�&��m�!��v�@�h�t�=!J��KZ��/ܮ�Z��p{1D'�)��޽{�����úu�L�O�B)m�P�裏J�K7�p�=�Xך���`W ފ`U�ԃZ�.ٲ�2ȏ5��1����c�=�8oj+��B�z!�B!�R6L�ǿW��`tȴ��7�C�e��_��v'|�R���;w�č7ވ��z�B)?z{{q��cӦM�����ӧ�j���sٷ�<C�}M�r�=���	�+=@Ց
�0�3Ln�D�8a�r�gBdp'�&.��(iۋPEe�H���Su�=�6��?��n��+gE��"Pɷ_y��z�hjj!�BF|����i��ˤk;7��s�׭m^�r")\	V�XJ�J$Ī���CX8;�e�U�K�B!�B!��W�ǉcZ0�Q5��b�����@@�˟Q�e9ܮ�GZ���av��^xA*���� !�B�����k�a۶m�����|Eu���G�]�gh�g����)� 2������}5������	�x��?"��;!6��#��5!2hn�,�&��ͦT�T��S��m_�m̥K����CUU!�2��
�/�}�ᇒhu��{��!��d�Vʂ���k:�} e+��`e(Z%�*e+CO�A\0o�o�1|O!�B!���S��+S:��ݗ�+4�Xf��z,�����b,˾�N�]��nw��#�n���Ӄ;��V�B8!�BFį~�+�������kQ[[k�G�]��gh��U�0>(y�6c�/��_,�1L?~��D�g�����X�{4g&#�	)��N��P#�������4��$R�X��kU>b�����V���!�BF.����G}$M?x�I'���`��U�UM��wu�ݬCA��p{j9�����ƹus�t�$�B!�BJ��χf�!�ѥjnW.b��7(�c��n/�?0�p�֭Rk���Q��!�2�~Ճ>�M�6�n��������J��ݾ��g����
�����[1�2,e�=�����pW'Q��*��>2Ra����?9����T�Qs��􂁌����`6�`��ۋ-P9-H)o�RѺ�?�	��� �B�ڵ?��q�%������4��ӢT.�C�2z�vVv��3�\���к�p%?GE�=��mo��Ś�!B!�B!��X8o=�͉p�N)������>���J��K�`1��B�z�'p�M7���B!җޮ��\w�u��׿��t���	�d7�f��v��)=CO��r7�˖��9�y���ә��� ����z��ȅwB�dƸ ���Ɛ�o:���(�����go`�;ܮ�(�v�����-�c�����?�O>�$!�B����'�����_��f�rE�2ڷ�m�llp"�n$,%��n%��J�2���E)^�~��*�Ww�������}QB!�B!�48�}�{PQQ�[�U�e�g��{�4����#�nw𽥥��z+�z�)B!�����J_~۲e~�ӟb	���v�Av��x�3T�+�%���B��f��,�/Ly������8�nVs�g2Ba���<8�ڏ��6c``H��]!PemoO�SE��U�����^�r�WL'����~�!!�B�X�n���j)�~�i��E�b��!w-�s
����6�~���T��ah^t�i�*D"�݁����e�B!�B�6_��P[#B�
��v�G����,��r�;���+��o��&n��F�޽�B!z<��3���ǯ~�+|�S�*�g脟�g�\�#�n��kו	��jhm�]{\�_��1��g���]��ȃwBr�*�Ws�����%�t*K��z!����Y��R����*�"C4��oVvww�B!�
��Iܿ��o��k���/K!Ȟ�6χ��q�t�=��{RtҊU�N�5�rQ����#���š�S�����B!�B�W��� �:��bU�x��Y�����Y1VΥX�۶�ʱCCCx�Gp�m�a`` �B!f������}|����e�]��{��f�uz���,���u3`��]}ݧ�eQ�<"������!�~��}\�	�O����r'#�	Ɂ�/����<��FPO��k`HTV���{6���v
T��zzz��=�P�vBH�"^c���v�z-> CA����GͨZi���ae~�AFq�x�H���h���G�]��{/�mۆn�ӧO/�(et�B��-X�r����Ě�n�ߖjE+�k<�K?�X3=�B�����{Éc[���$t��B!�B!���	AL�	_0`\���;�bɋ�g����c����ۋ����oGG�T��z�jB!�X����ӟ��Ѐ���7n\^�v�˞��s�_^!�gV��L���tP=��R�d�5~��F�YC��3~�r'#�	Ɂ����ڒnW�܍��u�uE*���I{�R�A��bTV���Ԅ���wظq#!��xݭ��AeUe|��^�+*+��V�ە����4���� B����_�gE�D�����'9,��M۶c��G*5�+_W����2�����M4I��F㷓�`��il@�9�9Ab���!��o���}�{R���'��(��y��=�b����ۭ�U�ǣZ��R������l�F�����W���=��^E!�B!�x���8�b/�P{���vc�PY�����e�0�R�R�;��3��e������ZX	!凔�P̰!f���X��t��\�3���@3jg�w0*�@�L��4kphC��%~[�
�c���I�9b�eBʋU�V��?����㎳��e_;<C��s�wt:�nt�1��b����)g���U>�|��qi�Qc�[�~����0���ȀwB,r�<?z[vJ�G�p{����:��n��2��:�
�C���^x�������B�7a��j��֢�v������&L�~VƷUUWI�fdF��r��xL`��	����"�p{�>~K�S�:�Gs�����c�QuR轿��}}菠��}�۽�=���	K?	!�k�.\����kp�WH׊^�̶�-X���+䞥�A{=�K݂�҂�,N��*�sd܇R�J��ub��*<�!�B!�B��j?Nӌ���~1��K�g�W���٬ˬ�����l��W,˗/��7�,��B��xm�Q��,Œ���vQ��L���m��6_vlo�G��nD�]�`� ��s0����0+"|¾~�,K�?E"�m�	�6"����@�,X�q�V
��ٶR�[E}�S�?R�v3�0t��(^�O�Њg����8)p'�'�b��!-P�U�Z���T�`ZA����z�
&�%��X%�eQ�����s�=X�t���hBH����ѣ1f�Ԍ!�T�֢������ޝmm��ݎ�8�8s.�����:���`�O��=c��q�`{F>�����3��}��Ĩ�@uu��(w�)���8F_o���{z��FO8�t���>��L�Z3:-��%[�lI�|sB�$�����'Ɇc @��l`CH�$˙d�KHv��`ccl�C�-[�uߧ�?�=�]]]=�#�)�ߏ��S]]]����zߧ��BgG�QM�ID|`A�Gy�\17������ډ�@=Ҳd�b�kZ��*־��0��f��^�?1Xe	�u����
7��{�⼅���n�AAAD*��Θ݉ޮ>�Q����)V�)t�,nW��r1_8�����Ʋ���?�0�{�9�z�h�M����'`x`Eӧcڌ�F��B ������Y�	�75cn�<�lp���^�Q��'�E�9ϴA����Nlذ�!���P��Q�0�<��^���]���E���w�%��g�0��Ӄs�s�B]Fu�:� &$p'�(,-���Y*���W)pe���
FPq�1 %���a�^&��
J%3� USS�q���o� ����/S�OCaQah*��:u�1��v�gYu�'ڳ��܉Y���򱺶k�B����]�D��O*W�Tu�n��v�Ƶ�jY(*��T:{�n�8�í�9�ww���ۘ�ԝm��n_�}�+�����z�_�˖-�{�IU7��7&��OGu��=����Y�*�# �@��Víu8���5�� � � � ��������{��#Mf�0�0�
:\�#���<��+���s����&2��k�.�u�]غu+�H�z:E�#M-
�M1{�����MF�q"���s�g�TL������=l����'�:2L�j�H4�~���Ǟ={p�m����*�B�X��Ĝ��>Rΐ����!�tqgm�?C,�0���?{�y��|!��;Z���xi	܉�	�	"�Xlݔgy�<��r�*�pmz8/d�w� �,nw�08���hq{�T~�W[�l�w��]�߿SB��L%��>�N�j�3#�1��m����x��|�#�'��������y���yv]E�#���hi5&��J�� ����'�vĀ���v�~���툡}�q.u�e�mس�Cu��]�]����YZ�M�fL��0�-6�!sy�7��P���)�"��y��˶/���Lض��+U��T�֤�z��}oll�5�\cA�v�ZG�$��D,K�z��܍��A����Z���;X%׳�S�IX��b��jlmAAAA����-�F,��a�#?�qo�M��s{,�X���&`)��1V����)?�'w��?��0�jkkA�]ۘ}���(�65,d��E"9�� v�٤b���0�b�wf���م���Щ�S�DeӦM���G�|��8�Ӓ*d�2��X�%K�I�B�џչ�pNWN�/�G�m�����?���^����-1q!�;Ax��v�Z܆���q/�Reyܹ�=zpJ��Bv98E���.c�o�[�������x�G�����|�L�ʾC��w��f�&�M�Z��=UwC웛���3�iƌ�z���Q�k
Zp�]$�vsŎ�6#xR\Z�lג�;�o��ڝ�P�d��<�v�cWu��B����5��]��"a#v��,s���\vp���cdt��������n��H��R��g�<������d�lh�T>\����[F"���y��nP_��׌{��:1�gY&�"����J�����>��k;28�9�U�9Ȧ�!��>����n
XAAAD���� F[����>�"v����y�9COs,1o����Oq{"���<��>��Sx��ǍXR&c��S*H�)X*Mr�w��G�� '���5�4�2��S,�Qn�#&�#̭�Ә�
s"���0ͶR@g{�v�Iɶٵ���C��	�Fax��9�s�X����=n��L`fY��YOf3��Il�8��,�|�wફ�W^i�W��3�3��,�����I�.�
�����v{9��y���G���k�a�7�^��ʫ�N#��ALLH�N
؏��UC�m�����s�-r�;��r�N��385���P1�࣏>�'�|2%hD���U�%31-,dg���mX�x����%]|c^�t������vE�B�csm�.�R}�I�\�v��_0�7 �ӽ���>y��]��ڎ��Z����o {���t�4��Gttvt������>l������x�	c$�o�%%%)sb�� >�+"wi���o�%|�F�'4����r=�r�����������L��ȝ � � � ��� ��j�)?�0�r�y�0`Or�19�;F|����D�c]��Յ�������;L�Y;������"��`�4��G�K)=���PR63fcFq1��^�%�=t�	�S�PP��3�W-�Iɶ���q��s+�d��u(�7���bn��mm�H�̬�e%�+��y~O0�̙2a��z��� uuu���PTT4n����D���5-��?[b��D��ײ�z,�Y�ݭ�3�#�DAw�PpA�������؜��Ђ^�Fs`�<�S���� U��R��Ǻ�СC���	�P���o�Kf�����Be��{��'���jk��bjM]�ol��k�[d��k�bM/q{�]�5��:�-/�^�i���E�\��ܖ] ��2�G�T��*{�^跌��W�T[�����r��-�hi>�CM�)u '�t��#��ۇ���cٲe	��uY:����͠�5����D�r�E����wk>��n��9��So�������]�AAAAĉ�),6bd8�!f��7t;��e����۳�|����#��eR�L��`�e������;�i�&�`v3f�4�졉�
��P�{o�D�D�a�SS�O3���F��vwv�����	ߓ1"4Ad2����iܛ���(g8�u8E��?�W.r��Et��F��2K�6��4���!��9Mh/���>2�"&$p'��0�R�����:�G^P�`��󲸝�s2Yܞ��۷cÆ���A�	�3��Y������9��Zᠹ��{�\۝�jaA����Ĺ�;�����]۝�v�k�)$�kٕ����+�O܎���k���hn�r.��hj�1-XXc������͇��Ԍ��0�Bg�H'���7���r�-8�3"o�rT��,�V��y��~��Z�^�#�<��W�JX�2+��T!z�����C�=��tM>^�Mw� � � �HyAങm���4ƒ��y(�۝BvQ��-j��S,����[�kN/��n����o��;���� �MaQ��C���3Jf:�������UF�3���C�����H"R���lٲ_��׌�ᩧ����a�e)g���M�s-	����,��T��l�9C!�444�O���o�O�=DL H�Nk��۱���w2�T�۽��5����I�nϧ>�����xTlH�{��b� &3�:�Q%����M�"�`܀K�񤺶Q�]��{��r���%nWu�[^���M�i���������暳̽��ޫ�]&���u<�]-++Ms�b�Y���M��`�7���ALV:::�`ss���+�{�x�=`e<X�kµ���Q$G��y���]8f�pq�Ԧ#���C�`��-�pFu5^�K�^AAAD<a���W����!nF��b�@��m��@0�1V &S,�9�w���3!?mi�������}� 3�X\Z��ٳ03�ʜڳs�A�B�s����a�nAkhb�A�W� �C������W_�/|����3��,�y�t���푞�Q�a��W��K��ς9/׭bĜ!o�O���:qAe>��C���ā��bZ �G��H�%��]5A������r�eׅ�C
�Yܞ� ��?��{��"&%,�T:{6J�f[�(M!�v~�Q�Rܮ��we�jܵ��\ۙ[w�I��n5/��p�R��C�c�O�vCt.��vy;^�|Yܮ��Q9����\�y��]�pIhZ�ب��ى��8x� �����L��9~�a4���k�����IX1����K��]��DsdP�sF
XY'ɕ������X���ű�5�{#Y2AAAD����im�tn�:�s�����3�&pW�b�yC�cw�p"���������������1�	f���-S�ٳȝ�H:�ww��9��`����:�d8�3�;��d���=���ߏo�����O��a�6Ɠ[L���|�ոG<F8�Μ!ˢM�����y+��� �		�	"DaN�+:���Q��#�T�<H%����/A*y�A!h%��?n��v��.n����<�_��W ���f�a��}��2)�)�زf;�k�umR�,h�צ񺶻���������e�T@�ڮ��?��:s�8�ݧ�Eum��O�v�k�k���'vV�<�N���ӧc��%FQOw7��1�{K�!�d�����׿���q��c�ܹ�@��%ӱ!=D�Z���{l��]���|����M;`�Kx����01w6��ˇ��2����&AAAA��ӫ�l݃��W�З�]toL����Y�ܡ������a��!q{�m455a���x��A�v�*-��Yef�pz�G� ����r�lZS����f�55�dlHL6�}�Y�fݺu(--�؜��z�[_���u�6	���f����eR��Fݱ��i���X���"�!�;1�aOX���Co[�Z�*FR�������T��ݿ��ʅ��w7�4e��
DeJ𪹹w�y'��׿� &:�S�P~��tV)��k�
YܮKK�VU�v�[!G�\���Q��a��mJ�E�ф�*!���<�i7��.��Usbvmw��%<�[�ԩXĦeK��{[��1��Cc�~]�u��J���z�~��[oŲe���m�o�x�#��ݸJ�j��*X���z7wY�΍�y�	�@U��d,���!�ݖ�����AAAA��e�A�u�"̎*n�ruX�vٹ=K�ǖ7�l�%���q��"n�G��߱c�!���AL�u���g�)S�bDf��Y6J9���\n9��߈�����C�BbR��k����ظq#�,Y��9C���>{k��%�U|�g�?�3��(n��C3����6��ۆ�-?Ӵ޽X4sv����DfCwb�s~����C��풘ݽ,,l8�ݢ�,O�����\��LM$q{�쑖�ڵ���W�����C��T/Y�9��hjQ�ڈ�k��[X�,�v��.��Hb�q��]�V��M���8\�M!�%׷�E=�]�8��;�������bgE�sAگpG�,s��1��N<h>xuu�ݽ�� ��FCC�����[n��g�9�U�e�,r���D�R��92DO��nl�2^��Bw��*���M���8g^>���3G� � � ����)YX܏=�S�)���{�3��g�6�r	�yC���63!q{�˘(lÆhooALd
�LAY�C�ΦS,��TD�����tک8�Ԅ�����1Qٽ{7���:�p����>��9C��'r�Ж[����q�Q���P��l-�r����:�{c�X�} �eh�;��TH�NLjN��P�oq{80)Pe��;�����p_P�0�^��@9P�Qd���,{��׍�)@EL4rrs1{n���bny��TzE͂��Esmw
�!�U����xK��Z;�k;�`��O�./����-�wtS�,�v�~�H�k�(&W�_���ݵ]�ɵ�т���x���4E_���<TU/M�8��G[�a4�գv�^���� &
�����{��e�]f�c2��#QcY'^"w�9�M��V�ۓ�ً9��)n��y�*<���ۋ4��ƹ5��nAAA١?�O�Չ��G�0E�.`��Àe�������b���y���2"��)'���`�z,���s��_��_08H)�ă��O�6'-[b�~	b2�����U������4��lj=�QgC�HGG�!r��w��K.�ĥ1�w��O��K���s�G6���{k��?ԅ�!,)�����l��3fwㅺ��1�������,�D�@=4/a{�@U �`��K���[�.�g�F�Jp\��VV�څ!Q���(n� 1Q�RT�y��7>���R��[M�\�5$͵])$��!nK�����'�N��brm���
��p8�z���>j�5��?��]ؚR����cum�����\:{�1{��ho���z��p7�6� 2���a<�����;Z���%T��Ht i,������k���<�U���)Xe��%G�p�<������j��G����h�A� � � ��˧�G���a�ۃ1��Y~P�Ypo�k�%���ڕ�X^#?G��SN0��,_��� �<�b"���U6s�S~A>�v�!q;A��:}�1-Y������C���݇��A�3������~|�[�2�s���F����c��?{߿"l�%�c����?u�0�н����)�Kd�Ed($p'&%E�YX3�	Cp�ڃ�80X�����`���^�A��9V�omtq��d�G�ǞN{����SO� 2�¢B#5��ųJ�r[��丶C!n]��]˔}�uy��?V���b|
ۍ?_����G ���~Im� �0.�v�X�k��,�k���横�u�;����j��>i�:�eF�cZu����`_]v�܅�#��D���kmm5ݧO����X���^�ږ-r_����=9X���,h���#ݟ�e�m=h��EΡc�JP9���$r'� � � �h|rA�-���*a{4q{0 ��v>Q�3s�ޣ?˂v�(K�b��+n��l�v?����ꫯ� &y�y�;�a�U2{�k�I� �0w����tdt���ذ����& �_KKn��1�#-�$���XE��,nמ7���/�e�%���=gȄ��������QD�Awb����]ރގ�1�����T�H���,�}AZ��ۅ!ҏo�瓵~2����O&����Ad*�)r�bC�M��Xf
xn�.|����н��pmR��.��ua�HZ.w��!��ro'v�P�]}<��L�k���p=ͪ���Q������%�:ˋta=sU�Q��Wy�uW?U뱾O)���+W����kOcC�|��{k1:J��ǟ��'477���FEEEF�)r�X%���Э�2V��TA+�����n���&v�PY�����S|�e���c�4���]���AAAAx��,�����|a���XcS,o����yC��a���bv�}��.ng# �[�۶mAd2��3o�a�5{���8�
�V�ߧ��ߊ�v�������� �L��:�6`����3�:�j�6������϶���t��v|��ãAv�aiI5v��DfAwb�q�B=--�����Ә���<wY�)@�r_�DA�Ӆ��8���Bܞ� �I[�~=6m���4���	�+��[��Z�'��v��]%��E��>�;�h��p��.�)�s;��Ph\��*�v���X�ǵݽY��{?uE���mW�4Kq�I����5��4g=(]��m��fwGjk��ݵ_�J��>��jj�v?}���E͢E�480���Z|�m���N�K�]s�5��}ɒ%��g�Q~�%#x�G�.���e汓]ܳ�C�����*��'/�Z�T��}���*�ŋ�S0��]'� � � ����� *�F	�an�	�CY��*W��f��M��X��!뵙/t����D2A�>��`�z,fv��"w��D�b^U���>��A��;sV�1�>��nAc�>��v���� 2�͛7�;����.,]�4�9C?m���]Ŀ�=��0���ʣ?k�|a�џ�W�9V�������j#�����X�݈�eh�;��H�NL*>Z���ûMq{����)@�}A��n�?�p�h�vU��{��;w�4>{����-���A)��la�7��ڮ�%nwmZ�����M�D��C!�v���%$W���Mu���]d�]�U����bn�wm/ѥ2�E���͸����4���|]��b��T��#�]l+7?K�/3���>���aǖmhnjAd�~���&6n܈�N:)��u���-r�
j�E��u����B���)�ٞW��ay�J��6|M�UO{έ)�ov� � � � �� pjq�z�=s�^��\��;4��bsn��s��2u�0��t��*����q�w���ĉDf��UL�^Y����<�onI�{Ǧ�����6c�}���QAd
,gx��Wǜ3d��`},��K�.�����o�?[�>k�Gfx��l9�C0Â�<!�
���ϟ�Յ
1Bw"C �;1iX83�i�{�%�������C@p_���GT���C2b	R�%($����X�mݺ��r�m�HxP�9�3���h�)��\�3�\ە��Q��x��C�'[�m�K�k�K��,�v�$��C�����n.-(���+VS{{;�|�;�mGWg'"�imm���_o��]�6�n~�e��ݹ=y��!9�_u��U��������v+`�R�S*j�AAAar~�0zۺ��v��ݕG�	�R�P=�stc�,���*�x�c%#�7���/����Z��ߏ��<D�îs����s�8rA��3���9�nj6���cxx���^�o���K|�l��d�/����{�g���U��6ms,����'�ź�\!�z��p~u>^� Ad$p'&�9Y8*�4Y J�<ە�(�Ђf`�����Q�`U�;0�zn�%m�{���-(�����Ђ �t�}�K�f��f�+*��L4��]����#\��+;�ʞ�v��
1��>;���>(���z���+8廉��&�jA�?�v�v�;��G껣�(_v>�y<� ����}0�������u.������]'Jߥ���˻z7��ǟt"�;��:���w`�@�Joo/֯_o<�q�e�������XJ�<{�;.s^E���M��W�";���(#@e;h��G�{�f�աrz%�;FAAAA���k���r 9��Qs�*��@8wP���X~M�����C4c�v��)��&Q9��l#��D���4�x�	<��#�<A�3�PV>�q{ @"4�HW�o�9e�4r��ۏ��z45��J��=������6r��A��3�I��ݙ/4J�yD�8������N��r����=���tD5���[������������Ĥ`mE?z��L���k�A1Xe/p/�Z0�
Hy��;�ܮ����|JEP��:�c��K/�� E�)�S���T��j��
F3�º�D��b]�Brg�\��^[%�p
�]�AW
�=��Z�v]�w�k;��O/q��OBr��v�L�hS)܆[����.��E��s�\���v}�V�&���/������2���vg����?q%��Q��z�a�Y����}����� ҍ���>�������m��fZ�*m�E�Z��Sts���5� "���*�"i�xpJ
PAz/���"`548����g&(^EAAALbV��{]#=��Jq��;:r������vA����ܡ��$k>�ǫ���z�!<�� �tf괩���6��|a� 2vO0A�1���������Bb�HGX���DSS���jCW��9����D�>g��X*���Q���P��jΛ���rS�.��8	&YY]�XZ� ;SҐHoH�NLx��d���	���� �/q{@b09@ɅAv\��VV����L�.�t	>����z~�ӟ��G��(�S����WV`��j̜Uj��S����n\�a�9�k���n��K�n����#�g�;wS��/C)��ݵ].��)���x���tm� ̏�w��;�k���¾)>����?_׹��O���Oe�5�����v�ל����U6�KJp��?�Ύ��`;>غ�== �t�g�A__n��c8�LX�m�$B�n��o��!W�JzPu�|u�2��O�X���Ἢix~7�� � � ��Ɍ�,,�:��`��J"�H�v{�g��=�1V$�v��nq��SHD�/Q��T��\I��>���7"������
TV/��Ad>��X�t	�Ο�C���{j���"�x����ڊu��aʔ)�y2F2\�Ǜ'�wn�k��̈́EJc,�G���q_�#?��23g�p�a�;/NG#=[�B���h̝��A݈H_(�MLhV�Ά־���AQ�.�\�)G�J�#/�e�|�����@�xF"��J�:��B6� ^� ҉¢B�*+��WA*�x�]��f<*q���) �����ׇ�k�R��
���߮F#��K�g���)X���FT��p	�!��"�ve]��]*�$lw��r��U�N!���x\�UsN%�Uյ¹#tTފ�37��ӵ]:?<��l_��A�i�g��SN��9	���a��7��;�V��W�BOOn��6et�*��r��YƯQ�u����C���#92�a��`�����Lv��.��ҝ�v����gTW�ս�0(AAA1���N?��=]C�e�>+r���k{0<�37�
�D�\��K%h]�Ŝ�#�0���d��Zv��a�_����@�Ƭ9eX�����!�۳1!�RX����}՚��߰u���pS3"����~gc�{�3f�4�7�u��E+r7s�,_h��f=��?��k!	ݝ�A�K*��/�?����}xn7�C�/$p'&,��C#��vPJ�<��f���v��rap
�Š<�qo�ma�q�_�1���u�S�������/� ����[1Ջ�pjz��q�?��nV�!��k�Y7��Nնk]U�L�_��J�,���r�NY�C®�vH墛�&W��ס�U]�{;Ϊ�|Wg����!��?wW=�a����sQ�����z�黠]�� <���Gw�qm�ͅ�	�+�0��2t=�m`��� A��W_}�8�����dt�*��,�m󺠇����<J�`��t�2��w���b��U,XfMB���w�bYi5�Ӱ�AAA�$��ݭ��	c}��d���s�����?�"l�h�%�Y��i2�����x�8p 7�|3�n�
�HX,oμr̫����� br�tGl�61�@��=�ݵC�� �t��^õ�^�{�eee���1���*�mE���l,���������򽬘/G~�-�r�QF���\���zkk���rq'��ÁaN7���� �jxA��/�T��])l�>��%hU� ��r�e�It�*Ձ�X�a����/��2"�L)*D��E���Fn^�Q���k��7����}�����Xׯ���:����06�vsYl���Ϳ�-�>��t�]�U�Nq�s\�U�w�p���q�k8ޮ��j�YO�w|����[y|�z��X쥭U=� ձ�%���*��w�S���vT}�M���?�{҉�W[���mAݞ� �T��o��o�ƍ1w�ܔ��E�!x��d���,|��$w-�������]�y��+8�%rwM�;��l6��,t��	� � � b�qlyC-{|�U9�@ `���GV��,c�5Ų̱��!���D��D2-��ZV[[��n�	�v�A�3fc������Bwg�i�AĤ���:�h�X�
�5b��8t�	�j6o�l��+++Ǖ��[/Y"w�D���2�u0�^.�zޝ3�.��{��{�-��<�V��s���A2�"�����#90��T�/$q{�����~�t���v��=U"�T�bY����peOD*)+��E˖a��2�rݧ`]7+������;છ@�vQ ,���b��sA��(�D�b}I��Aֱ
k�>~���T`k�������w;~��ȵ=r߅�9�>G��R�n�9�]�-U5ա�---x��M���mA��M�6��3VUUU)�'*x5^�
���(q.�.�n���Y�tqĠ�3@��9t��+)X580�O�����|+�FAAA��)����E��=j�P4�
�"vU�p���Ǳ���.��t��ر��744� RI0;��U�Y��fLA�����ü�
cjomÞ������#$4%R����q�5���{�ŢE�&��=тw�����}=wq�yC������_{�gu�P��a�)�/�G��`AZ��ɝH/H�NL8�/��P�n����y��tl��UkR�kxA�{����u�ReZ *��>�[o�o��6"�?6���\�b9�N���c� B��}��Q]�b��B��|sQ�Z���[��^sl��j�����;�:ŅΉsmw���G�;����]W�K�k�]�9��^:��}u�߬6V�vm�}�W��Jq����wն�����8�3p��>�w����|=�� �d��,`�D�K�.��"���'�6:��.�7w��IRq�����΃V^�`P=� u=~��ނ��U�ov� �� L����n�<����t����-|�����=����Q:����!���>�ͻ� � ��?�O+mG_���;������v���+�)�h�%������#1Qr��e���[nAss3"UL),D��X��u� �/l���N>��;�{���m;���	"ٰqX�����ի'��=��]d<"ws���P��,c�M�<F~�9Ax�ew1_(
އ��p��.�X7�d�E�$p'&s��3T?f�q!���C��CR�:��;h�z�Y�-tO|`i,��td�߿�֭�֭[A�&� Ջ�f�"���zֳn`�����f��7�����}���n������rmג��W�5�~&ҵ�YW5����;�ێ�0_�^O�c�x��;���� ��d|7�Bv�>z�]�^�w���ꃺ���C���T�q<��煮/��9��>
{w��;}�(C$���:#`u��wc͚5i%rIa���?��wV�ְ@zP����yQ�.��T~�Vb���nۋ5sb;HAd8L����_�I�+��\{ɩ�^��[~�rҷ=uJ^h�y�Ȱ�{��/���¦]� � &7��9������*�r�jq����1�����ͱ��He~1����o��a��F&�T����-���J��AD�d�dc��%�M��k�N:��H6���V��Nr��&�V�8E�F�s���;߮<�2Ĳs��s��\�"g��=m8�����HH�NL�C��S����sdLjq�-f��T.1{�v�z�=V��OA{�Y�w���7ߌ={�� �Iq�Lí}���)Sh�f�����)6�E��b��B��|���qvm7���S�\ەhH�k���ǎ��졦,soGCl��
��b.~��vU�s��~s��zv5]:���y�]^/��[�v�O"uq��.�=Q��Q��o,\��B���Flz�]�ڹ�,���p�u�)V���K K-r���]l���vq�2DzP��u�I�r�<��+�F4̡a	Lx9<2�ށ!&��9����	A������'.Kq;����C=����"�L-�ų���"��` sgNE:��݇��A�!/'�iS��G��>AaN�������A)o��/��@x�g��=�O�9Cٽ��ˇ{�ʵ����a���Y��#֯_���>D2a���h�R�,-AD<a�s�SG[�!t�W[o��	"Y��������ߎ3�<�̰b�h�e�+󅬢`����s��M�n��,�'��z�4!��o�����0�W}�����r���vu�*�s�g���i��L��S2��~�!n��444� �EɬR,]�e�ч8�Dn>�9����]ۥz��Vs�e��D�������$�b�Lخ��T~u�^<\�]
k��Bl� �%����>v��x���oG�?�vu=W��ǵ]� ƶ7�����8A��r�7�r�q��8?T�tn�rm׌o�e�,a���}��3�s>�WŻ＃�����QD����7��N�+C"E�"�Xi�F���ӭd���]re�T�,��;�;�+X���*.v���a���"����|����՟Ƽ�i����v��?���^~ã�/q������p�E�`IE�Q�x��<�[����{�������5�t����o|uM� �xS������4��휛��	��߂��u;��3QE�9�<~��q�q��4�t�[��k|�	di��O��`���������{� �T��x���9�s{0,j��oc�H��	�`����^��Tc%#/q�K/����CC�02�<؃35K��y�{�$� ҃���8���`嚣�k���ڍ�!�ɡ�����s�!3,�nc,Y�6�
���ݾ���<�w>Qe�e9��^K0�hv�&�H=$p'&ǖ�߲'������#�b^0"v�tj���ܹ���۷�h�w�	ڗ��pn��8n�=�����˵=\S^ٱ~b\���IqmWvJø]��n��v�f	��#���\۝N����w<��=|�|����vݟ�|.H;��|U�u���\�}w(�.�Aq��e��d��������q~���יQ<��uN<�d���&��λ��!X�[�w�qǸ]�p�I]��(�u���T�\ /���W/w��O��U�+COG+�V����{���|�/W:���@��=w}�l\u�q��~���܏�E�����Ū�2Gyy�4<}�e�����g^݄tᴣk��-�ή����<�t�U���'Q{�/����۾��WT"a����ع�0v�o&��=����x�p�'�������G��g���*���ጣq��V��_���W5��	�0a�>�PԊ�^&Bu;�g�$n
�v/��(�l���!�R��X�t�G�;�����^0��### �d���ՋaѲ%���AD��/��QǮ1t�{�b������h�a����/L+��H����m��Y2S$c���.���o�g�Y'��<� �2�/�a�����~/����)���Ǒ��}�����=z���|��k����#���T���|�o������"��]�����������:�ͩ�����y�+�ӥ:�C,+�U�g%��/�Z��k�����v�R}��^�vYoK�Ocpm����x	Wv�[���?q;�z�sm��bu>פ��E��y���4i�]�����:b7���pHW�]�V��H:�cqm�z@zo��E9&��w-�]),,�)�~Ǟp�mق���-z�H(�����l䀳�>;�E���r������ŝ��_m'w�#C@�Ƞ[.�^w�ɝ;2�ߏ��a����L�/�����ϒ�]dѼ�������x���b�s�'��_?��x���q�v�6����kj��͗b�te�̩�9t��?Ǉ�� �.�b��8n�<d2��9x캋q΍���~��D������D�/�u%>s�hh� ?J�O�S�.�ы�#K2��mW���W��w�A��_=���N��Q�}:�[�C������"ve���m��HA{<s����Ƴ�>�x�F�$��.\�Ջ"+�FM#br��k.]b<t���;�lCwW"�0��~��ƽ�E]��o�C�0Q�_���Bwݺ�����W1O��G�/�&p�Ŝax����[3���H)��"0��i����9�vo��� �ۃ.q{��r�da�+P�)l7zQ�H���x�O"�dmٲ��777� s`�Y�KV,Gn^���L���^���ZU"�����z*Q�؀ ��pmw����4Kծ�
'x=�X^(W�5��:��a������[E�K
!�s��um��w�&��u>w�s}򹠉���k?� �U-Z�P����wm��>o]�����q4���+y�k�q'��k�`�����EoO"���l�ڵ%r�$xO,���H.�r���ێ����`���Sl��t�.�la� �rg�{���Ŋ���!��0Q���L
���Y�)n��/֦Z�~�1�>���vά�xq㕸�'I�N�&X����ql���9˫f�o���=�"�Đ�"�t�s�'���*�Ǒs���m_@���u�:~�iB�� &='��F_K��7
yC��}�v�˯{��/�G}�̱&^�/��_��x衇H�N$���%X�r9��+OQ�� "2잣�z*Ta}v��m4�"�8��9L��\�/��Ҵ�{�:��QK���Z
��x<ͱc�F�{��BW[^��7�hID�H��AD��� zZ[� U�����]N�R��L^0��X�ڼy3n��&���8~��
?�=Y��=RE*�Ͽ+�D��l~uj/6��b����PԶb�ctd4J��TXnQ��ha���O"X�����кYf�˷���@ +����/�Gپ:W����*��έ;֮r&?�qe�dl�튦��pe�3ʎ����!5��.��-�V�s��c�}��������h�Q/�_M<��ύ=�=:��uٵ�ѧ�����st��}�L�;~�v���xpB�3��GFGB��/������y|�4i�'�Q�d�R,Z��v~����d&�o�����u�>�,`u�w��\W��H*K����%����Uve��T�1�e^n�^.�V�:��;�n�= ��!�	"��1���s�-�_|����@"w"v�P�?��,.�D�SW�/���?�"1d��=��&r����=�}�H�>�_:O�r	��� ��Q�g�S���ͱ���ͱ<��nc�(�����)z�I�p݋t�/2X<�'��~��1�A��	ۗ�Za�	� 2v/1��Ҙl����C[K+"�{�|��^q����$:��Dn�)r7J�eJwV?��{��a�w1�(�ٲy��7���d�E����~��������Xbv9@���G�J=���s���r�2cx����z��w�~�z��� //񀋾R%|c�3U�r�l���g7@�ھ����;sV)f�)CNnz���)���#�L�<���)L�PiKU4��H˭m۳�ѹ���$J��zh��t*�u]]nm�7�Gt���׹f�?�v������sn0�p�[��k��
:mvN57���w��6]�Q=M1�t��@cc�}�v��Z�>���j��v�w���]�]��<4ڊ7��ѫ�췣��A���<T>x��$�ϡ��Qt�����Σ���a�w���C~~��7ԇ�o>`�\R�[�ީr�a��{����=�������k�g>�q�"zR-N�׼����o�f~sٱc�Qte�B���:U�3�틎b Jpl�
XqW��ĂV�-qzU�TG��Μq�"<~��2J�αD��;� �2mJ���
�h.&"�|�ll�sИ�Đi"�L�s�1'��I�>>}�r<���d�o<A��@�o��fu��+�Q��	V�%n�#B���Ja�%^�"w��-ng�g+Ѣ�L�/2X��?�)~��g<`��M*He<����~:�RU�/�6���a�̙�����?����m���a��;K�~e���;;12<��޾�l?��>22����m�����[�J�N�}������$� �������v�kH�'���s]P�̩ؾ���T��c����x��=]��ݾh�%�ew)o��_�y����/s�f.P�e�%����!�1����;��,(:Fd$�9YX<��р��EG�H��*W��3@�v`H�z<D�j����2��;:��7��8�Ͽ�/50�z�����qO�O�;��=�D͒�X�b�!d��o�8�۰�݀�|Y�`֜2��)zSiX�:�RD��jn�����d]^5_����&D/S�I՟��A̫�p�Ŷ\}���y}���6��n�Kf�:��ɵݵ?R���0*j�؎�x��[��b��ja]�ٵ�%@W}nBف}�Q8m*�M�f�I����Z�Spc�ك%�,Q�Gҹ��y�Br=j������e�<�7��QM�H!l�I.3��֑����ĩ�lۆ���/F�<Y��]��}�@
�����;φd���.��D�>E�&�`2�ijw�`-oG|��#��:�+_�V<@%�1�)�]��P�F"w�HG�Б	��1S)�6/l�"��	�0q��q���3�����g^���A$�L�g����D�υ��>�����{t"���Oĝ_:�tj#"&�� =�m֨��>G}���b�0(�����\�?�v�������;LF~��rK?�����c�!��8H�rWl?S��#�d�w�}�:˙^\l�SJf�J��y�:'/5F1욗�m�z����ܜIy�#,қ��g��HY)2"Sw��H�hJ�_:�,t�Eu�"��p7:B�J�f����բ$j��o]�`#�����+_���l��э�4��Frq�m�r��]����`0���.	�{�[pւ*�~/��ɇ�DF�v� z��M����0����AZ�.� l�����ʅ����XĽ�؞���7�4�흝� �xR�x!��^���|K������̑���w?2�K�m���y�=����-�b��^� ؽ&�r����B�+mǫ��-nW�ý⮺J���7��ۅG�C$��ˌ}�e�U�ե��9=J=��!��~)>_�9C ��z=�}W
୾kR���P�� ��)nW}w�A���!���p}�=X��#��C�m�yM�X�6���^�+W`������ X@��{�5~�>���&$�$���x��}����bpc��/��]X��Eq��R�1����#8v�a��,��h��A���v����c{=��	o&�s�HU�<�������8����;�»���=���s���ƫp�m$r�C0��{��W�},���Us�1ں�l;o��Aר�YR�0�-lW�`��v3�ǅ�$n��>�C���?��?�x�>����	�X��m?�s6U�O�3X��[Lоb�*���Nڶ����x s�O���l۩�>s�RX���))�~*�}xh}��O����;P8�����T{3ޯ��;?��Ҙ���m5���E*���>k��ֱ�'C��x��G��x��ER��׼h�e;����^Bw�C���rѻ�kR:���A{ ���K��acɅ�D�qFuݭ��ӝ�ク�A�1808VQ�����)��+���T{,A�M�6��[o%q;7�w��r>��gb��eVY,�	�u�"x��J[���:8���C+�ϕ���m�I ,�����*�/oRզB��*��+��
�=l�s�@\W��Z�c��OA#�藏�x�]�k����R��q~hb�z����s�}���Ƈ��k������Ֆ.���<���v���n<5i���Sף�	o����x��;�#�(�R t���c�r�Jl۲y���O��91�`����ϸ7fN�vU�Iu *�~���G�"�����1�n�VG�E7w/76��t��ixiWj��$��yY�G��ف��4E�W��۞$�;�dza��}T͜����p��y�F�+V��*�YT>�6�?y9�|�����z���`^�Z�Lႏ�0��~au��r|����y��A�Ω�k�ܙ�{S�ܽ����Ǯ�g���9A����jЈ�@�!l��ޮ���g�F}��da�Cܮ�ٌ�̱�C����x�b�D�ۉ�Mn^.V�Y�yU ��,̞;ǘlw6���/����_�*���K�n��R��~A6�b.�����B�aV �0�\6�R�#����+s��/�����N$�E� r;k�%
�E�����2H���m�AU��^��j�/�x��A�͛7�n@kk+"̚S����iӧ���ݖ�ݿ���e�zItm�b;
�xF��{��XW�)���U�-��]MK�
vَ��\��\m��ޡ�������.w>w-�����j�N9��z����U���p=���-]%Z�<�����{��%$w�]�ﰲ�C��(?��8?T�)
��ڮE�>z���òU+���w���H�S��ą��ٽ�\�T1z$R#`����i���iJ��j�A���ܙ��� �{�H��E71`�xN���_�zA��	^x�EJ�Ι9���3'��A�EL��E��.������������0~ے�>}�e�Ȋ�q�s�?���w�ǖ=�*���u��[d
O����������9�.N�I��1D�w]��n}�D�
ʊ��ԭ��t�#��Y���>h8T}��l��W�7��\�y�P%l�m�gL(q�L<�eq���G$n'�ʔ�)X�r�#q;A�����yg��~�nڌ��D<`"wvo��/9a"w�T��3��3�}��������n��ϑ��9�5�`�5�߇s*���n�Ƀ�6"c�]��+:��^�rk�
R�V��=R� ��u�[�.��T6*��4�2���֭[q��ד������kV��d�U6�]�òXw7#	��6����>"
����Cخ�OO�v�G�J�v(��k���[�n���{�]S�E��.���<����d����Ӫ�j�1���Oa]���＼|�t��X�z�z��x��M����������kצ��B2�=X��r�5�};��,8$�2�`���۴E�b��^�D���2x
�E'!`5s`f����"U|�����5!��#*0��Kw]e�L7�N'e"uL/�3ܵc}��+�?�?����w`����Zw)>zԂ1�ÄΏ]w1θ�1����{�s럊Y�Μ���+R.r���vN�ܙ����uO�����e����m_@y�T16Ψ���	9�Q�-�`��=�s{Б+�D.q�۽G|�f�%��+��I�_2�*q�O~����?Aă��,;j%�V�׺]{@1�a�%�A���P�{/�oي��~�x���7��ϯ�⊄��3I��c,9_��K��9Ckh#ox�a�%�]9C�,<�۲�V-�kud�E$�ù�:�Z�� UPREpa0�� U�%n����rb��0q)n߾};n��F��h�T�X}��q�}�ĸ�×^�*d���&صݵ}�(W)�7�
!���{
x�y��S���S,��K,=�vc[.���?�O���յ=�~T�v�s
1��<R�����������wK���h��~�.���}1�)��Q�x�ßk;;��_O��y�MZO���0�h*�\�)w�	x��~�1V���p�=���g�yfZ���u���M¿��¯Ztw.xw��Eѻ������� Λ�-w�jpp���๽ "�\���x�;"��!w��ڌT����:��پ��f���~m��K1s���X^5��:�]}�|�/�iW�]���q�ݿ��}��b�t���'��L�����-�ണkb^��W6%���[2߼�C��&r>����'�ߨ��Ǐ�ƿ��9��=� �FŴ r;�Q�-a�Os,y�g�e��˿{;�	q�r��H��=��S�����1^�)�ңVb�E�
��w!��,�{���QQ]��;vb���1<D�ネ���/��҄���
ʓ+Z��͈�X�\�c,ކ���'s��˞Wb9\�]Y9��S��S�p��D�D�!�;��.b�ew��\u�*�C��
#�ۣ;0h^����C:Γ|�&ng��MM��&�{�s�ꕡ?�9n�3���) ���%���WJ��rgOm�K+���Gj4�vQ�X�tnõu.V�g�]��s���vR�ڮ��q�\�5Y �X�5�k��ϱ����{�:���Q�X�� ���8]��:�Ee͋�����3�q����	���?���Ac�9��_���-��'?I"��+�$�j1`�_�C�^�*�2_�XY*���!j�WG���8����`A$�>���gb��t�"���J~���xrݥ�W:��:3�����3'�]��>an�/l��p6�˾C�t���ݘ>�	L�~�]����\jY��U�:���8����&r����йq��"��͝x���0kF��u�/�w^i���o�d�g����v��� M �w�	���ߣY�X�ܵ=�)�רϼ�;wY�M�nbF��=��X� ��E�xꩧ���?��ILl�w����8z5r��2� �h�{��+W�z�B�ܶ�>�a�.�X`���c$[�az$�3�6�r	�a�y;�+���e�.c�.�G�xb������씙�x���8� 	܉�gJ���&�cR��vS�΅�{�,n���1��Q0� JO��]�ߵkn��8@	kbl����eK�?��sW@���S�ڮ��U��.�c���(���mE�;��u�rY.��\H�k�����>j�e�rx;Q]�5�W��<����|���õ]�S�Br���N�{��יl�r_�k�k۪��~���z:7�v�mM<n�`hB�xϘ;>.�WaǶ�x�OBwW7"Vp������~�� R���ɞ���Ќ%cv���@�s�A;h�P^NUx
t֢r�Է�ȝ ��g>���Ӆ1�ߘ`���R/ngl�kƙ�����9|dE����M�ó����p�&��X��-]���'�{�104�+����8��cj�9d_}�)����A�'SD����������_�-e�v�{�c|�M��앳g�^oIE)~u�U���P{&_=�Dl�ҧ|�l�͹5:z[;g�l��=�)V�Q�M1��Q���+_(�Ϳ�U�X��K�y����'q;1n��+����)E��#� Lrrs�꘣����mނ�u ����J>��q�|�%�P�з1��8���ce)^���9� r���]vr�r�R���gWO��{�A"����H{ήF[��
z�Da�������gx�D;0D#�L����L�~�uס���D��"k���/(p-�/lO�k�R���{�`����v�8�7�\�\7�MC�?V�*�v�=�������r]���vm7�";��c��O]Ѧ����'�ZW��D�*�v�8[��v�1V��5���_
�����rm�r����޸��������L�]ۭ�T��{Ͷ���X���,��o��7��W�� b����pr�����'��cB��H񜏴��ί��;�DvPR�6mA���Õ!�ҝ.�`�J���<�㧵a�4�R�� ʅ[�G�sᘜ��E��i��3����y���վ�3D���L����Sgg&~�KS[7.�����s��G�����Oo�<>y��1�qř��__x[�!�XHw�{�:��44w��c\3w����+1db"w�;1`���^y�y�� b|,+b�u����5�s�����]��QG}vc��Y��yD�����yղ^x��?��c��d&V����?0KA�)�:'��QZԄ-߄��vD�����z��^p����t��z�)rg�Ǉ������ +�1�S�.�ܭџ�������a�5�V��3`w�("Q���HkN(�FoK�ہAZ���a�{�R��^0]b!��6��ۇ�n��x%�X�1�kN8ť%�S���<�/���F��õ��u�z�׵�-���k�������k�S�<v�sޖ�<�-��}S|��z��{��K�%ӵ�%�������1�]U�e~��:�P�v�?��%lZ)���j��3�r�ǰ�c����M�����X�n���pL�<�(<��X�k�5�"m�[W��T���=R����]܍���+6�vv`m�4�v�H_8�h<���M�HGq;�	|�������&����|�[�����Q2m�����w`�o���?�:84�������ŧNX������;�$l��+ b#]E���.�x������������^����B�{��?��"w�����v.?s��A�r�0�;W�gyC/S,[�p�����G}VO���W��I�y*��/����^���8����)S��أ1��AD|�5��<�l4���w��@?"���q�=����sN���W4�:Y���smAX�ȷ�����2��]��|��34���B�Φ�ZP�>��*� H�N�-�Y(i�/a�5p�/���'�C�HT?>�;���� �X`�,?zj�,v����k����*��"Xq���W)P�M�.�]��1����f���
a���K�.W��EBre]���SW��)�v�I�Tۚ���~�Ӑ�Õby(����{i����.���������/��5g�z��q�qlT}ڒ���Y�ӵ=�-���En�:nN!��������?sHe�}
����_��)����g��+�Z�W^��6� ���ى�o��pfX�bE܂=�h��v��|�}ݓ��<`��BW���̕!,xծ�a��Y�j��KKj���Fx �x3��"?��7����^w�!��^��i�}�~�Y3
���+Gg��ߥ|�E�_�9���#�����ǿ��9�u��׿�S���Ͽ��J$�J��ܙ���?�3�[�Lܾ��@�q���8ƿ����_�W�6n���'��=1�m�y��p�G�� ��sN��[��������b���AK䞌Q���1�<_:��㙻����+$n'���.\��V�]H�B�(ؽLeM5�++���رu��B��oܸ�����'>�+?���x���c3Ɗ$t7G~s��P�=����B�nc�t����nDB��|"m���>�����T��]���],a{��)nD��ہ!�H��g"�[o�;v� A��}�Vc�Ն����ο�o&�z��,zU���F=����\݀-Z�k��O��X-�w�G!(�ۊ�w��ڽ;TN�\~����vI�5+� 
�ݮ����v�}7߹�Ϣ�PO~����ӵ��٫�ݿk����D�&��#�Q��r��9]�=�7�nWQ��nh�����k����O�;m��ֶ�����:��D��r\��/aۖ-��W�����)< �{��[n1��.\�Dw����@�S����,(v�nP�vrgx�ۙ+���]��� U�`��5�<� j���wFDt���_?o�9|w7ο����KQ1۟ӯ!2]�!r�D��o]tJL�v�??�g��·�4�h_��9������ĥ1�[���sNZ�g^�"v�������W�~�������˱���ҏ�� ���19�?��i��.S{����^�������xn����>���������y���A��5s���9��]�����}��>K�X<W��!�W .�.y����7�����o��"��+���Ea����� ����^���*����qp��_�~�z��OW>0]���cTc,�w��	Bw�����\����N��������qpp���KQD��X���Ob��~&��t{A�[�%ƈhc,1�رDA�F�*R�(W����3�3󴙝�{��7��vg�y�;�3�;��g>��/r��Y4����Gk�z��3�m���D�!�;��;(��[}<����]������#M�x��܌+��o��&���AA����&O@�JU��k{x� m�iT�vYt*��U�f��W�;"DU�tEq�{��vS�S'��t`����)��6<��3Ko���.t�6�v(�T��\��퐘k�鬔�&��YyU��ۿL[�m�m�.l]�\_�x�]�FHȵ��ݳ��,��b���l7�!]�w���~�v����E:~ŵ����د�|��P��CǍÐa���/��7���ƍq��c��0`@�N�����䞏7[�҉�M˝Nuq����w��}o�����c�@D�3{<n��r^�n����;-'�ic���S�%�<��Ex��u r� ��~��^@G�9��w�#��_�btt��$�N"��j����{yp��������^<��ۗ����v6��7�y��l��������xnX�+N�Օ���l��H�.%��p R,�ꆶ9�W�woq��	����#���d�۳I �����ۖ1ց@A�\Qa	����� "3�s�c�ƖM�-�{cC#"���V�����=Ǝ�qy*E��ZNl"w��S7���\���C�k���y'w�џ���&�|��>-��V݁H.$p'��>!�7m l1{�����=| ��*���&���T�td�(=Y��]xW_}5�.]
�BiY�0jj��>����G.�X��ڮ�s�k;08m�fS�ڮ��%��,'k]��-�C̵]��H�Y����/���W���_D�����Z�ݐ&)��!L3M��w\���"��W{l�!�w���&����1y����\��,��]����	����sg���I;n��Ǔ���VD4V�Ze%���{uuu���{'��dw��g�����*���IX	.�19qr߻c#����ɑ� �����<��0��W܏�ߙ�o�41�<�J��𒯑�=�a_u���/l�]h�M�?؆�-X����|���<H�DaN�]~�"�Da��{~s:��0,�y�����<��;?����)������'�=+��gcH�*�f�߇杭�{{W?�����v�{{&F}�T�.Y$3��?����џ��;���>#ǎvrbADfa�i����?���>짛ֈ����㷿�-n��&6,�&S�ɾ�����!�]Ï���|��~"w��.�
�ڠ�fȮ�t��}��avM+]Mrd"��Ed̩pz�.47�(..R����RT�;KL����{�	�ˁ���N�"V��9s]�����3π �0pH�%n/.QݱbumG\�k��?v���ѩ��K+ί���?T���	�u����$mw)�e�q"7]��<�S�rrf)T}[��W����M�>��m�D���
R<�45v�g�sm���ziں�+�,~�v�_��4B�X\�����ƦG��͵]Z��S��Ը�ێ�rLr?�^��.�e�sl�~}���V��.���������zp����ҥK�D��{=���C�+a%'��iz��;�`4w/�;��P�M���7�Z:�А 2Eiq!n��]��l�Մ�\z>ٸ��p៟Ƨ[�qŷf#�ɛ��o��1�����?>޸�W����L�~�����O�>:j�U�v���,�8L�~�s��G_>2m�<�������ث¹]fQ����������4s;g7=����Q>������� �Ì�B4�Xg��\$�ci̱��aaH5�*�ܨ�:�������֭�DM[�nM���}�����Љn� ��:�o�cF������[�|sn�m�Բe�\t�E����z�gb��t5�w}�������K�n��lJuC{���X���1u����nv!�	܉�b����$�Nܮs`p���v�J+n�=Q�i�hdCRJ�}y�z�X�d	"]�Ub��I���y���T���n��b,z��]�Mh����µ]GZ]�q{j]�݆Fd�I.ں�Z��<-�B1��kE��Ivmw7��Ov?_e_T�3|lhb����n��˓��������'v�Q���4h��cCwA��k; �d"n7S�F]�׺�?w�˖�uΝ��C�7��sO?�O>��ǲeˬ�����Z˝+Ӊ�L�ٽ��"ww���Vr������%r�Vm\�JrP��p0򷵥'؏���@q��\�\�����c��:��_A��Ҩ�+;��Oִ�'�����̺���3�x�۸mθr!��4�Hmi �<2�<�*�v@q����q�϶�����K���]:� ��P]^��{�[�>y���3�r��B���:�F}֑5�T=߼y3~��`��� �h���4� A�ݰ��w4�lڌ�����͔� �Y�f�%r_�`z��l�fK]�����sK���!<j��߰ȝ5���S74#uC}������l݈ne��s/�DI$�@YC��!�v�C�-h�PEA;�����ݝN>y��u��с!R���Һ뮻�׿��}G�א���e*	*��bHص�PE���zi��S+a�BaE�nǭt���.	���Ʈn]Pn�h��3K�$��݀# ��CX�n9nGB;S�N�{?K����Z�ݐfW��~��V��]�u���c�������.�3"q�X5��u��<������e���Ƶ]]W�7� �y<��د-l�	�v�S�<�?Ye	ݛ��@^�����?L�Ά�tB)�DO�c���c�qc�V�����}���7��NN�D�V��'����L!A%'�t���1��P��e?�H-�(n���۫��܃�.:��v�m��L#��+��B��D�?��c��z�r��Žۿ���p��`1��l�?�����n�%�qh-��t.+A�cf�&4�jci��^�f(�a�<j�Y7곎l�'򼮮���Z�
�;������nn!� :lԍ�_����a�G�� �X�r%.��b�p��֭��N�-uE_c,��uJ[�S��k�����;����Z�%n���k���[[Zp\�}xd�G��@w"+`����w�y��$��^�Ђ��U�A������ rǁ!�.�'���w�	��W�>?e�u7�������hFo��k{�m�|������kgֈ[���Z/���N�̉����e�:���Vl�퐦vm��k���ѵ5�.�C�/	���.W�|���D/L�vm�֋�������F�0v��7+��!��)��=f�� �D+$�C��u�)qm�n#gk:�(�+�p/���uس{7�\�:'�|UUU��l�^��QM�.�;Ye�ݳð���_YܮzP'r;3r	���#����Α�~�&|R�����@�䞧��Iq�ͪM;p���]�>�
zq�So��O�u��v���g7?�K�z=������Z`ۮF�m���v��Ȝq�a�tH�8�~�1��O��BHO��F�ƈ�jD>s��B4�oEqI��v�qo����υ��]��T#�,�9�"b�z��ЀK/�+V� A�Qٽ�5�s�U � :&E��7�R�寿E�X�/o��6���J\s�5�ԩSƅ���S�[ߠ1�Bd����o�g޵ݒOp"w����ꆼ�ݳfx���3L�7�6 A$
	܉����B4�ׅ$���h��"r���u�Ar`�|�ҥ�+���/-���.hƎ��Çjߏյ=�`=�ފ!a�vM:[����sm��wm��Iڎ=Ů��[�tN�,u��v~}LCޞ��r�յ]��1qmwo�5�6е��%��$vg�ܿFH���Ǖ���<�=V���|��Cjd W]��e[7���eC>�	s�X���%ر=wExDb��~*++q��
��Չ��.?G%a��5�]��I,�����E�vM�ud��T�ߖ�V̮iţ�)�@Db�j܋3�\��ߙ�o�4Qy��'�Ꮛ_���l�����Z���|i�(��Ó��b��:q���IY_v�˵���<�
���; �|�{�tٻm�EQG|V!�9V<�CY؞ͣ>G#�u���V̟?˖-AxQXT�1��Ð�Җ$� RKe��8d0���������_�~/�"�N0�<�%��X�)���s����t5C[����n	�պ����]/��lDeY��K�=�Ty&2N�J6 ��]#nW\�ei�A9)�� /�����_Q�9�2�-�� ��{�=\}��طoBG��}-煲N�a�c�#�L���M��ڮ���յҙ�S��.'~�vY��N���r[9N?�v���k���q�֬G������ns>����s����1Y��F�����`�ُ�8��v�����NM�6����k���o��$M3�s
��	m<�ùI!�k;߯rc���v�y��E�~���e������Ժ�%�[n����8餓2��ʤ���ا��KXy9�&�9�s�FU��{[�폃���;6��>C��r�%"1lÅ~m؆k�;���������%���_v7�� ���S��?��u��~~�Q��YG'����p������@pl�f4�<6Ɗ�����{{dZH�%�#=�C/�v�G8�ٱF}�F����7�|3�~�i�=z�Ąi�ѹ�ADn�~#}�����^{�?�
���F�����?�AJF��l�%�"�0�{���0Tc,�����}�5B� ˴����B���]7Z3�---8�_�1� �gFu�w�(..SE>	*G�n'�
݄��P��+Bw;	%%�\�d�w�JG���?��S\xᅨ��AȰc�9/5B��-l,n�,��hPvM��kD�B;,��mՋ��0Uq�:gx��Fl��.x� %v�}��#t��CS
\��vnx40M��Fb���JqM�(���>_Av��fx��vS�8�x"�;���k�C��]=���}�8�Lӣ���M����ekjL���4�6P�p+����\+��ҝ'����,"W�>m���ۇ��L�y��'}۶RҊan��Ȯ]�bڴi�gR��{&7_���M���9NL��ΰ�m��=t��C2�����G�������������>߉�f7�;�F� ��'����jވ�u�L����V�قo��;6m�� �i5�h���%���vχ�s{AD��ݣ>g�Η,���~.A�(*.��q�bȈ�q��� ����i������x�o��~*"*��s�U3��׿��H]&�ꊉcI���b�e�4�3�3_#�k���=,n?�u�(.�RݐՀ�vlƤ~C��f���Cw"�[BC�������$�Tn�AA���������ޮKT%!I�#WE�۶m��_��>�!ӧ?��D�>������ 8?�����+K�P�v��FT�Jm�\�����R��.^=��r����hp����'͵]3��$��.Ϋ���.']���x��έ���F��ڵ���p��#5N�硉=�k��=L�6�����!hc4u}k>s6�����n�/�{]R��n��r>]����������?�^y���	6���_�?��=ztƓK��MhɎ�C:r���eX�����$�=�nPv��������=�`�_;iղ�'֚xl��v#������A0��H��J�9|��˯�(O���}~vڌ�����m�Z�� �M�ʲ�Z6����1��=���uuC}�0�{{�G}Nv�|��O��nA�`B�#�MF��rA����Cѫoo���ױ���	l�g��>g�dS�0�uE[���ٵ��Y�/,������eq�m�řbEj�Q]ܹ��=�_�&���FSK�o�%����<����F�����'�d��B;!%&��\<U��v��&��T*�E�HU�����%}��G ���b��2	����M���GK���DU&��O\N$BUt*�����{��.�vy]ൎ^�=��J�N��Ĕ"�vqY�g�r$ߵ���MH����'���ihb������n�c��#i?T���i��I����*�V�i�Mb���~m�ѵ]����E��~f�6��5�.�6��q�/,,�Ga���x�n����ĒV5559�tJ�o_G�?�IX�N�^Cڂv1iŹ4pN�m'�X]��n_��zÊ�ɑ� �H.e�E "��9n0�z�(.
!�a?��~{�;yr�}����w>��Ͻ� \f�ۋ���(f�X��~�v�n��e�{ �v��%��k��T�ԓ�_:����K���,�F��)*.�������A�Iy��8*���������TK \��0w�\TVVb����f^�.��cYF��g���Y�U+��c��p}P�D����h϶)�麵{���hiiŜ�xtU�獈�@w"cݫM������so�%���۩]NT���;���v_��Ƽ�G:D2*���~X̛7���:����O�6e�ʴ�̵]'�T��d����ku~3�O��P�nq+�gXCTl���4�^+���k��rL�޵=��Aq`�v�ێ�ą��ŋ��vIvm��|�l����x�ͮ����R_[ǆ܆#p���"�,��(�caߐ��X\�}���F2�����~��{Ӛ���ǋ�΅�;s�}[l��4ͱf۽D��gajڨ󙦦/ݱyC���F�z��y?�>^^�b���ͦM���n��&TUU�=�ēM	-�|˝[��uN�;2D��#��B�;a�qqg�!�-���-�!� �e� "{�2������~���־��_��g�O���;q�5b�*� x�(D��uV�Ppo�e)�nX����������9�5�l��������+�w�^O��}0��)V�pݪ5 � 򛰛{���kؾu¦���]v�5��ȑ#�R�Γ�Z��1�S7����j��z!���L��Q���(Ϧ�1�3_/�\ܛ�o���C��gt3;��u$����P��%�Jr�(��]v`pU�DU���˽��a���D#��)�J@�}	����ǳ�>��a����b��C�?��ƵP��V�4��k�j��rm�Ϥ�[��Z�fZ,��i��fDTۢpZ�'��q����������a;�z��Wi�Z��1��%ϵ��A�凧��ڮo#n� Br;ص]8^4}����d�m���9 �p�2�e;�aM�_ &�v��-lcbE�cf�!Æb�#��k�.c�ʕ�ꪫ,����ҬL4Ų�d������pn�Vq;2���&����U�ZN���܌jM,Y� �H�:�� ��`�!��eg�Si*0����7.�>X���{���A.%��z!g�U$	��q�[���fXќ۽��M�k��HG�q�����K����&Z� ��_�;�c�YX���x��w��A0�o�nc1�{���3*f��Z"_���	9c,�nh8}�źaA�^X�&:����{,.�������Z����i�[Y�6�G[a�ց�NJ��0�!7Y�sm��W~�����;0���]~�h�"<��� ��=�0q�TTt�}���sj+
���?�y�6� ���z�`��5��b�J� X�����{	x�������v�^��˵J�����!��4Vד�Hk����"i�]p�v1�3/�sh�Eqm���nv��&����>֔��v�җ�3�/��؅�H'n�쳺����Wq�VH.k^Bri_�ɵ�	)E�����������&��u�X9S��h]
Є;��j��~�C���g�Λo� l�o����o������V�]A�����'w;a���OVX�GΕA�����5����Q=o? � �HU];� ��3aD,��l�����
L�~ӏO����p_�y{5��`1�[@���-�[ߊ�bo�vOq��n�������Y;��4��&�͑���T/��ڙ�}Æ �h�C� �`9={��/��]�;A�O?�W\q�U7���["����YK���	axG����>�uP�O�fh/�]/�k��������Q3tD�]7liه��U �X �;�v���;�P\\�80��0J�цԹ0x����줔����7a�QPA�?�������`��gب�=�P빌�&?Ln�v��+z��"r�5��e`!�03�mլc�iU\�*�U�OMԵ]I{��)n�c������ ^v�T���P����sC3���څ��<vg�;���S>y_0����Wi�{6���p޹��cP���\��(m��b�v�uyz�}�\�q�ǲ�󰦍�/���.��v����h���y��&��)'c�C��Ë-�g�X�x���p��M������X�s���WF�I����	���'��_7Q�2�ޮ��<����Xmt����	� �Օ "���/=��r_�^*��~�U|q�!	�u�o಻�����9�_!�v����ݯf�<��a�X;�cy���bzs,F*�:�%z�g�---�7o�5:A0��	� B�KeW{�|��J|���q�f!r���~�_=.��2���h�'�j�:c,�t56��{�uW3�E=|%��,
�M� �K��y���5�o��
	܉�rx�"4֭��9�ǽ�ׅ� ��B!���/�&�d�v'Q��b'���T6ٔ�Je���>��JR��O_8й��fi90�H�k{���sr3Sjc��T���V�_����R�v�vN��S{
۵Bx9&/�vS�3m��ܼ��y�rm7�MWT�l�\�5면K�k;?_$��������M���=���.�^��|e��ej�U�6
�Fخ�l/Z]���Q/�ר�Muy~}��L)�aÇ�����=�֭Y"�a���7ߌ�}�b֬Y9%fO�?��gw�92�U���a�����JT����M{vcVmw<���AD��Mw��$cj{㑫���Υ�u�
C��W_ŉ�G&�ρ�m��g�i�2��Q\��h	���~#?�$Q{ac,�v���˵C��fMܞ��]2�H���a�X�� ]�`⴩��C� ����6u�X���o��M�� ���z
}���~�m�,���d�Zy�K�1_?T�^�B�z�-~o3�a����m��R3�����Ë�⣂�8��	܉�Q2P[���v9)�9� �P����ON9mb*�$��l����[���+���$��kpđ�QTT��g���#�Dm��H��R#Ƅ���sm�*��
���ڮVUQ�:�-4��5XO������{��n��bqmW�����׳���@\�<�}AZ/����^��8_���}Í]�A�	�vV����;!%۵]����Rn^�z#��<��~�w��q��Z��i#�Y��&���� �'&n�WL�qη��7^}�~�_օ.���$��W_���jv�aJ̞���_L�#wHE�����:���î�+����c�As����-AA�0��'��Bh�O�)�nF���!�a登~u*�L�P?���;�?����A�9a���%%%��ݯ~�{�"w�+�׫n�-j��Q��G2�?���X�h�1pH-�<�:^	� "^z��Y_<��&6|�q��Z�?�r�)Y#f��|-�U!��0v;�n�U3O+����|�P#l����u�����mj���xj� �`�U�6N�5�I��(��B�D�΁�����5�톒��$l�Da���6�}Ē�
����f̝;�V��߰cm��0t���c�ۃ���E �-�Ř�����R[�4l����g��=��i|���W��!l�
�5b{h�Ŗ��(�e����Js��d��r;թ\��@r]��J� ������몾��5�h�Ь��.�ؕ�Hڷ�Ⱦ-�$��G��c53�5r��Ҿ�k; ��S�=�,+�k�܋�Y��6r<��uOӹ���s5'l��n��B폩ӧa���X��Cصs��eϞ=���Kq뭷b��Y�tJv�A�K�#������D�)
܅�F�~P����bz�f<�P� �H��]:�'L����:�H̹��W��n�/n�TZ��.:3�M��u���׮Z����QAxQ۽��ִ_O)5�"��aa�S�7�
�J�0�l0_Cd$Cl�|�&z_�t)~��߁ ���0~�D�� �H�eҌ#ѫ_K�~`��3ƚ?�e�u�Gvx1{���ͧ7�r�u4Y\ݐ��}��H�P7��j�e���Ba�g��}�z��Z�M��&�Cw"-��Tk�����E�CH���%�x'�{Ȃ7�t%���G���KP�X����H���bd
��0t��� �랬嗔�b`� ���a�⛖�Q�?�ٽ-��	��HZO�v��TC��=�h��k*57�D����ؿ�}�[���գ����O���ʳE&�޵׮c�cj�=kk@umwE�{ڗ�a���K����߷�ِe�564�M�W��5=����F��~'>]�Z]��צּ0M���D�s��0;����U���U�3|P�T���X�u�YW�ҲNڮ��ZYe���M\���G+?�ϧ���M��YF����8p� �����J�~���?A�,u�l�|+��mFqQ�FA�?ނ�cžt��[���wV�E�(�;���G��Wb�σE��ߊ� ���%���v�܉y���n@EEE\	�lJh�ۇ�}��;~���]N\y&�"�v{�A�V�����$�l�;{�P�S�k�� � �g�%/��F�ICTD:8lH<tE����vљ����}���p�Ջ�}W��îa'tى憐֭������a�h�ŋ����џ�ڡ"|w��:q{���td����?�F�ۿ�����=�,b�
AD�8����y��W�4�������+��m�݆!C�䬘=�X|�P���B�w�f�ꃦ��]�ٮ!��aj�n<�;1�!����H��D�@�
*���d�ށA�k��n��?I���ʄV�E���]w݅%K� ��d�޽���*SɶL�{2�_;|(ƌ;���'�k;;�*�wCIiI�"4�N�e��rϙ��_� �S����.�T�B;/�mX6��}�7�ك�޽�]ۃ��v���J�]�d�oݏ>5���((�՘���]9������_d���	/L�Ɔ~}tbg��4�bIl__Wg���^]-��S�)��/�bl��#ܚ9��(�����͐c��ئ��������C���؎���L�|�p���6nBE������n�m�{N�nY�2������6Kx����X\��I��`wӰ���}Vs\��KwR4\�;�n5��PVV�����0�e)��04��x��3q��ч8}��*����I�o3v�axoŻx�ɧ�^?����gɍL�ѿ���vg�e�~c���[�+�W\Uȟ.��L�!��;2��aDqd�v�MV(�*�mD���=E������"�:��Ž���[� "�`�֘�Wv.��~x�%%"�L:d ��,Tt���x������Ƅ����k��G��V�ͱ��а�><�s��X�C4�rM�x�,YԮ�*Y�ꅆv�]L��U��m߾���<\"�Xl�|^��Z��,w�	2iX���LpسOo��|����n�d�]u�X��e�k�km��;�2��Lo�L.����2�*̐^&ם��1Xk��'̌���5�F ��ٹ;c۞��z}Scfn�ϥc~��a��V���~߰ߏ�]�`��ڙ�ms�)�477c�ܹ�1ssOTp��Qk�"FDN�j-���Y茱���a�F��,cYm۬�a[[�qs���ȝ���7������xe������H9�*t�T��B,I*>A�&�D����������O&D���O~��SOY�d���2��n�Z~&�=�峡���:��(�E��X����c5TH��G�*����l_n����qS6��N����[�.����X�P!��k�5Br� V'�5�y�27��{Q��l��]#�Ո��mUq���`78�Ķ�J
�#M�־1EVH�*h��l�i�_�|�Y�)��~������w�I2~?Ҭ����\w�v�s3���`��=�]��=���~h����y��^�$���qG�Q�8Ӵ7}�/��|S\\�OT�e���i����#�%;��ISnc���k^�	� ��,��ذ�l�N���-Y9�h�=J;gy�1���w���.&��]���lʄI1�v��B�ؾ^��I��=oǐ	���駟F���q���	�t��y��G��ud��
?
\A;����+g�A3�����ĥƑ��ef״����HA��{{u�OO�x��'�w�0w��M�����/�:�e� ������W��qC�&�σ�]�_��8���B��v*KЩiL�s{s,�^�덱B��]�:���t|�TW;�IW/}$k9LTĜ3W�\�Daۖ�ۛ�23�Eii�e��X#�dj�������f�u*���G�g�^q��Ď��A�X����򙸞�w�v����3��3��m�}��]*Щsfn���3���Ϸ�oMb7t��w��R�<}dr�3S��=����2Qr�g��[6m�[�,�jxe�J���"S���]���X��2�K���u��u�]g-+��l�%��X��#����s~���ڡ�o�Ż�[�Y[{h�nئwp�k�e�{��z�&���AScސ��H),IUޜH��@IX�C�n�!u�*Q�0�'�d���|�Nt���{��L&v��R٭�=];�`Pq{�GS��&� ��풟��<���j�Zi�-�V����}Z�US�S'浻�������eA��>�~==]�u�$6��#�0e���i�5qX�N��%�E������� ��ɭ���&����:�t�{C�F������['nw�<r�r��M �k��e�x�����k|,��&����3&C�a�۵]\VP�vmD�[�ӝF$�ۛѶ��t6��Yj����]�������K��� ���I'���	(��R*�QX������k?x7w�}~�A'iIJ��q:'w>QŦ�ݱ#������@A�\s�QZ\��}iJ�y�����v+^�p�H.G���/9她/n�TZ��.>3aq�_��~{�S��A����;Z	�)Vpq�X7�넺�ew�ڡ�9#���#֚#��_�`^}�U�K�^=1y�4K�NA�O�~�u�X��˨�1�"r��^z	7�|3~�_8f���w�Z��1�>bu;c,�f���G�cq5C�^h_��uB^��F�=� [����	܉�2���cKR�%��$����5Ġ���/Dsqg$C(K�Tӓ���m�p�UW���D~2pH-�O���Im	���v��@�v�8TO0�vA���,G#�׵ݐ���SbJе�#vOq�S�]��ͥ��JJ�cS�·�Sd�$�t��5�a����(Z��h��R��NX]/����@[������~�ˎ�9���.���m"��uN�Y7eWn���gB��M�bM�;8��X>�F�,���pmW�1�x�y���Csޓ��n'�>������d�x��+�"<�ȗO?�C��ǞH�]�D���_=jjj0f̘�K@%�_,��m��g�5��p���>䄕��Ҹ��!A�nZ����'��e;��膃$�!� 8���s��R�S��}Q� w��8��w㳺= "9?a8���i(.JNq�݄2��d#e%EXx��0eTb���ث���� ���[�ƺu(..�4�ҏ�vjwj��zc,�v(�<j��kH�v���&���x�KWmQ~�p�B<��� 򗡇���G��� "�uꄙsfa��w�����O-Z�A���NK��=�����u�.���P�������=�wq���ᑞE���!r�[Bw� k�s(Vn��?���D�8�O!wĞ���U�%IŻ1�ɩ���DU���:�)1��7ʇ9��Y�D�Q�~�>ij5C��,�  ��IDATE�c%���t���m��M�!�k�( ���%����Jۣ��C����DD�o�s�ļv�IrmW���5b{@���ĵ]#:�����.��u>��.�vx�3�?ޟ����	�qe>֥�!]����ݞ�)���daz� ���y�S�lϛ>4�A�gbqm�۸=z�$�1#;�|�̵]�����i��j��1I�t�y	���|�Ï8�z��C�?�];w��/��ك+����z+z��v1{2Z�����ב���V�k'�����i'�L+Q��3��� 9�7�ٍY�Uxv-�EA����q��p��ӧ�^~6N��/�ݴA$���q���'n_�����g����"�`�F��[}"���+����� ���2��%�EL��b�Y������ uCK���b@���^�d��1_�k�̵���n��0�	GNA�� � �l���;~��{��W�ak+��㦛n�D�'NLj�'���xbvtK�1V�=�1_;�k�|��wqgӬ�ad�g�-d�#uD�^��a�uÑ���Q���������H	�@m�s'I��P�T�D����$��\��R`�DO:����J�KP=��� ���z�t��߰��������h-��#ҏ�o�u/�{S��TH�)��2=�k�6��N챴���J(�vm��]�j�H�k��/�����{�csmOf쎰�;f��� �C�I�.�9�gݔ�]+$��3��O�/̔��v��)����;�%'������,S�G�G���q��/�v�D]������v~"yq����o�~��O~�G��0>��#��ڵk��1���Z����U̞H߱����s�{�g{��9	+{>Y�n�������`��d���ɨ��)$�G)Qe%��l@U��knAA�l�~��M��[�2L?�6�<#j�-��s�=��-�AD|�2}4n���(%���~Z��pÃ/��0���f1�����g��v����@D0Nl?���5���4\���7�*�������ꆱ�cE7��MKU=1��R�ߺu�Q��A�Tv�)3��sEgAD��w@w����K�M�Xy�޽{q��W�[n���B�k���1�^bu;�n�W3�녎������a{�������=�=�
O���!�Bw"%̮-@s]�%6qSEE1&�ć����tI*��#r�%���ǻ�T;0����~�G���0i���;F�۳յ]�Ih�*}�u@�>��6&�=L9v����R���O������f=3��.
�����c2ܵݾ���2��ɢ�d���䷕�@�]��]����b���rkn���n�����7ͨm"W���M�umW��T��G�GD�R<�,?�k���L.ve���K��w��ƞVVV��}�,���X�or��7�.]��o�?��O�"`O��=�>�ik��&��s¯���k �C�V^.�,Y��c"{������d��� 	�YA��-X��A���z�����s0�`�L��貳p��Eh�Gn]+_�9��)I��c�'7/��/�D6RԾ�w��T?aXB�0�>��	"8}��@����D�VX�c��n(
��ڡW�PW+t_�)7[�^��$ې*��%Rglhh���۶m�1�M<�:�� "[�ܥǜ8o/{֮�_lܸ���x�(//�j1{�5����uR�>��Y����.����P�V����C]���Yvrg��ףW�A��H�?"$p'�NuyƮ�(��'�
�$�޽]��RD��4p�����3������˗[_�A��D�0b�(�9�0�QX�\��sn���1j��]����b�T��+1�ѵ��	����n@j�^�ve�힀�n��`
�A�������]���]d#���PHn�o��_sG�rw��o~�!�)��y��/����y�@\�1�VL\�@2]ەs�&�hm����g�a���?������~��1t�P|�_L��=}�2�_[_G�KZE^��ܽ\�CQ�U���;KV��mڱcz��[� � x��9W/£W��1���3u�@,��k$r'���	G`��N�����mg�u�X��H���-?�2�L�P?�=�<��δ�=h�m��B�l�%��5D^���������=�\�H�ks��MV-0���u���_o����?�LĠ�C@A��:�����xD~��o�w��.����@&�&Y��CG,�X&���y��puC��F�Kg���j��Ԋ۵uC� kF��x���Cw"����;�@�v�Ђ�I*�{�_�� @�J&UB�t͗H[�l�W\���&�CaQ!&9���h�	.l�V�v�V�_/m�Jb�B1E��d*�r+Ź��@�J�ib7����{�[�>���z+�k���pcu�[:�]��5�۩�kYo��ڕxwve��m�
kyvu�|��z��@����Sb�F;חt�"ޭ+ƙ�k�!F�x2=����$$�nK�k��I4�����I�C9~#��H���y8�<߯���=� ��TU��S��%�h���x#�܆��G2g�s�|�	�۷D~����Ϸ�<�0�F�t;+��G��qd�q�Ǣ������n���.�z������<�$��d������莃ts
A!��iκ�,�曨��=�<L��׋����=h��	���'L���Iж��-��Z�1��f#L�~�_���1:�~n_����9�I����~�8�s s,�Q����'n��V�0�9#�fX:�A�~�����'�����S����� � �����Cѥ��zeZ[�!�x���1r�H�~��I�󤻖�nc,��ϲ1�+n?��!m�PW;�	����>C����.$p'���>E�'�u(.�$�4.�k{t����T����&��xS�p``B�y��aÆ ���8��е[%75",n��3����Z y���\�j"���b��^��ٱ{�'ku�5�ve�FDx�!n׶�b�tm��'2As^���B;S�W���-�� ��Ϲv�]�֟(qn����Y�(U����	���τ���t��qr��#��}�����T߯f�����g��O2�c͞��x�����ԉ���J�y"�h��K�Qo�ќg4Ǯ��nu%�@|��7D�������97��m�sy��U8��YX��;��Ï@���͸��p�M7�gϞ)K@%Ý!��b�Y���ܰ��-p����{$��u����&�tɪ�s/q{$YU(��76����z�Oi�A� Be��F�v���ǵ�B���@��8�O���5��ذu���N��_?.)}����;�!�j܋l�����/��3�$��#K�#q;A�HQ�@?s���B�ݰ@��۽=h��5ȂS/�oO�x=u�D�x�p�w��/��}��(�T� ��0��'Oć+�Î�;@��^XSS�)S��]̞�ZbPc,C��o�E[�S7�����.���1ƒj�^�?����E��Q�����B�$p'�F��$7�x;���Cz%���T���T�k�_�*�O�%��ξ n��v��� �^}�`�Q�PT�������\��`RC������Q��$�?�صB�@m��99��V�]ۡ�k������	��i��p4��r����	��i=M[�-�Q�m���@
\۹�=ۄ?y�Fÿ_g����.�F���}�����u#��?��ǀ�������G��ˊ�՗�[�����#�"�>F�;�#��3�6����N���E8���ťK��g�"?ظq#���j,X��r���w�lrd0�O®u��Wwq�'��d�=Y%	��뢦��,�]{I�NA�lܶ�]�7<q�7ѽK�@��Wn�!^X�6+�ܯ��9l޾�	���_�1�<sfR�{j�G����b_�d#l}�K�9��'�Ͽ��?�y�.%I�s��=��������O�.�]���b����k�D�X�f��k9p ;��Dj8�GL����� � ::�7�I���O�n�Z�3x������?����O�=��X�K��SJ�5/����NB����v[�λ��5C/w������{0���]K5C"	܉�q\�����J�*T��IHRQ�T��y&���Ɠ�>�{�9,\�D�0b�!3~w�D��������3#?���L�k�����ʵ]��K,�YN���t[��mL����k��[�,�6�yU�z,�G�r�:�k��;�>V����.��z�/.��D�y9�K�����	��!��)��=�k�sN	Я���C�ε]�&�6�va>�yB#���qΝ�r�c4��ؿt�H�k�f�	ʹx]����ie�6<��cQUU��=L��<��_�=�܃��??�T2�b�#�mE�3���a�C��*9a庸�n,q�0�bHVqw��jmi�1�Z��j*�v�C��\�\��� Ad�6������^�������0�HyY1κ�D�	��y�bo�;�|���,ڲT��~������&$�ϊ5[�����e�H�����ϳ�`"[�.o��ܵ^[+�3��?D���� 2ژ���U7v:Oo��#��Yɘ/H̍��֨�uuu �v̌w(F�� ��%��τiSн����U� r��۷c�ܹ��{YYYRM��YK�Jc,�uC�Ktq�G��j���{[�������,6�{��o�� �;�$����a#��!}�TZ����$�d'1I$+I�7�d$��90\w�u�#.O`���'`Ȉ�´����\ۃ��|��ѩ��C+��,��*a�BaE�nǭ�+N��[Irm��h�S'׋r����ůlcu��}�79������v뮄�>'ӵ]�A\w�h|h�C��R��4B򤹶s���G��͵=2��i��9�v�db��=�~ma�N //[�ڮ�[6h�����c�?ǻ74yl5T�6�,ʷ����N>��c����j����D���rfΜ�Qz�	� ���VLV�� �uU�+����?a�9-Y���Ѓ{wlĈ��x;ݐ��̙4��kA������>�/?��;�}����ҴQx�@���q�_��G&.\c�+���߸����o��|ab��6�V�s��Ջ~��ϕ�݂�?���[����8@�w"C��݌杦�)�}��m�%��l���!{΋/x�,��Ea��CetD3�x��{��?�˗/���`��3Pݫ'� "W<|(:�����^���V�ϛo��;�?��O��'��*���ۖSRn�Pg�Ů��i�U ���5��\�Cj�PW/���5Ö�ݷ����9`"9�^@$涷�����Ib�un�=I�ﾐ�$��lIhu``��ܹD�S�~|������``q;|���l�c��ipm���Ԭc:]�MgN�?Y쫛�����"�u����Q�61�vW�.+�r"+��k�</�|���wm�9bhe_��=r#���P�Ӻ�b7�IB�n�����|�������;����y�Br�1e��k�t\�; �ṮBnmL�^�Nx�yB#"��qΝJ?�\�u���H�]�����D�^�+�@�6V?���>j>#Sl��{�޷__����o���Dn���ٰ�������I��=�>2�6�#��h��{;����N�#������j�U���Nu�����|EA��\�s�y�_�5K�ۑ��'��k��q"�t�T��.>SGL�������Ó�}�l�s���O��|���3~x?�a��e?�[��u�|���x�h޷�j�S�ƺu(..I�n(��,��Z��������uD/�-t��|��O<�ŋ��JJK0y�tTt�� ��uz��cN8���456��}��~�9'�pBZ����RUK��'��8���n�g�e�Y�Ю��hk�|�P~��6�؄��C�c�=$p'fXUa�IELR�
cb�@��������^I��lpcHgb�~�7bŊ r���v�L�m�n�f�Gpa{Gvm�I�âO5LU(���N=\�#B_^�_G5vu��r;�E���Y�&��z�4���c)��v��]L��:��*���<յܾ�h+m�f	��K�{�إ�#(q����׎ݧ����c^�8�-��\�+�k���^q"i��J�\o^�����˶��:�������
�})�qͶ6ܘ���cW����� �����m���.�ML�*++q����<��>�n�8[�l�n�dnc�a��ΐ�dT��+���$�,�v.i�'r�'�dG���<g���wafM���dA�����Gx���+�����r�����H?x߉���r,��l��;�v5��7�y�>؀l��g১N��a�!��&��a���xqŧ�M6��A�~%��&�lCKH?�s0a{��@�!�G|���YvJ���mRe�K�d�����`�� ��=�0t�p�AyE�ʮ8�s��җ�c�6��G]w�u<x0���:`�}�2_<m�5ƒ�^5C�5o��j�^5� �X��{�ctY>&c����D�VQ�����+A%&�
<W�JR�Ȕ�=]��K�,�D�SճG}���`܃����c�mg
��ԋEe!�!�e�Ipm�W���ڠb{��Ib_i��Wa��ۃ����x�����5�����*�1y�E,�qm��	sN�´d�����MSE�q���}��G��h����cwmO�G+$��3�M����ř�N�v#|�����;u���(ˇv�|um����v~ZiI)���x��g���/��m�z�-�~������c�T$���B�j_;B�J��b�k|�*,x��ŝOVَ]�mFyqo4��ʆ ��f��+-��?��� ����Y�[��/}D�QS��۷}>Pӫ]~��p_���Ys��M;����� ��
0q� ��3����t���;A$����\׀��OS,�;W;�j���=H�PW/t��<�l�K����k�.̛7MMM r�AC�`����]O�|A�Gq��ԣ�?�{�u�_�)��f��ݘ;w.n��6TTT$\��Uc,G[y�����B�Цs��ŝ��"�B�fشg���zD�Bw"!f,D��z�����ޮ^09I*��,&���Lґmn~mW�\i909�ACc��I�1�����"xF�sm��k{X�)k,U��{`�v�O,��ж�d�m�M֌j�4؞�1�z�v��sU�,�vA�m5zP�D�]�kcw&��sq\L�إ�Ҏݯ���L�6�vs��p0²�}�Ǫ{�����x#��<Q$��C�GX#m��<��ˀ��s�o|NL]��`�s���]��/����~0<�H�F_�憄X]ەx4�M��>��P٭;�||�u�L�.<� F��9s�dm2*�|��̑��~}�����b�����l'��]�-[���hii���6,Y�� ���W��K'��#s��'a���:�h87�/�v��VQ�\gdMO<x���SU�p_l=��Eؾ�c��t*�/N==+;�+�G�>��ӽS
wo t�X����X!�~�=��\3,p����X�xj���'c>�9�Fgu�?���Q���-{�� � ���q�������� �T��trl��/�8��_�k����c�]�����ۣ>����vq�j��QҼ	�%}��B�h�Bw"n����ʖ�8XTNJEN81����e��D�Tn�JLR���$U,m�:0̟?��� r�cFa��q�s���AT�\���M�� �����������K�mg>E������{	x�NW�����sm7x�4�^P���	���_�.��\N\ۅU7����J;e�s�`�Q�cMn�Y�Թ��q�?M�q���n��\wAc���wԘ<��A]�M�4�<�]��bqΝ�r�xLu���2���2�ڮóo�h�O�.ە�#�N��O�|�T�����އ��� r����a����R��e�#��*<�;wY�F���)9y�VV�#sa���n9��~#�T�bK92A����k�Z^���6���b���3p�/����	yo���CYIr���⾋�L��{��5��u�qoǸvb�oQaDp&2 ���8㊅ �D9�o+��ڒ�ޮ�٫n}�g�:��mfX��M�|�93	xꩧ@�6�x�|�4���AA�a���Ν��˯�1V��裏bԨQ��W����'��bi�1����n�����cuq���1����8c�-$p'�f�@���PR�{{d[Ĺ=SI�l��:���p�7bݺu r��>y"����!�p=���E�:���*:�y�`5�{���0Uq�:gx���k�(�Uc��ĺ��9�v}[�@V�Ƒ�$ͨ�@���c9�LM�d���q�N��0��Iqmw���&�ؕ��?v^!�Ǥ����ʉݧ���L�6��Ո����r_�]�ݾMi���p+���h['��E�@�GHν���~m��k�]�x�`��"q��(���nM ��k��:-���r;!��wذ��q����{；n��a���q�UW�O�����J*ś�J�X=X[�#�;��ǫ}�A9ae_˙N�J������{6��r�$� �s���-A���4�!}�,��7�}���"
��\p������|r�3{�p���SQZ�x�g���W�=��;N���I2&� �H�!�Ѵc�����¨�vYܮ�ٮ'1�E�{�t�a�fX~m�����{�����`ڱ3QU�AA��T�N���_�ĴD��4sÇǘ1c:DM0������ȝ�Y4�j��"w�nh=صc�vȋ�[�7�o���l��	܉�`C��7��h�qo�ەU|��+I�̾���4���F{��'-q������=��)@;�]��E-f�\ە4m�����3��*����rm��DZ���]����.�uն�A@����ۅv^�튃:\��?�2-ݮ�B�L��+�Y�)e����CP�!6�v7$�����ӵ�_(Ǐ�qmW:P���9�t}A;�r�34���t��!�h�+v������<�6	��kcҋ��i��~��sǝ������a��\p�1%�:��Bl}q�+ұ�;�	�D���n��udЋ�cuqo�ۂ1������AAѸ�/�BE�R�5k:*s&��OO���~	D��ѵ��W0��Z�_;n�����?إ�����ぃmh޷�Jsߩ� ��û�F���+Ƚ]��5�PLuC�A��{�,��a:��|uuu��k�?]{�2�+:c�qǠs�
A��{u̜3/�g)���@�&��l�ܹVݰ��2�z]�u�\3���a,���urg5Ķ6�����l="�X�V�cM�n��{�+!�;G�mž��R	纠�{&�
d7uhA]b�Oܞ�$U2O:2����Op뭷��]���t�г�����҈��֎\��刂u����]�)\۹?�4u9�ؕv��]�]ۍ��U�����d��]�7M�b��f�1Į�7�b��BL������N�4�X�n#n�,pm��,M�.Hm?���~���yا��� ��v;a���>1Y���<b�&��B��34�|�F,�������h�u�]x�j;uuPU���ɏ�{�ņ��A�&l��C=�f��ɨxWA������
7�we�sc'�l7ޑ���῜�]��PIRr	+[�>���� "�{�W�?�n�8q�HtT~s��X��3<���s����NEuebfL,�8��ɘ��9��Y������#/���ʶ]�Ի���i��H�#���~;JJJ���Q놼9�ƹ=S,�fh8�<��\7-�a*L���]w�����~J�X9L�U�s{Ii)� ��KeWs�l��ߥ�U�Dn�j�*K?w�EE��udc��my����� �ˮ�uDo'w��\��b4wf�5��P��F.��	܉���^���Q\\�8�j�vI����E�^I*х!�I*�rcH$���@�7ov��"7��f��.]���;���Nx����.���R[�PU��5�q���tI1�5�A��^^�/%v>6a�V�/�����9�05����>4m��x#�rx
���������z�,C#�v7��s��K}mr>�����)L3���v��?)&k����X5�۸�MwS ۽ɑ,�vML��¾i��ڮ�kjڨ󙦦/�k؇�ԗ��F��Epo���U!9��qo
Pۤµ=�	�$};nZ���������Ea�W�Ax�#,��#0`���AAخCtd��p���=���]k���>"w�I�vd�\��߂��]'n�]t"��]�8r@^��1DeA��O�N���%�y�c��v�� sm��Ÿ��3p�������Eq�g���[/�2���l�k ����4��;+)N�?��	d3l���۳�ݓ''�מ�|{���һ��#��?�q��ǀ�ܿq�C �x	���lG����ۣ�c��v�K?�3/n��{���H�Y9u��a<}i�H=�G�F}&r�^}�`���(*�QM� "(e��p����ŗ���- r�ŋ[�X'�|rR��T?�֒!����.�b�i���Bc,q�g��]qr�pqY�]ú"o �;3*�XC�B�0��ɩ/q����O�ŉ!LbI�lvc�4I��<{�=k�*�}�-X\R\����qڙ��sm���k�4]])��$�ڮk��̵ݔ��b�Ȋ����z�����nM�m���,�k;�Ů�7��r���K�C�3���ʾ�d�vg9�}��� b{�BM~P n_�Y�ޯ_ �\�=�o��R�����(�SW���a쬯���Y��^D�m�6̟?7�t�u��L6�,��69�-�dM��΍3�ލ��^��$��aC���wqw�T�=�yz܂����� ����NDM�J��~�FlmmDG�u�A�u��a�оxಳPեS\��n��Wp�e�D�Dl����?�N�6*��%�%w=�%�|�l���7���2}t�}}^߀��.���~���O,�Y��a`/rq��֝�8����n�sLm��{���$t�Ź��ꌱb�z�cu�a��~�!n���ˠ��1~�$�!� "6
�
q�13��+˰��u rV/5j����<����1���\�ЮF7�r놊1V�=�sHk�常kF~nڳ�kz��ۨ���11�O��m��U^"��M�Jp`��r\ $;I����1<���x�!r_�U�{�Ĵc��~`ǂ�ID��'SigJm�����'nk$�pm��r�vL����r})��ӽ\�S���_�I]OS�N�=bvm�׷�=�ߵn;G n�G~���^�k�kh"��E����+}i��z���k;�:�k��wy�����q��7����웩umc�m#)#�vq�Yv4��i��\Ѻ�	�vZ�yd(�bWVO�����6�4Sm��k{����ݿ4�Li�M�rک(++�KK_ �{���k�����|�C$�R���U�9�~����v9i����&�Z�)��]qq�$���}{�0��'�^C?� �c�|�g8�����o�sY|N�SGįΜ�k>"8��;u*���p_��⻞���|�J������gb��~	����8���sf䀽-����G��:B��{����_�g;�� ⥴(o�����#>s�>茱���b� ��l��������d ��Dnrȡc0zܡ � "~�o�I3�DIi)V}���c�Ν��k�?Ym8��]��e�1�Xӷk�|��K���������q;g�U�j����]?�j�Ņ=�J����D`���
������U�ƿ������r�C
&H#��@�QP��S���g�)>�PCB�"�  �#%��!���{��gvg洙��;{�?���3�9����s��N\��	K��T�4���O�>�k#U>�1lٲ^x�u 
��	㭡���pEO�"5bL�[����նjj����\u��<�N�wm7 ��U!E�����VS͚�#��7v�>vfitm��)�Gl{9Z[����J���]ە�ںK��R��:h��@�|��qb�?��n'�w_�{�;Iǵ�-��R�_I���vn�X�	⡖e���;�dM��o�d��|>Mݵ�;FW�x�|��q˷R%q{�\ۅE=�M�/n��}�|�XT��#�D�z�jx��X�paV���J�q�<�g�ȧ~#�����%r�l������g?G����.��Ka6m�ЊIh��� "��q'�q�_p�/NFiqr�����R<�n#�[�1���z�|��
e�wy�G�c~��A�����W��ǭ�8���r^�7�~y��QH<��&�ꆇ�/��Rٟ���Ӎ��ޅW�ߊ��݊�ތ�#�%�H�L��U����^���]3곟1Vq{��]g��Hg`����'[����/�Q����þ��AA����棢�o��D���k�����g��e�O0�r�C��}��X?`d~?'p��u�w��P5�bn�:q�`�I�ܻ:;q��"<@�X��Y>���!K$1��0�E1���qJn����O��7R�ȶН���Ӄ?��ؽ{7��c��)Xx��@C:7#�5M��dE�š�S�1De��!���O�k{̍ٔ���G˺yj��J�FخYO���Nщre��k�!����
�5�Ǘ��y��+��垟���Υ���޿��^�w�ܪ��q^���p���I���k��e���Η�
��:*/�8�m��d\��� [*K[?a��fjˆ��͖&�v+I*�y!��������ǉq�L5&����ǎ�ˁ��hH?ڑG��AU��]w�(,���q���[V#G�L��(Wb��920��}N���b�un�s?��he=���)���Hr�ˑA�Gһ�{q��^ܳ���&� ���>����}�8��x�:�.����{�X�T���A�(/-AMU��`>a���!����DZ�`��﮼w?��¿�>1k�e��r^�e���f����f�}/ZSX��W�����,��zz����]X��v�۰�Y������� �DUU����US,Nܮ�7���dq�W��W��o�YB����0_�}��Gq�]w�(<�>>�"L�1AA��}��FIi	ֽ�J\�>����kٲe���D+��X�'I����7����ɽ�3Ų�ͦ-V9$r���Dei�5�`�ƹ�n��f�Ht_�i��+nGLX�����ah�ґ.�믿�>�,��c�'f�����"��q��J��T]ۙ�Zjߢ ҍՉzUQ��d�fK�Sa��	_[�-��&�ij9�
�ڮI�|J�k;��)N�}=�=i��Rݳ�ڎ811Et�]�U1���-�w�B�Vl��|�����]�{�趑��̵�Y+}y\������8/���}�G�.��umO:.�^�{	�z�k�o����tt饗ZB�d��<�l�JG��|7]�n �sC��m�*�9��#ߣC��V��{d�س����Mt,�w>ޝע�t��bƄ� �H�;{�ƍ����4��x�7_??��>�y3��3?�r>�e�(+G ��*��xmJ��PUY�|/���Ŗ-Q�3AWw/���w����|��%�q��?�W��?܁u3[;@�}�]xw�nl�Q�rg'��a�]訇�oȞ�>�?��5��v{�g~����3��)S�fX^u`m!��F}.<��h�L�<	AAd�i��DYY���t?U`�������=�O����ڤ����?�,���K�3�r�<��#{�*�&w�g�~C��	ݻ���||���D�Cw"GN�GO]��+D������SQ���f�~��H�x,Be͚5��`����ܸq�`)@��V(c�Ce1���t�vU���k��)��G�:!�*浳L�k�$�t�5b{x�����
��ɔ����Z,K���x	��q�:j?�~w9-Y�v�����=CSW�u������J^����oۿ��{�u7�^���h�m��҇,w��B����u\rmw�SW��fj��c�8M^ʺG�Rum緛Z-7ͫ�Z!x�'�Tc���n�?z4L���$�>r��s��o��5���F�!
�x |0�=�ج6Fe��)����J���ЃZa��9�H�5�`�5Ԡ5G��92�D�asS�����������2���'��� ����[ǾG�S���'9�?�:^|g3��>�[�@���_�Ýxr�F�+�{���C:��/����+�P`���ۺfY����*A�M(+/�>��vI�^�هX��E��8�3�W(��E3,�Q���X6��G�L^Ab�ϬM�.��={@�;d�2�W� � 2�ĩSPRZ��|���
��;w��/����#S�X���1�"a��B�o�1��:�s�>�t�Œ)��Y�oh����L��Y���M��� 
�qVY4n��0J�^������UR㔟����@��F�t��ә�Wlkk+.��tuQ�D��\�g̊�L��ߜċLݵ��_�ӶjjSqmg�+u
�k;':W��b5�t[�-��&�i����Tѷ>��ԕ�Y�v؛Q��z�{\��X\��G��!�����z����b��}��H�rm��;���ә���f7���;�^M�\VԵ]��d̵=�(�J2<c��Ja��]z����k;԰��l���g̰D�ׯZM"��������2eJR�B��ؔ��h�t/c����]��.�C�UE�Zq��Ƚe�N�=o�� ���3�t����0{ʘ��g���9e9���Z�aOcN��-xs�N�#���w�_�Ԃ����ۛ��oEkG7� �e������v��]/rWG}���F{֚bA�Fd��͇~�t�h�-�܂�Da�\d=r9F����	� "[�N��G��=��WQH<��c���q�'��'���X��%�1�)�3<��Ϫ1��/F.r��t��Z�;3�ڊ����!�;��zѹ��奊���E��B�V��%r�5Xɓ����'�	�����A���꫱~�z�żE1�3}c�փ�����kD����WY:��r��sm��q4���J���R��V���]ۅ4�'#&&���|B�!��7ky	ĥ���4ݮ톽w{�]ُ�};]�u�y)�ȶk�������SW��fj��-=���f��F�������>X��]x#n��f�1�um��(w*��7�;�������6��Ι��ի���	�0hhh�^e��S��)G�l6\%3_����� ��&7T�C�V�C_�5�`��Ƞ9Ȇ�7h7Zͩj�ۨAA�	����߁G.>C�+^����`Ѭ���6�^6l݋��>�Հ|���מ{�Z0#-�=��&���ۭ}� "Y�Ֆ��a�5�,n/��s�X¨�na�ϰ8��]~6�3��"�}����������w}�pQ^Q��>y$�
� � �˨1������z�d>ZP\y�8������R؞l��L`c,��19c,n��1�_�!��yc����3f:��E.�	�	_�.FW�f�Qʧ�J7Ġ+t/�:0�6P�'���5���T#T����?��S���;A��}f�wb%"Xg�M�k;4b{��7k�������ea�.�Cܮ���-Ŧ�ڮ]ayC���)�Bq]۽�n8�
���.&�:�r)��[q���u{�uϪk���),gW]�������1Et�\ۥ��s��v���͗o�?��o��:!9����Z��Z���o�dEw��ȼk��y�u�J���#l��튰]:���(����RX�eh��q'M��g~��ttt�(�}�Y�q�8��Ss��Hl���3�}XkD|��� �2XS1/lw��9E��~��ū;�� ��w5��K���?;�j�L��?{0	��̿�݂�~w�ۑ��Q�[~qrR��:}�|�w���:��H�ie{��]�����>�"{�g�ɝ��B������C8����ܹ�:?yy��گ.�����絎H��
��$n'� �2l�p�z��#���D�CKK�e��r�JTT�����?�Krp����XŜ1V��+�_ا1��c�X��ϳ5�-T�(\H�N�r�.t���T��*a��"w�Aѱ��ӵݯ�J��S��r����'���*�V�v���,����Ҝ��Ⱥ���oTdaӆ�R~SCc��T�4�����zl[Kkdj��J�bB��8}��nR��O}�"��G��PY������V���ݝ]hkmX
Ww�j�~$C^>Jc]=�wMAЯ[V-�õ]�َlV��:������TѺ�v�W� 'ώX�}�޽H�7�����{��o��]󒅫]��8`���ڍ�ֽ�U��_�3L_��6\^M�MVC{EE�Z��e�x�H�y���k�N���J�'xd���ղ�q��C��=��9���ȿ���_����D���&�M�����m߲/<�^����,�!l���:��ް�"1�d~	��D8d�x��/[�1O����MUUn���}?���p��c͚5�?>fϞ�5a{>96��U≺(�o��*�F+~�Ag�A���;�Aލ�5^M-݋W1A6yy���s��	�&��g��VaOc��">w>�ι�>���!�5y.8�3?�&-�=F�v� �Ē��hil����>Ø�@��Ήܭ��?��9�~C�Y��/�Q}�:��e��o�������
X��]n�����\�h٬�}��Q=x0�R����a��~��}9�3s��l�9\��o���?��{ֶ���ތ���9��t�����6��|fϷ�kj��#���OjG��=_�\��{,��_~7�|3��o���	c�`��r���3����X�Q�Ց�������7dϗ�џ���b���xe�y*$p'<�:�m{7���<�Hk��5R	UE���/r�7X�7R�+v���F*�h�b�/��R����J[[n;�rU�-~����0�A֝��]���L��1M�R�:3q��ӼJE&]�wnݎa�FX�Ysm�����L�9]y�.�Zw� �v�BN>L���Ԍ1��i�Q�u��tm�Ҹ����6�������L��~�����nHu�%n���'�f�StVVHR��OV~_&0g7��ǎլS�������ob��k�w��vLS�Ѭ�]'�uҭ�[��Ü�x����K1ޮ�R}4y��G:lHdqE=��bt����}�_um��c�AĲ�󄜏��?wj���I�N�����7���s�㜼}�ĥ9�}�����x�"���A���� ?�Z�M}����>g	��$}�����ƆF�ܱ����, mRbq�.�5�_���Va~.��}t��g�v�����o�/�W_}5��N�l�,�3�D��tVJ��*^����M3����1�9��e7���,�8�m!w� "|\p������5ytB˕D�����_|D������͏��>�|�	�%�i��_�l����=�)�'"<G�����BW�?��3���F|v��ɣ��K��=ڳj��?+�Z����^z	w�}7*++֮$.S�|V6ۿX�D����ee�g�t�6�XS��������}�Y�֦f�ز��%�sU~G{������rA��}.�omi����93���[�}.޵)S474�쏶�\�ߤ��=9�?��|�η��o66���b���{,v��{,v�+c�T��ڵk-c�y��eM��Hl����}�����~C3j�U�:�������џYڔ�x��Y	�	OkE{��@%��{5R�SBcU�!}��O���*H^?�0��~�;-[�	�'i�7��2��}dq�)��R9^"Xi��|QZ�r+���uub���Ԋy�,�dK�*��v�zz�(�׏��\S�=b�)�X]OS����-�*G#X�t�B�(*��d@�|nx���3�P��M�ۻ�iĄ˦�&T�KS��q����)���M�:Hߝ���8��4���
W��ԗq�}YF.O�y'G�:I1^ǵ!�7����+��'l�XE ���+����F~�+u��XIܞ���;Ǝ�
�uy�j7��po��`��֝8����G���}C��(���z%o��c��[g���/���"��o��n�g�yfʍQ�uIHn~b�UjC���{.c������n���F+ޑ!�|�r�o����{)ƚ�Pl�@_�:d� "Yz����5���_}%�e�T��H���|���亍�w�%ng��_��/$n'"->��-(//wG{��Y4ǒ��,����Xq���Z��T��G��н��]t��7l[��FC�6�o���)�E]��O�m?��
���rnO]�h����	���~�����,���lD��!Æ�����wo߉��T���Ps��=�=سs�M������n�qֽC.��g/U�5�`T혜��K�۬�oǌ�'~�a���{,���=��ٔұ������^k���������J�h����u��^����ϱ���س��6�*��-c�g7��{!BwB˾�Jвw��HU�i�����8��C�'<�[>�	4�F�x�ݰ�μ�oߎK.�$go����-=�G�ߛ7N/rԔ�����cz�y��{���8�|U���������q�,���1q�R''v�����^r���bE�v��'N���5�)��[w�:��py�N���ݽ\�Mn�h�*І�{b��鬻#l�S+���� .�� v�:u�����A��&��þN+y�/����ߒw�1�'�;�,#u�v]4�=ͱk�I�~��Sm���q�D�^yi�K/����M(i�tm�.�[sm�>N��P���ر�cq�����/�\qr'�ɚ5k�`�|���llJ�|�gc�ΫїO��^�̱�k��>G�ss���!��*{�A�(�ڂe�F㉏��� �����51o���Dr�ߴ���;�yW#
L��_�]�t�DD�C�w������r�a�=�Ї���L�t��'p���+��>�Db�%�_�r%>���A��jv���ȝ � ����<��������BG[�D�D�x�w�j�*�s�9NZ>�zŦk~��X�6Ag�e����X��B�h�c{�r�X�1֘~f�5���
�Z��nBG3�@�5�7�`�ƅ�gx���Sh�JW#V��3%tg'o&n߳g��c��'NQ�^uo��To��5�v�d�_���2O['VS^RS'KY���g(�|>�P7*:��IYK��5+��n/�U�d %�v�X>&�Ӳ����CF�Ʀ-�6��r�tm�rU��vx-�y)@�}�-(�sI��7�2V�Cm�tǪF�ĵ�9Wh��������rXk���<U!�['�:qQ�!��Ju�
G�.��smwʉ�D���v��.Mү{<�v'�K=z�ɜ�W^"�0'	v}�uס��:m�M�#\6_==��bG��|f�~����8�n��F,ٽ���F����QZ4=�I� ��y�J�㮜/�m�i���n~��N��cC��������GGW
$n'"�9�u(��pD�}����E��%n��;��o(bpSz��tdZȞ��֣�>����� 
�ʪAX��$n'� �P5�ˏ>
O<�:�;@���n��2�:��CD���|Ay�|R��bi��B���1Vt�g�K�7dZV�+j�Պ�'��c��-�� �;�0��-��Q^^�
�97uhAۅ!��λ�;�ũ	�E�g���5�/���;{�1���ŋ0i�%=�`�9�͞k�Nڞ]�v��Jz"���>'v$��k�'nc+��k�!�%�|�Õ���\ۡIc�ޯ���eε]ZQ����+ʏe��kҴBr�r�K|��P��-(����ė�r�r��6�|����`<��N(��A^w���O�qm�뮋ќQ���~�E�I؍���]q��e�e��0�]���V[[�3�s6nX�D�ٰaV�^���NZ�\r�0�W?1Fj��~�~�jCUl�Aٍ��_�;Ϟ�#Cql�����)�xhcn�'b���D����<���`F�e�*�@�=^]|Ǔ�(2�iv-(H�ND��*3Pּ��!����Ms�
�~� �vm�!���Lp&�\��e��P7�޽�{;QT�Ï>U�� � "0�����'������.��"̞=Æ+���Ԍ�T݁�o��1z�2�*�:��L��џ9c����(-�EO� j ���P�V^���R��ʫ�J��^$4V��z9/$�ޮ�a#U�n[�nŕW^	�0�w�BL�!K튋�/T�ȝk{t�ZMS�������㺶�����i��XE�K׊�ݥ�*j]��b���zF�ޮ�J��8G-ĩ�kY|*q�:�{�J�a��Y\Z/��=�I�ߚP��먩;�]ݹ�$�[�K�\��U���+˽N�|��a'���.�\۵Ǌ�w����Wٯ5��]���ï�]v<����
)����IQH��ɣ�@�y���������4�������gƵ]9���89�HԵ]�&���ƍÂ���g�AgG'�ps뭷Zn�-�HcP���.���CN#,�]��*�y.d���	�9n�#�0�"iF�VT��GٸA!�/O��������F�$-�]8�ҿᡗ��@���Ad�����n��X�7��;,Ҍ���%�<ڳ�g�?���k`����^q�زe��SQY��>�Ճ� � �p��߇}$^x����?����;�<'-�����w�E�O<c,]ߡ�o���
��Xa�g�!?��-t���Ċ��H�B������hi��1k�
4̠�&M��P���4�ܔX#�.-�������@�&n���L!-�`�9Ƌ��,UѦc�C����f��V=]�!���\Oq�R��>A��'o��]+nW�6�sm���n3��{`�vy=bqZ!�	�0޳�r mw������|1�:De����]KC�����v׋�uu��@��v��܏!�4�i�u҈˕�b���դi��r���\ە��p�7u9��I�lJbwnI��ג�r�r9��S*G�Cp�vC>W��v���k|<AzPѺ��K����v^���4���n�Yumא	�vS7�f0N��Xu�U���^Xc�e�]�U�Va��#1�� ��l�O���{�Fvc���rC�W�#Ck�*
�P�>wu��*�� � B�3olJ(���xw�n|�wb��z$H�ND&Z��4}y.����"w��]5���;��GQZ��ӥ�k�������?����O��Cj@AD8\S�IS�ཷ�AwW�ps�wbɒ%X�tiF�s-l�W?Nu�!p���}�|��)c1��~[�����)�bYi%(i�F�X	�	�q؍{�A{� �E���=��X����v&8O2B�x��ٍ�����#�<"��p� nw�D�*�g�ε=&DU��
��yJ��zK�&���IF5�d>]��<�SsrfY(�m�vE��H��89M��f[���k��fH�خ���%j�����u��i�>�Vwa;p�r���A���>ism�21M�y�A96L��Rum׊����~KS�����c���C����+�,���.�7>�9�xM�8'&���n7ϼM5&��Jݳ��nh��0#}��n���S&��3���W^�����w���7ވ��:K� ��Ʀ�6f	gc'F���=ܠ鸷��EG���{�v�A;�Dh��6V�i��'������ � ��6���vf/-)�s�?���s`݋�������A�d��^t�����\�3�?�+l/*�o���H�_ȋ�S�ӑo}���֋�D�)�(���k�AA�ƺ��O=�(c��G�r�Jx���1V���ҙWN���?�zO��P�7����r�����E���Xv��m�%cu��������
��0���&TT$6Ġ3��5���D]2�H��F�d��*k��ݸ����E�?��= 3f��T���k���#�e�]�����Uŭ\���b{���x� W/KzF؊f�L2���+�Պ���W���o�m�vC�#�eҵ][^��k�sw�<�����vO��'������:�i���C�ε]�&����u򪳝&���Q���~����2�_���/Ɗ��>�c�P�Ѽ��)e�v�r�1푷t�s�RqmOPoh..��	�,4?�u��ƥ۵]7u�}��3Nǟ�����fn��&ˑa޼yy#<ϖ�]l�RNx�=�t�����z�8�����E�؝�t��1w���n�:bp�� � �P��/�:�1���ƿ�݂���ćD���i�)��٘g_�7���h<��C|������ ��3�����3,��P�Ct�	��7ƲӴ}�|?!�=��ܤ�/}���O�~��p˖- �MYY;�H:AAC��ң����z=��e�B�>��իq�9�8i���:?k�XV�~�g���;T�M����+�+�����mS,���Mh�F�X	�	�q�t��C�Z�R�Hh�*�3uapO��T�\��ǫS���a;w�n�k���X�]�P�傊���v^�TH.�n+}ե�� ѻf�.�N��m��(N�N��m�_G~�N�˭��zʢ]N�,e���x�m�nw?a����k�����B������lx1-{��B�|�߶u��A�EN]���Hu���3���$]ۅ�\�XT�|�
��.}�v>��])KSv"������Y�sm��A�;/4yl��b���!��m���k��@0��',mǩ�]��m�;0�/i��3��"��3f�?��_�a��A��q�%�XV����,���wi�V�Fl�5ܠ����1D�)�#ϓ�1W��"}C/r���d4oCu��vӐ�AD������j�߹�^|��>+e�ۍ��v����`B�E�&8����6⫿�]��b-A����}�CB���1���@ߡ�)����?/�}�٘��3���{�n�$��8���AQ�9K�<O=���+��v�mX�l:� ��0��X��D�o��w�>�s/B��X�����w�s�������� �;aq���65&��n-�5R�\	ۡ;щT�6Rś�o�P��?��x��@��I�L��E��A��1^d\�a�;5ǜ-����<E�nih���=Ĳ|^��;�IU���vN�n��B��M��qZ�v)����&�|�����ٹu�_e_T�3zlh�$-���\']�)I�����>�����)c���;���%��b����/�xݺ�ǉz�Y���9E��[�����Qʇv�@��bz��O��UwUH�َ��-��ڮM�^�
˵]'��s��8�?���o�DxY�~=֮]�o~��ƞ\7,%���26q��F-��
���*Sh����|�L�Rc��p�ݥƪ�'��!	� ����G���^������-8���h���_�Z������^�@��7��ݎN���V����%c��"Y�n����N7�����4�J&�\�oii���^j�N���/Y�#F�AA�ɈQ#���C��O[}D8a��]t���zTW����?�=c,Q�K֐��X�)V��H/p�0�b�@���
�㍽����:18�TE\#U�\���xRmJf�\ͯ�����p3�f0.Y�|�aTo�׵�O��!���&�Kл��BaE�n�[�4��J��L�T��@�rrf)}�^ +ocu��	�!��+ǀ��Ų��-�v�U2�P����h+1N�޵]\�%��y	U���F �"J=eq���,\2�ڮ�G�� t�'���S'S�K��������u��Bs������=���8q�N���M���_�v�N	���'4%�OqmWҌl������ �������DxY�f�.]�ٳgn�����D���rc��A�������"O��wc�VT��G[��p� � ���RQV��"�Z;�?��⢤���׏A]s{�;����f|��w��� ���|���h���T�c��j��=kj'p��<�����L���W^y%6n�"��}x��%3�AA6��cᡋ��g���&��lذ���;�����Z��	c,y~\c,��t�c1�����y���w�
Y���7�r��&������X<�-���8.n#U��*��ʷqJn���8��H��<�=��������A���c�`��I�}�(���9Ƌ��n�j='6S��U��q�A��:�3'���5\OjEܞ�k;�tS#Xw�)�]%q}]YA��pc��Nŵ�]uw���^H˵k�U��.ޏ�u�^s��G+l���따k;�oͱar_��BSGSS~����o���I�g�U�kFr���cM�;�E��=�d�e��<�h�9�+ŉ)���#o��ν���]�+yk��� "xum���C�8.ۮ�"�[qԑ�����>"�tvv��/�5�\���2+-^�O&�g�1K�?O��nP�ˍUѡ�}�u.��'��� �PAw�;Mm]��G'��,��v;򧳎���Mx��(D�z��[���� �L���{>v���
}�v?bQ���еܔ���L��|9��^��w�"܌?�LAA�IS�������2��r��7cٲe�;wn���0c���ÐF~��2�*v�
���c,��=f�U,c�l#c����ס3Q�v������C�Bwم���J<A�T�\;+d"� �T�=���^�e��X�|��%���7<�]�%ѩ��*��h����D\�U��	5S/����S�����j���[2��.�O�n��(˺	��,�k��jƅ��Hٵ]~K�g�:vE�}���Y��R�ĵ]WwC��Oݝd9��\+nW�+��>1�F2=b���v��5�����oH�k;���q��
�w���_�#l���C��h�Τk�����\U��W�ȼk�P3vĩ�]�R�Zk��D�Еk���m"�殯��L�m'���c>�)tv��ǟN֭[���'�|r���1K��3��*HW���+w^�n���5V�V9HA����bTU����׷�^z'�����I<�<����J"�~���ذu/
�����6����A�������k���X�;���n��eO�����퉎��3���u_����с�+WZ��Dx����}K�{A� � 
�i��DWg�~��G�+dzzz,c�իW����JK�+���cI��ee#Ic����ݚ�ѕ�����
�pO(AkSC ��"n�x]#�ށ�cx��❴��%�L��Lv��Hu�WP#U��<K�8�q��#������]���Sqm���=���!=�j9�n�b��vmc^#-���++h9�|��2G���z���(���R�'�ڮ�]#����ѻ*u��S�{h~7M=u�U��Ǹ��NH�@�c&]����Y��Ԥ%�ڮ�C�./h�Kε=&$�~�x�������R��si��)�A�������}�hlh��^>�����.]��'�B؞�2�Jb�i���<���L�o�*�L��+b�T��U:��&| � "d��c`��1����ڇ^)8q�́��%��;0����~�����R���C�+q[d�������ЊB�����_�B�v� 2JM����͊s{P������-&����/t�3�E���>B��7�x#�}�]�e���a��fa�R�A�@d���������p�~�z�y�8��R����|.�u��E��+��G~�`1a{��	ڣ�����hَ�����8�	�8��Б�{{�F�D\Dn�|�T2�dc�ڵk��*ĔW�c�'�@EeE�Xӄ�����ѩ��*�o[۪���T����TU����.
x�:z�]��b�?�sm�qL�+kF'\Y�OS�1���.�)u����k�f����[���-Kֵ=u��&�����;�V���1�Ƹ�t�!�/K��Z~|�v8y��v�Ÿ+���>�y�C��mq��[D�������ܥ����#l��+�j�s�\w��HU�_�Fx���]Y�D����.ot�?q�u,l��~q�l��]�ߓŴ�qn�j\T�{�i����|��Fᣱ��V���矯m�	[�S2��k�29�{"�U��]h�*r����|����^5o��*� �����|�q�A3����O�1���=�k���es��`���9�z���S1e찄��8z(n������n�(���{p������Ad�#&�讋���7�>���Xv����v��]���dK��}���n��&�e��i�oށ � b`3�������?N�1�a��)S��0]&W��ɩP,
7�3�|�?�}���Ϧ��9���XEE�M�lc�#&�1V�!�� f��R�46�<%�v��a�I�*?7��$t�����*İc���Q]]�g4�k�c"KU{(ƈ�T)6�k��CJ�햴j�ᬧ�W-'�k�R!hE��t[�.�BJO̵]���5qirm�Y����|����-FYAF�,ʽ>`h���d�j�f�������|�#���\ۍ� �?��j�Ǹ��NH�;���:i��/n�wm����(P�v'��Ƹu��]�#n����Sz��=��Jޚ8;6��rm7�8S�(����f�!V�k�5�V^^�o|�t���Oؽk7�����bŊ�TOk���^BwY�n7^ɍU	��G����:qsq'4� �PP\d��� ����������t����s��ĄM�=h|�������W_���D9`Z-V��E�����/�/�m�ی�Ͽ�� ��$̽��qK��Ŏ1V�3��ϾCO���gܽ]G����W]u�5�3Nj'����� � ��`��ֽ��;A����6\~��袋�}m�"l�d�d<c,Y���=S�c%���&2�
7$p�L*�k���s`���{;�He(U^0�*��r��#��T��r�J����l�?��e>r�o�i��&�dq�.9�Ft*���*Tw�̸���Yqm�V�R_)�]N�,����n7���c8�ʂ|�ZN��J����v�����0�:����'C���o�������'Pwq'��;�꤫���v�D��G�n]ۥ4�~X2�ڮ��-����������-L���@��v���$���/����	๪�/�CxT��	�v�\��k��K��:�v�hs��z�Ĕ��Y)	����TUU���9�^t1��@�v,���bȐ!����g�1˿��m��j����CT����{o/�^B�UD�2a�JK�-���&c��J�o��w<��{��Yh|������;��9h��Ə����]��r�g���,�eZ:�0��Њ/��F�����h�Ą�?r�t�����\q��o�/�}� rCԽ���	��q�X��X�s�"l<���M��ԇx���駟N�����-��}� � ��-z�G���"|<��x��q�1�d]�o~>c9#?'`���yW��)VPw���rq'c��B�ʂ�%hi�Gyy�{p�xQܞ�{���
j���X�T��Y&Wn��w�y��d�!�0v|�oLT�/����+�NI �um�3Ј[�<�Y	V//��Rw>�C�.�Vź��v!��v�صH�k��D]��
*�&��.�"Ĺ�u7��w��K���ڮ�ŭ;��h���Hڷqm�z	@�N��vy��5�cZSǴ���u
(���F���oajb��,�1���+uJµ]WwAH�QwUH��1�KjLJ��X/q{�8�е�[�ƙ)�A���k�s/96�:�L\v����	"\l޼k֬�w��]�F�|l�J�2�J���X���[�^�U�96��P�:#���I���XE�5O���>��
;��d6~z�
L�.�;b�4���[��f���?s���S��o�l���C��-3zX5���C^��m��76�v������ϗ,�z���'{A��;�B��Q׌�2&�����AD����{���X)����Q� v7%�ޞ���t�w�^�^�D8�\m��\RJ�� � DJ�J��#�����D�`��W\q-Zd��曉U�c%��n�)r�Xd�^�	j�2��%��0�:���*�{�,b��C/J��*_�t$�gCCV�Z"��7� L����|�"'#K<���p���Br>Nl�5�vM�Z�n�2�xq�R'U�kIU�FH�k�4/��d��٭WC%.��	q�&.ݮ�8�����O��ƚ��i��I�k����u���쥮ʊA�T�A�(��|��wf��?R�^vC�3"����n���F�����r�ܴ���a]/���"��RkYLyd~wOtxy�sd>�E�|K�����:��Յ����Չ�Ύ��N+N�}ma����7Y�vΑ\�7����k����|9v�&F�p\�5��@���k�V��#X�]�]ۣ��_�L��k~�X}D!�u:�
у
�����Ԏ�ӿ�-\u���y���z+V�X�9s�d�a)O�,��XŻ1��X%���t/�;���k�*nۆ��q���n#�0��+��y�w�����G!QY�c���N<�&���Ԏ�{~{��˛�~�.�AO��('9#�T��e��a�ܓGUEb�팦���bdGW��f~�Y��&���'-���͸��u 2Ϥ1CqǯN%w�	�O�\������"��=�v�з�Px�4�I%�����o�5�\�]��8����C�\���
1�`״ʊ����#�GG�g�[��/Bww7����Y�_�kA�GEe%�F���#��۶m�7܀s�9�IK�p*���d�e��ߓqq�ͱlc��'�$c��A�ȬQ%h��k5R�B ~�AU����ۓso�?a����=�XW_}5v��	"|L�1���㷟�"�Ћ���/:�c��G�v[L�&�bY7O��Z���]+��딄k�����Ă�����tû��]��J�ڵ=v\xם�QL%��++/ð�!�\��j+�4#7��0��g����hmnA��]hkk�&&�ʦM��أ�"U�5���
���<�G��¬�k���(vg"��Hݙ��n��o�p�&I�k;�����	ۥ�D\��"yE%m��q>�����B�8uW ��1N�Fx���n��d˵=V��T�q=���j���3�A���k�{��`�ҦϘ��N=���D�`��]v����:#�vdϖ^D�:ȍU@��*/w������ϭ����n;2tuva��"<�)��� �@iI1�;�8�ww��u���`�	��;�Ì	#����U?:KϾ
Da�?�L�ńQC|�>�p���i��ooC}s;�ʲ�Zn����:t����/��-8��	-�ne�x�g�������g�ԅl�g��5?>��� ����$�ִM�;}��bw/c,�_���h>C���X�\���ه�5��^����7���8�kj@D�(�\�BU� TE�V�~���43f?w�6����L�^QQ��.�0��?��\��B���	��2����c��e$���2tv1s��h��i����s�$3
imo��cvt��=���j���#�ӏ<F�X!���o����Ν�R�\������3��xc,��P��{�������cՂL��	� �մ���k��pq����f�wg�wo��d��6P%�Ho~>�5x���q�=��#ǌƼ�j��+�hĘ�5�1ѐ��\�*"��H�õ]�rBaW��;* ��cˈu��s�Z��<ëRV���p���u��f-�O�n���+��,ȧ��,8+$9����3���nW3���\���q�=���bjנ�(Byi9fΜi��Ʀ��>t��[C�n��c455��"�_KK�5���#F�@EI)fN��\���u�5p�76���YݟyA��ES��.��7{��=�@<Z��#�+Y���N�tm�
�u��g���+���=�v�pm��P�Ο������K�̵�>#��;�#M#n75q��=����>"\���+���{q�����)��v��J����� .�ȝwq�����]l�������B�1
}q��"l����Ɵ~_�Ƚ��?<�0�}��(�ܳ�9y�s��үn½��_qŰ�g����N��-ؼ�ac�Ա���'&��ۼ��n� ���ꆇ���??�Ȅ�-�l�?��%|�gk���p����G�ˑ}>�h� q��3��:��O2�]߃rf���z��}�Ŏ{{q���a�3��M*�b|��2�����^��'�S�`��������KDn`��Æ[��!CPlĞ�b�����1�x;Z�6`g�KH��9�����[H'���̱l���cƣzpuԔ��D`�^L�2v��5ԣ�'���D!2j�h,\�/=��p�^,Z�r%V�Ze����vI�a�&���X�wC2�R��l���X1s,f��tr1�(mlD�0&)Fk��ȉ�<���o��M�Нo������*z��n�bd�q)[�$2�=D0�D܁���=$�|���˘&<.�<�8Tc�1Q�~?��n������n�K������H��׈�=��Z!��E�(W��ӵ]���%.�k�X�O�\�_\��������u���/�_S��p�;�k;k|*��Q#��'�fo_�f�DC}=6���%`���F$���������%�c磡C�bܸq�6aJJ��@q$�Mm-���CgW�}�R���>+o�[�B�ߵ�s���]Zέ��c���iA��k���������v�sH���wu���r�6�+���83`�U�4��L�v7�[.�=���Ϣ�����e�5T-[��F�J�q�{~�]�SYƻn��"`c����m����,w�"K�9h5RIn����V,�P��P�QxT���柟���x7|�]����N���>3'�Jx���R�����8�o����Z]�;m���������>؎�0�v8n��)<�<�对�y"���Y��w������p���2��S����=M�w�
����8���ȝ�<���?�A��b�De�N���(#>{	�3���L�&�YT&_D�:�чx�-����>��;�&N A��]�ƌ�qc�b�0vl-F�n5�3{�޽عy+�m|+�:Vg�_��齵Cf����&��������"�Vl߹���"�L�g
Z"��;o���"�[��2�=���.\�7?��X:w^��cY.��X�n�1����=��E�ZD( �� �Q]託��i���\a{L�^\H�.7P�����T�¼��.r����p�޼[z�(/;(�x�Rum����
R�X�|;w�Z�-4VoNLmy~by.ݳ��v�Ny��.J�=ʉ�P�\�c[͐����T�e��C�>|E��+���*�[���j��N�H�غe�Y�&����������a���GCC�5�_��Ig���c�b�ĉ�0����7[�z�������h�
��O�.�=b�|c%�^B	����Y'.-��h���IU��q�ܒ��ӵ�TӴ���q�X/1�����vII^�C�-+%�z��vq�����I۝5 ���S�w�l��1��'��t�M8�s�������BjJ.�B�{���<��G��C:��In��%g��i(�)-)��sO�D��?�� ������g%$H�).Jn9"�a�'��V������~�V��~�5�{�����ב�Ԏ�;��Ը�^l�݈���NMk��2v7��s��F�
ۇ����4�v"Ӭ۰�=}I����Y��g쥦�,Q�1q�P����X�oj"���}���
� �ǲI��ljGyy�22���4�ﰘspWM�\q����k�����(�0�J��t�u�V�́S��}��A�ePe��P>nl-J"�(�oX��1�{o��?�[7o���L���^/MUF�]mm-�?E�%(++Eqi	v�ك�w���Ad����֖Vl�h�p�z�j~��3fL����3�e1ƲRݨ���(rf�Ż�k��Z��x�h<��D8 �� bTU��[R�  ���������;1�'!���
��*�|i�Je� y2��뮻���!��ߋ�/Cu�`!�4�{3���bL1������0X��U)+Kg˵�� �R����S{
۵Bx��g�@��m���-n�r�ܟѣ/a��g4ή�>�~wM1J��8Cg�7CSW�{P������1���Zמ��>455Zo*3q6�^؍>s|g�p�ԩ�>a2��ˬ����	{,������$�x��h�&/C���'^�r���浜WݵB�81N�FP���.	�}�؅��]�c��C�]�_#��=Z��\ot�ڄ�q�F�n��E�H {Y��o���~�A����G}4�̙S���t7V�.���i��<���,������Bf?����Á�#��j�"
&r���/��7?f��3̵������G��Os�;���چm8�w��_�W�̄�l�5y�_�/������A��}Ҙ�_���-��sw�y��wq�ooÍ?�rܗ#x�k"˰���<�����s�}X���~��y������Ww>ܞ?�&����c1��"�~��Q<��C�=F��Fgq��_�3�E�Zc��"!�˹�S��Y�yI:�~�N���l�&Sv:���k�J�p1r�h�_L#�D�6d(��2U���vv�hjl¶�[��Hw� �Pl�ƍ�dî�#G�Ĥ����}c�Z�[��Mhj�kAd������V���"<���c�ڵ8��s���8�g���3�3�]��>C&rgϙ�VaL�ޗ�1����Hmj@�� ������E��p�1��#���m��D�]i�R���L&����/�믿�r$���E1z��{V]�!��|k��Țk��'���=��)nW�ԉ]ˉΕ��X{%��1��!|��Tˉ�P\�v��ԕkz���q��C��������׵(--��1��)����ض�?��ըB䆶�6���[��`�x���iӬ�{J����Չ�;w����m��!n���1�.)�v���y�vM��(i9G�-	��k���ō���~��m��s���|S����jjj𭳾�?]xzzz@����^\q����+���vTHG#S���l������9��Sq���}V�V��s,���s�Qь�1𜙈�s4��iGb��1��GWw~��Q3��r�������ܖy�e"w<��&|�¿���91����-�A���3.�+6�ʯ�m�v&�N���ڄ��z�?ϼ�N��Z���S0�&�5���&��g\t���I���(-)��g���}Ƅ�x���y��ͱ�?{	��_;_��´�w�O��{�A�c��R�67����w�g/c,�+�|'��U�v�ȝ�?�bpS���&����^x>� �pQ=��,_f��A��oj�hL�0e�l��$����FKK����ߏݻw[����1y�d̛5Ǻ\���Y.�o�lj�����F{[�p��m�1�QG�y����a{`c,+I���Wߡ�gȄ{��X-��8p������� 	��ˋ���qtH�X�0a{��Jpp/vE���:��l����y!�e����۸뮻@��}���}fNw���x�ε]�_�!�+������8Y���S{
۵Bx�7���e�v7NW'���{�֥rM9ΐϴ��a�9��Hi�zj7CSW�# �kl���L7�G�B_o:�;��G���^!W�<�5f�رÚl�{��30a�8k��֎��pi�n|�@<��<m>�qK3�)O:��'N�nJi^������	�|�4��:�v�|I�Htn�I��M���N��EȞ	�v�t��c�&�פy��}�õ]}1�Ą��_����Dxx饗��C�3��LV��3�rRuq���ƪ�.{��#{��s\����ݘ1b:6��� :�z�����d��i�����X��ﭼ�7�B>p؁���~�F��媿=��y�����?��5JA<�;���[��<��L�����TL��s;��+�zDƺ�q�O����=�G?�w�ll�݈���/d�[�������}�r\}������uaoS�;����k�=s��MK~l�o{Ad��Euh�̰����,��H0ƒ'�(�C��-ˉ�4�ϣ�ϩ���2�gfzp��W�H0d���a�G���A�FyY9Ə�q��X�X����K���Kd���
�z�}�f��"�ע�Y#�E�%v����M��L�"%**+#����?AOw7�p�4�~����Bii�����v�vq���=�7S7ƚY�D�X!����'����q��*n�AQ@`;0�N
����J��bv��Jm��O�2����]Ԙ�#=���1�j1g�\�sb��O�l'��.d����ѵ=eq�R�]ۥ��]�iyC�fo61�D�\�c���乢h�Ȣk��um�����q�P=�
��ￏu/�L����w�^k�1bWѵ�4e2�뱧�N:5qCݿqm7�Ӈ�>8���Svm�-'��n9G�-	����n��g'm{�ܥMJ N���S�.��
��X_a;(nc�v�������?��c�{����,]�C�Q��KcU���2^�U�}��X�!r��w��y�b�^ϲΰ���}��6l��Nf"�����m�<�f�OK~��3�\�M��ȫ�XpOcn�}fM����G43�����Ǳ��W@>���>�q�]��/���D��E��y ��6#W0�/;�G�N)&�߲;�\��[��3�]�;��+�Ĥс�;�K�����	���ܻz���ǡ�8ywW����?=r�g��W�ӛ$+����,�+�Ғ��v� "��7�Mu�{��G�na�X^�v�y/]��:�Я�h���_�5�p���Ň/�F=%"q�14q�L�0��?lokǦ�>�3o�"�a�[�l�&���;̜���
�E�m�lh�T�M��!X��<��S��/���5"ӱ��p]���5Ʋ�⻸g�K�3l�ߍ�#��:z�8�!�� �,�+�l�K7R9U����w`��ۡi��5P�d۽=[Bwy�?��<�<9�����j�lIT��%��ϵ]C���r�JYYZ�Rng�>ub�1�%5�q��qm�S{
�5�
�vSZg'.K����)���Ҝ����Ԥi�G��Ѳ���j�?`��i۰����
���A.uuuسg�Ր���oc���<~J�ˬ�hˎ����Cs>���J�	%��D������g3n �<�+�N���qm�+��<h�z�ӥ��{�&TV]o݅@sΆk{B"�hj�8�4q��ݵ/
8�4qb�џ��oێ�^&_Xغu+n��f�y晁�����;'j�n��4X��Ѿ~ΑA�Pe5RI�ڍV-u;0a�4lm��*"�hh��q?�}��8�Ғgq��ӎY�/-? 7?�*n{t�۲���(���[��_��B,�*|NA	��o�'�>��I�Ł�C/�����]���D��>}����E\�����ډl�d����/[��T`�m��ч���-8��kq�/O����/���-{���3/����7��э�?:�e�w�����N�4���!���p���3����/�80my��Χ�[A�gVu3�{K���8}�n�a���^\�������ޮ#��0#�5k֐x)d�p>Fצgd�(0S���Lǐ��V���m���O�� ���A�{ ��a��sQSS���^��4����t���c������A���l�2:4+}��#l����z"]�aƍ��>C��ԥ����$p ,�T���nk(���TE������X��ޮ{�P����L�	���l�իW�%�%8��PZV�-��E�"���p]��r���)nWꔠk�RM�� ���[e)"xC��w��\��;+~�;�[w�K��}���DEy��3�e������o��Gz��(l��w�yǚ#G�Ĭٳ1�f0����������)�!��rm��Q�Ը|sm��\SVPq�sz��54�X?ز �I	�)�u�|�(n����15�X�%lW��ow3�v�D���W�c�v�ܾD8`�O}�S�g�}�.8�T#S���j�\ܹgC��J��VVC�Ƒ!޳�3���ЋEû����B�����߹�oX��6��kG�ƣ���{�51:#尉��Ճ��^'�	-m<sn�XSU���g�r���(�����Ҵ�[���߾�xr�F&6>��wc5sr�v̈́�?8q���!xw��k��G�𷮹�z��-��7�w�%2�E�wv����>��Ӄ"ϸL�<xP����1�>�R��a��J��ĄQCQ;���ʻ�w�'�>"y�y�?�7��D,�;-�2��U?<��l�m؎L�^���ooÚ�|9e7�Ic����)kjl���V4D�6F�����ȹ����{{���Սp����~��+�JQ��F��aՕ�>>"���Ze��n}�����>S����n��+<D����N_�6V�+�g��l_%�̪U���2��g�>S1���� 
v=_;�m�X��Ptuv������������Gcc#���K��Cuu5�O��A3�QVV�{va���8� ����~hjh��M�A���;w��o����='-_D���+�c�ֺ�W3ۛ{A�/ԫ[�������� �V�T\CbPq` <��*�l9&�;�D�a������0��=G��e�v��>�?.��>��Ғ��ݬ3��~Y��0R�z�<9�����}/!I=���ڮ[1�����-�.���cWX+l�f����Ų]]]�uo�"L�.)����::�#S��eu56Li�����푸��N456i�}ut���<�{��(U���*tF���Ǟ@kk�5��y�Ɖ\��;;ߖ���|&�@+����C���lڴ������g���Q��"`��=���҈�5�� ^ �9��ݳW���uo*)a�s��C\���aod}�[N��rP�4U�h؝v��:�w��W��kU��8I��mؽs�&;CyK�v�ruҍݡƱ���n�����P��f��u�׋���m�mعc��=M��Rj�m|����>r~�weu��=�ݩ���|�����.�����D�r_���*���K�.:2���~ˑ�s���o�'����n�VLEc'u���u��7^�`�%�7�&��W��X#"�l��{[q��wa{�zd|�]|뢻��G'�3�0��i���;{,A?{	�H�-O����_�q���;G���/���^�����o|��~��6�^�HC�+�)_�9"�,ށ���`~��;����8�vow>C��gR��t���O:�y�7p���C���C� =�2s�t�5��}���&lۼO<�8���+\�n����#L�<�Z���blߵ������%���Ԍ��F����oǧ?�i̜93�D��,vc,��3�Z<�m��Ld�8�+E{�����q���oq�F � @����l"�b�E�U�9�����ɓ<�嵝�Mlǉ�7��:�dK��%Q�����;)�"	6�$z�������������������������~�6dddH�SsaP��7��i�T���`soקUTT��w�U�m�Ѧ��7��|u�+`@�O�<	#G�BwWW��R��
ٰ���� `�b��=��x���4�V?�/>A��S}J��BX�ݝ�����ZZ)�[,Z�����L�m�p{�����޿9\�
=�g�G<����\�Mk���;��==��W�<��qIȘ�='���cİ������hn;وȮ��M|`e�]�]e�]>xv{��J�ng�,6b���Ŧ��kܩ��۞�F�b��{�{�Ɖ��یx)�bf���]�����{ݷ�C�
�Ƶ]H2VI���++�p�����F(_�@",�fnhi�����D�R����V߀"�HQ���c�
kwI�K�{�����X=.�\�v�l�`Sȭ�|��ʵ�|;�/e���G8t�V�^=�U<��U��*++�i��?���'�^�ąAKcϧ�E��2�ca�������?�<Z:C�}~�1��ŝ��<Al>|	��d�;B�{��?߄+����G��M���#K-mS������K��;�Ǜ�ת��_��7��5L.���������@�=��B뽛HMM�O!���)��1�"�/�:�C�7��#��D�Ň��ۣ���z&�c�>3��D���23��6�U>�K���@���i��1{&j+>�Kks3��o�X�3j�KDj�3�8Ю�;�:���@բ%��^���\�f�ύS�����!���TU��$�lև`�1v�u��Zo��7�`�6��	��:xP�������c�NKG���5wj�>O�`�5��,�N���v`�������v��Y���E��#v�c�FD}��u�~��������(d_�2Ɗ�1�1ݍκ
d�OBsW��">��}�S�ڈ. ��_��" M�.ua���}P�V�op�Hs�Н=��Q���v
.�,_�;0�d$��8K��|8k��� �=}��|����+n��r��,�0�Jd/�c���ra�I}t��i,U��)TT���1y���P6�ӡ����!��'�onh���_��s�ȏG8vE�&�I=��'o��n�l~aa M�/�&�_��%/nnΝ���5�Ǎ+�+%CV�~_����!5Սi�� {D�::p��yܺqӿ.�G������FӨQ�t�y�v��eÆ������?[�6�/¨�\�{�U��bbm� ����{ܭ���S����X"R7
�=a�h����{ow�:cŔ�ӂ����kZ&��pߵ�$Bt�;��\�'O��aÇ��	۵�Iru�i>��>}��qص]Q�G�Y>�[__�LfΞ�_����d��g6�>`~>k��e{"9�!��Z}g��^W������ݮw,vͳc��+V8���M)^RR���Na{<�U���U�"Xe%`�ڧ}.�C_�8 � |g�_}Ъ�
���	�`����~��h)�����b^��]����]A��4�E�/l=����[�c�_�|3�k���|��6����������)�q����������?�����ę��z�𱲰=u)��=Ԭ�����+�s�L���|��-b�S�9�ivo�s�N9r$&"�HaO��*�����Y�U��+V�%�J�7&/��1Ҙ���v�S�\��o�3:��m+����P�����f�x�{v-M_����p��p��ܺuK]�b�c�L�Z����Փ�]���<vv�c���gBܼ�<KF5M~M~~>�-Y���L�ܩ���e�pP���<+���卵���}�����x��H������fw�������~�����ٳ�ڵkcއ����c�}��5�ZSl�¡��}3%׍��{HOO�,P�.\�ʢs{�E�����x�����?u�v��"9����V��KD�$x�߾�,�N.�@'��ۥ��F��¥�yė	���/'���g"��'Bw@�:ydR?S!�XM����ן�r����̵�@\9j},�ݟO1�i�v~/�Ǹ�QܮK����׎�<�|���aʄI��6�Ο;�{�� �E[[~�sj�����%KT�{cK��b!� ]K�?�e�t���	��l_��<|5��>!]��b�(���ZYKE��mR������ }� ��R�:�|���˷�5��'{5���p���9y��p�6mڄ'�|�A�x�xB��߷D�.wrOᖠ��������
���V,��j���nBvÞ�m<�se����z
����I4�?��?��wPy�	!�������o�u�D"w&����D���w���������r�����o<���n$���|�����~�|���1�8r����p��A�G�n�2um9�f�e0ƒ��M�!͇�[|$ʽ=V��v�&��/�& bu���[��U>+W["aQ�2�u��zI��#$���~��.�ʷ����gW�Lp��x��<�S'MƤ�	�xO׮����#�uf.�j�69��so�Lv;�=��*_+;��X�����'�ϓ&M§�[�=�
�ߺ�[��b�y����z{]��[;�L�[�qE�1g�|��gh�;���cg�v�mV>��i�ʕ�0��6�pqW{%}�2c,S�{�����p)c��	/$	�1Kr;�Q�2��F��U����(^\�}�,X��`0�������_���)av]�X���=^�.��+d�v�ې-��D�.#�w��K%(l��[�����w�K2�ORw%�h�C����=$u�	���g��X<N�d����  27v�P�_�Ż�K�򐺶����4����V�o.�d��۝����dg�NMvl�F�."�0���W?��՜y��FyU��t�����=�h�!F�Ǘ'�hݲ >xK0䉗k�T�-y��򅯿���Y ��(�"��v�9QM����#����$Ͳ���|B|��}��O�j�-/E�W��uTWV�����a��^x=��:��l}"�L��Od�I�U�����?�`pq��|n���.�����_�-y$"8z��������Q|~�\V��������v����Dh��?���Ϟ�>���	���o���Q�P�W�����?���4�w�Z�[5xy�)$�^���o~�׫��g3��Z?xq'��	��7����1V3,��3�
�o(�;D�������m�x����a�\�~Dr0y�4L�91Ta��.�3i�Qv{w&f@(1�a3���+L�6�^���N��p� ���̹�hlh@��� ��ŋ�q�F<��S�	��K�/d�;;��jB*��1�!�� eTf
��k�#n��� �G̘�ۍ��@�&���c鼠O۱c�?��T�>��(AΨQ&k���˅����ɒ�z�]�}�v�>��Y*l7��Lx-�����˅�<֮����ȵ]��c�n���o�h�PE�������yy(�/ �B=}�::� ���b���ôIS�k���rQ��	>��	��[��\L��[1���<���ۏU�v-�����i�x���.�g�K��&�NH�,l����k;���w� ?���S�Φ��o�����`���&�K�����U|�*(r7��vj_�ߍ�O�
�����[��1o�h|\K�*"9hn��w~��N^ŏ��2��s������?{{O�<��u�����`"�dvr�����]TЬ	c���hn��s�K����g���'��6��k�jr���tu��/�{3��sA8���;�0�sHc,S�w�s;����Pt��xϭ�%��QWW��^{Dr02'�K�� �"ƍ��������chooA$�<�VvM]2331���\^U�+���>�	b�����u�hnj�l�����ǃ>��}K����l����ylJ���1�n�A�A�����y��v��/H�O/�2P�|�*�ta�qB�)�y����n��W����$aڬ�4m�����v�0�DH.1�5�]ShJdA��
�QP䬭��(_"0����v�A�:*�D]:'l��R���k�"pmαx�=�}��v]�>�6T���O��|*b�ظ�+���q�����=}���ܼv���{�X����`KAA,Z���lܮ�@k[�(v�a>{|y���a�(�H.O<]������D߶�1Z�vA�Ο-Ͳk;�|jJT�L�,����	�%?#�N�Y>+�v����B|�k_�+/�����7��g?�Y�?~H����b���`PJ�˝�mOc�*���

�-�����#��qm:"�xs�9��^�_���1k�v��?��P�L�D�|p������X�����a��2�e牫���_������7��BZ*�JI���q��m<�?�_��Ӹo�$7�����ĥ[w@�3XR�Fks�32C
�������f��r��;L1��}�@P�.�/.�i�!t�v?�楗^B}}=�ÌWV�_����P!;+��C�;W>��}��� �BGG�9�~�0q"�_�=}�8s�<ZZ[ACw��k�`����%C�SSS��_�>�lT}x���hc,���P�7�"�9�A��A�;p�Vy�#��]��)e*>0%����E�8/�$K��~�|�M\�v��ۓ���QX�l�dM���r���AA��7�k���}��� '�����k	um��G�W�O(���µ]���=��A\����K��z������)���҂㇏����L�F`Ͷ�sa鲥�5u:�5֋�6?X�D�)
�%e� ި��%̵]"��$�GV鶰,ngI����xq{��5b�<�|��Ua���*�KKp����!gÞ�/������>�6�]��*5Ű^�T�)X��S�ۺno����}�����Mk��Fa�4T�� Z,��6��)�5Y{/n�H�ؑ�Ă��s��o=�ov9RB\�N�9!��˻��&�C����/����O��>��z`<~��G	-���ǎ2OwOZm��%& ��^�o����礶�u���K���������z|���Iq��t����>H���`�N�uQN#�05��ݩ����b&x7�����'�'����vh1c��dro�~nܸ�6�H��Z���`�ݧgϘ�����؈c�F~�dn���Kzz:.^�ޯ+k�q��U2u#=#G�`��R=p��y��W�裏���hH���TQ���fc,���e�X�d��@H�>Y=х��.�[��s�\���b0E�/�k�!����8-��}3����_~�^�� &�\�~�:�'z�vN�n��X������]�k�v��vH*܁�8\����ܲ�]1�ת�=P'����!�G�O�D��mM>�յ]~q{aA�

��vl݆��~D2�\ݏ>�~�>cF���Ģ	�]Yaȗ�v��[�{ty�u��k;�ñt��pm���F1:�SX��)䋽�]�ϣ������k��n]�n�����O����(���|��x�'0o�<
V!x�V���ԃb�UZ�S���Yrd`"�^%�c{�^�Y��Ld���u�[4�4��C�wb(���oC��w���M�Z��l?	;�����=�o�;����()��d�����:�����@����ϣ������=�4"���:��O�E�c�����?|���ͦ������C��d����_���S
s��l@�W��5[��濼���^����O�pt��م�7��K1�-'0"3]�j��kUu��ߢ�N�R4�����:��D�.��ٞ�����`<Ÿ(��+O2��t?���/U�ٴ�4�f��b���<�.���|��6?��ΜA$]]]W��EEx`�Z4�����b03a�$ܭ���+4K��ь����!�F�X�c�rm����1��d��$H�>��C��< ҉A7͠��H�Sf�*��bD�-�>�c���o~�ܽ{��)�o���K�޵][��+� �tm�nle�vU�l&����	�?.�G�.
�9=#45�Dr'�v1ݪ�=&��|�$_�\۹�R_S0}�4�de���r�ܶ1)�z7o���#ǰd�Rd������T��C��M���=.��ϣ�)��x��C�fq[X�C�̊�k{0yyѹ/M<��	�}k�x4���{��v]u�y��R������_~���N΅M�����?��e�y������PdmH^�\R�a���`�*��B��j�F�{:i�NU<�������KX�`�asm��;�۽g��p������b�K���{�ǌ4�?r����7��i�t�Ld��߼�GJf�ϾxM��D�|t���>U�K����. #͍����w���k����u[�����g����ϞT���0����Vձ|(Q^ۨ�K����0oJA ���_�����8���o��?�����gJg�I\.��>7�_wƹ,�g����{N��G�Y,�UdX��<���l����p6%���'o'�֋���jz�i���M�o�m;}_a�vk"����ɓ'�k�.�'wL�.^���>�������p��1455� �꒕��qc�b��8y�4��i�#bp��d��Յp6�1����#�#c��c�u3?��?�(XQЇ�i��� �� c��T�46 #C��.�XCM3ȋ� �T�.� ,z�*j�e`���
o��&�3�x6
��Ңwm7���K��ǵ]"U���%K�Q��x~d�҂Չwm���XL���r�JrC>�$� ��1�k��p�`u<�܆Ӯ݃}�X�~��b�������xu5b(��mߺM\���"gTʫ*����� ���O�	�=b��\m���u�z���D�����DD��n.l7�v��HωGH�.�I�eq�\@�������/�$�uq����qEޘ<|�_���
��9p� �9��+W�&H�?Xe���`���tc�
)\�t�f"w5�D����������`��/��U|���X<�	�\�U�7v��E�����N^��k�{��xd�����������32b����j�$A���{����U�a� ��o��U�e�{�syy�)ܪm��|6#GY�=|��E�9u�m���E��\��
s���^��}�0f$��:�ܦc�r�Y�%u����}S�/�5N���/n;��^z��l������X�h�.����3Pq�I���(�<��+�j�T�Z5�2�ۃ}�b�a�i[NH�ԉtmV�dro��_�}��/~��>�w:���\w���&��F��ј;c6z��������AFZZZPq�G��E��3z�^��w� �}�t��޴�g�F8�x�����rc��˥cU!�=]�C��)	 �� c����Xwo7��SR$��������|K����N4YM�~^z�%��(PǓ�;
�hѹ����6�]���N�-����u���ks�vQ�������-���H�G�W�Z��0ߨ�ET���C�1�c�iV]ۇefbެb4����ӧ��:��B��v�ڥN�[��ESǣ�n-Ztׄx?���C�֍�v�N���˵]�BrѺUq;$�,�k���|J�]�%�: a�o��ඞOvB��E����a�iy.^�Uk����πp.����_�%%%��@KJ�*�o�d"r7wc3ݠ_�n�B(`ev�x������o��T�GwO^�}F]�Ρ�ԅ �2�_R"4�n���^�"��O/%���֣��1t`��{O_S�������GjF�Խ=lߡˬ�P��l�2/P�C�W�fǾw�ޭ:��g٪Rd�A&F��C��Gc}�ۏ��~�P���8zT}�3w�ŵ[7p��M�`aD����
� ��9x� >�U�V���7T��y9��[3ƚ���7h0�S �� b�pZ�j���jY��r��Tza��yAV�[ě��D��֡����>g�DF+֮Q��d$�k�o��k;?�D�{�]�a.��"�%q�dP�~[E��>M,'�$7��H�I]��O����q�u������?{�[۰w�nܼy'NAu��ȁ��#˖-��)�PU[���V㵪��nE�܊ܵ]E7Ї�[��ĵ]��>�F�4I.�̵���c|\�u}Zt�L�,���z�ָ��|��y�~�ш��|�I\�Z�� ��޻w/z�!�Jv��I\��X����*ƀ�&r�̑������T59�AA1xpy�Ri�����.��=Tߡ�oȷ����<�����;���/�v�~f�-f}&�d��o�͞������7�Į�4ؕ��g���/�˴�����5�t����&`ʌi�WC�8��������$�˴}��G�ͮ�� �	���}�S"
R�������W��漠wn������[|8!��H��鼜ϒ%���������ȥ��rm���B�(c����9ѵ"��SXBx� �Ӌ�����C����E�\^�0^�gb\�e�T���GH��ڞ���y3g�|�w�:�� ��>~�8N�8��K�B���*�wt��:�^)T����1�Qt1�E�0qm�vF!n��%sm%nx>���vs�QU^��[#6�����G!X7�g��r��`>�ݽ���^��^����տ#��x�;t����0�3M\����*N9�k��{۵��SY�Ϯ~�������a-8�AAA��w�������0�?��v��0�k;'n7.|�=H���E��-[���ŋ �ͨѹ��x!b00s�L�8	�=��'O���999 �VV�.��������nC>����D�d>ܾ���ΩS����I��`c,���ڌ�8[C�XN�����n��~����.h�(.� Y�
�EA$8A�m�>��c��A�����)��%!����/�Doѵ]-�#�{���n���ź+�W�*�	�e�p�w]��z��IZl]ە@5![ˉ�e�7�l<}-��RQ<s6��{���>BGG�{V�:y
gϜ����0{��WU���w)�\�RخO�u�zL\۹�,l�p���񣜴��]����g�fY�.�g"���w���[�G/��1|8��������\.]���[����=��}�i�! lS��I���c�����t������g6ژ�Sp���d&� � bp0!�m.�i��l0�6�8`��O���Y"n7������4M����/��2g�Nu��U�o� ����&cƔi�x�cl;�A�S]U�.�&M§�[����q��5D����'���}}} ��/�K�[�iii�w2Ʋn�%ӷFl�%���c�ц�Ha?$p$����܉�����9q�4��P������'	�����_��4Έ�l,)-7�W���3qQ���xѷB���e�vY�|Zl�b{M�m�k@$��ω��t��Z�;׵]�}b\�� w'T���O�wc��Ӯx_�\�3s�S�8|����AD�F��#Gq��	u
�YS��Bw�,�iq��h]�`-�?�"y��ۚ��%�)׻��uH�Y�vm�ϱ��{�v}]%k,�5y��XK\�z>��	Ο9¹0��~Xm�1�┐��oo�5��U27��x�_h���v�Q�J��µ�Y�mE��@AA��d���p��i>��C,�}�f��C���ͱ�&Q�Yy6l��7@8�ťˑ���HV�L���i3p���ؾe+��έ[��eʔ)����e�v���Dr�������� �KYY�j���㏇�_\}��1�2�il �X|���n5F���v2Ʋ�ƻ�aѵ]V�B	��`�4���=�/@�n�<NO�~�;�����p.�w�b�j��o�:Y�N{lUH���%����[��[�R��.VS�򺛊��:���a]Hn&n7�cE�����˄��r�JrC>�$_D��2��(Z��#�9��P��Aa���;�\ձ��#h�i�"&0���C���ѫV����B�WV��G���!^ky�|f��X����B�"�ܵ�w�t�k;�ٶ��'V��r�
�#�+}7auI����eܺq�M� �	����{�җ�dk��,-^��xQ�)>�_� sd���)��z��̉0l��.e,�<!/j� � � �S:��u)����Rhq�Q<R�-��3�Pt��d1��Eymmmx����E�2i�L�:��L�03&Oŭ7�e�f1p؀4�L�6�{ ��]Ey�mD�1m�L�Vՠ�v��y�2Ɗ�1�|�2�"i7�����6�d�C�A��l7Z�� =ݚ{�!H�2�1�"���휸ݸ���I�x��g��N8���`T��w��V�ߘ��Z�+~��k���~�:���V�����u@�/���ta�T/
�4q� WO���;�x��i�X'	sm��! nl8���S�"od:��&{����o�>�U:֭_��a����Њ@�.�!(n�%�H\�%w]i�"ӗF(n7�y��C^+�v���{����ػ���)j������Z"�2|�|�o�����p&�~U���琕�H�;X�� V����Bw�w1h%�nP��q��.��A�r�{WW'J�Rq�6��EAAD��N����:ҙ� m���L�Yt��`"�El3�8��*V�������\�g���� �d�pl��*��7�k�;�_��.�s�����ŏq��]D2�l�
��`3:�;@8���r�����l���<-^���1�g�1VjG���)�		�%��誋̹]&n7��%�Ԃ0�ۍ��z������}����	���Ɍ��Ys��u�:��ت�\�E/J���<f�v~[_�@\�%�A��ZZwSq;_��\���k}�`5ż��Q��,D�lh(�|>�x���|@��O�0����[P�����3q��y�<tAğ��.�ؾ�F�ªի��׃�u�L��V��rm�܈���vA`nL���o���G&l�t��@d�v���E���s����1pm�y0m��}`=>ܳ�3�s��z�-<��3�V�`���]��Tƴ�jS(`��x7��`� � � �����i�c��D����B���?T��!�W�XųOO��Z������p.췺|�
�SI>A$ÆÊ%��\߀��w�G.]��O.}���c���8x�:;A$l���W�Ý{@8���G%c�c����l�_��ڱt��*{@��В�TՅ�ֲ�B -���l��pn������ro�W��`�u�|�
��OO�]�%Jt��\gYl���ĵ��R"�6�K���(:M�nȫ*7��3{A�D��.w�W�k��>�O�������뵥���_\��������to!hhh��M�0s�,,^���5hmkU�yL�Ӳ����KH�k��B>�Ԕ��p�vm���Ks7vc�Y]��!B�ɵ=�5������K�����3aS��_@vv��ݩ������f"w��]�� �vPk��E�j��E���h�AAAD22Vi@��m�Kߎ��w(k�	�7�6|�a<S3�ЯhV/�oXWW¹̞7y�� �d��w�.X�w:�݇�]D"`��sgϩB�e%���=u��� ��_X��g��+ ��ݻw���o�w�w(*��XVL��n7&�5�2A�	ܓ�U��ֹ0D�&�/�J���T����*�o2�%�.Nvo߳gN�>¹L�9Y�Y�f�/4�q���\�e"k-�~[3q��]�C��T�.�I.���Wz> ��µ]Z��v1��'k��>���n���F2�����;s�eN�A�˕˗q�����b���v�8V���(<7�G#n�l+Л	֣qmW˒
�c��$�ĵ]��Do�	������=��<nw*���o�?�	X
��f��drq�E�^į'��4��V2'��������X�xi^*�@AA�tL�q���Խ�l௹1��H ��d��0��3��8�o0Z���ذa�=r$��A$3�M��	�q��a՜� ����ݍCDNN\�5U�t�DÄ�Y�t1��Ԣ��:@��믿�'�|R��0�+�1��g7c��ZfMCuc�	ܓ�|ԣ�saH1	T�#T\:q{�i��(���`Uh�����h�ÄC̅�p.�y�QP4� ����L\T%��������PBtױ:y�-e���g��.y[�K���=$�vUyi�k�c������Q$e��L]�����8���]۵X򔉓0nl�:�zru!G���G���ӧ�z�dd�����>��$6�C��s�`�_ [�=K�"��+FQ} �xێ�k;W� n��.�Lخ�9��c0�#�=A��f{��������#��,�n��)ʟz�!�
&�ި$"wM�n�������w��.���B������
�)��C�B� � �H2���A���{�m$�K�7��"w��1�P�k�����HD�T�oy��E��d���a�칸^V�m[�� �ill���;0i�$<��~��p��o�p0��d�J�ٲ���
sq�w�ˏUc,m�gK�X)�����,ۇZ@�	ܓ�i�n47�I]Rn���ǻ��+����]��!
�<g�b������̙3 �Izz:f�-&h�A3gT^T(|�BA_^��:�/kБщ۹􁺶+!�n*n��k;$�C��k����;/�O�k�$���0��Fdaa�\\�pg�� A΅ͪ�g�n���㾵kQ�Ԁ����z����v.ђh[����bw��&l����Bt�$-�7&�v]f��ٶ����ۍ�ʵ]�j1�髩ٻ���t�o<� .�?��@8�z��w�j��ؤ�׮}[3�+�̍��R���lf�~��u�>�#�q�3q�xWW'V��ay/� � � ��47��X%�q�L��3B�ۃ}����Pm2��ݸc�z��_���{��{��)�4#Ff� �Jff&�/\���&�ٹ+�ށ ��s��-���c��%X<w=�ήN�������sq��y΄���O��Xc�I]�����-���S
�K�Bl��I���Nt��S))a�U)~��@�ʕ�]����S��� ��;�`��?���Ԩt0KV� --��/�Z͊k��R����Pΰ^'l��[J�إ�v��Zs�5�K���=$�QW����!��M�����.�'=0���E�v��.��M~J`|>��9�̜�t�[u]�룩m"Y�s�6��6,X��g�V�mt�#�ik��"�<!���$ك@���|>����O�k{�"x��v��]ۣ�`]���]�r�M���vr���?�Ia�����\����[����??Do/	v�V=������V��`����Py�˰�RGp�^��9��J��>� � � �H�Lp���7`����,�Cti���>�C,I!�@�7��b.�X��D���|��7ɽ�����#���T�[���G��G���� �{�:qX�z���Å˟� ���VU���=΃c���{�ַ�R{��$W�`�4Q���1�oq���f�}!���~Cf�UZ��A2Ʋ�')�.ݍ��\D�vލA�j0d��T�P8I�� so?u�gR4y"�O�����������8�Y�v���,�Nt.�˫$<�<��O�ĵ]�ˏSVnT��]w�ssFaެb=rwjkADrr��9\�z>��:ۍ+-��KEےm�qm��Fat4�u�>�m�yC
�u����#I�ۍ�v~�yyc���㽷��<�`����o~s����Py�#MB�2�����.�v�>M�������i�i�!AAA����:t�ܦ3>��~�3>���Ӻ��j��a�C���q�0=�fXx뭷@8���T�ܷ���������ƪe%�p�<�ܦ�	"�������{0�����!:y�m� '��뗭^�]����Cy���Uw2Ɗ�K0�һ�{ۿ}C,��V�o�FaJ��>4���=IY]�BoS�%�k]���]?� ��`U�nħR��Ty<�4`�.�3IKO�⒒`�U* ���M\�Ec֠��߫�=�ϸ�����E��Z*����a�Bµݰ_]����qzd�$�#6��&�u�\π\�ŀW�+����s��m�n��G"b`ttt`�ƍ�2u*�F�Fzj:�{����8½]M�=Q�n*l�P��/D��<�1"�)n�۵=Z(�{�哽���!B�,X�@oR�uq���V�Y�sg��z�5΃�łUYY�����|N	8E�&��h�Sd�`pJ��td`���Y�J�^hlG��htn5� � � ��L�FksC���%�+��{x3,��v�;��%}����TN�ӋW����F���e���6|8	�	G���-FzJ*vl݆��~��TVT���
�J�ctv��8�pY�٘�p>Ο:�y�1V`MXc,��P6��K����#���f��-�P�5�-�~�hH����)��\t#HB�0�����]t`����k�!�����i��4zک,)]���t�Z���Ep����µݤ���U�D,:L^��\ص������j�H��:�H�ڎ`Q!��Qsc��Zrm���--�/���Sp`�~
p� ���U���by�r������ڿf��*Ҥ�	s�(���=��`ސ�v]Fö�|�\ۅ<�|\���!M��״�S:�N��t����em�/~�+�ɿ���4���`S���;�`U��ݭ��/��LD��E�� ��@�"���y<-5p)c����AAA$�Ey=�g>�W�w(k3�	d���c��oێ<ɘf����6l �L��b��� '1&w4�-\�ǎ�qB� �6H�ؑ�HOOǂ9s�����M8��s�QUQ��;��t"d���	o�e���h�H��3��O�n��?@|�~lj�`H���f�F�\$��.��L(`X�
�E�􁪡����1�vr_v&�E�1a�$�D�m��-lε:��a���Q����e4��Ʋ͎3>���9�����^ʱ���+͐&�� z�v.��v��d�"�VW���A^X�j��m�0aV�^��;5�û�ޮ&��۵�5|��\�u�yq����`����K�2�����p!%��>i^�X�\p?fL>���`��A8�z��1b���@�N���G�~!�o+�wi��_*�0����}yu3��׳�d�KŉJBAA�sq� }M5 ��@^i[�\��"�4��v�g	N��3K���o�[��׃p.�O����=�t�2�vucۖ��9 �AHCC*++�?���g��#���A�{o_��;7mE?�&��\ܿ�o$M_aB�� mT�K�Whj$�kO��ZZk�w��>��0H���,ۏ޺`'��T���2�v+.�`�4P5t\��:�cǎ�p�iiX��DP{��jɵ=�?�vA�.���9��*���@!\�����|V]�5q����$�XssFa鼅�p�>Q�JĠ���ۨz�m���~�����j�\��4�ʟf�G.X7������d�3��vq[�$-(n7B���=Ξ9�۷�A8�z����կ~5�A��m +�����q;�'
1|�b�Jtd���'N�h�	d� � � ©,����.ddd�S���?�c���!���5��,-N�k477��7��L�/Y�~L�����q(�>GFKف�`��+�>u���XW�
e�7Q^qa7Y#�Q�`.�>�y���+��;c!l�ahc,En��}���%���XT����= 	ܓw�x�iLSڈ�8�0���]�o�A#���e6,ӐpI�r~�*e��k�O�΋��ڮ+Ǫ�]�wK���vC�%�z�8]�����D&�W�k;L�)����^[<}�\���۶� ��saؽkƏ�5k�Cyu%����qmW��{9����&���u�d[k�v-_���H��d�3HO(�ľ�Ƶ�b^]��|L����~��Sg �k_|�_P�-e8�Q!�i�����~4���M9h\�-��R(k?Tz1��sk]-FeNAC]+AAA8�"w3��n���C����X��?�T��� ��&����<�DRg��ΜZ	�;&�f� A���.�3�2ұs�1t`���ڍ�`M�J:~��iۙ5�U��PG392�
|���g�e�m̷���i��pi 	ܓ�Ņ�hom�0H:��S��ȅA�Qsw��c�v��y|��G �G��BL�:9�]�K�r~tB�D��C���k�(����I^@�ڮ��k��H�ٍi�pmgI#G�`��blݲ�UU���AC6��;oo��~}#�q��^��dQܮ�	�O�����>�u+��y*l�ok͍�j��`4��������jM��ྠ� ��ضygQQQ�-�w�'�x���Ĥ��h�� �'D[5���2���I�*%��r��������~AAA�cTf
Z�� 5-U:����p����]Z�~@�﫾������+���6l �<�o�d�J�~�����\̘0�.\Tg$bhr��9dee�����3�[wa���ؽi�p l ��6�R��=c,��=�1���0\���;lk����h�r΀���1'lH{�K:B$N�\��`�n��M���qo'��������R�tWn�@2����9 ��ӄ�~Kq�_�pI|9F��_"l*�/W�2Z�v�X_f�8=jrt���O�|�E�R�����wmg�3�NG����y�F5�M������͛1w�<u�YQX��"O�˺G�g&l��k���$Ͳ�]k������Ͽ7�y��}0����{�~�>y�5� ��k����{,���@R����wQ�z1�PfV�vw׋܍�7��2גAAA8����z��Zǻ�)��1�����=�)����x�l����x�}���s��1g�|���A���������<r�H1tiii���[Q��S&NƱ�'@v12'�����s�p�o��V����<�۷g�1�L��c��f��z�;?���=V�K��} 	ܓ��i
�j�v>H%��i�1`&8�waЂUZ$J��ȅ!NRݸq����)������;UF��/W�{5������ⶮ�N���:���!h�f=�bf!U�s����y��+G�)���Z���e����._ՕI����ȮI�n�z�xKs�wi���2nb{}}����㧡�W/^
d�����K6f`B�����~q�:����W}�ioo��z���]S�655��͛����ݭ7���soױ3�<�������.v`米�\kk�z���k�NL�6]��o�D��5hjl�_T|X����D�ht޾U����o��ʵ} u��>盽Ϛ���ЋDD��[����}�;���7�:Uܾ�=�F���9s��Ҋha���h�5?��o�����~<��pjp)�4� ~Ќ�;��.f�
R����Li-��5&����	� � � � ��.�Y�!o�e���o��4��v�_����x��> row&#G�`Ɯ� �����}�+��s����+#bh��GAaa!Y� =����/����媶�p���:}�Q2Ɗ��0��d�g�Qf>����gZ��(H��D�,r��ރ�4y�{��z��=���sa��D��7��8L��a㋩ݎ��*?'w�.���M�\�����ѣ%��&��H\ۅ-}�n^)Ô�Ӎ�T�b�������#pm�'2q��Y3��HC'|}$N�fy�\�YBխ��?��c��L��zB�O�||�Z�¥���'_��9s��]���s�k{Ѹ��_�}{� 77W]L��Į�������rL�8v����'O�����F�ߜ{\W�<v�˿{�.�6��`���c���SũEEEa�vz�V�Z���
p��RM�ֵ���S�9{&��Ͻ��EwwF���L�~��uƆgĮ��Me�~Y��	�++*1�!_"\ۙ�}��حmm��;p���{�y��ڈ�����:~�(���۲����q`��߾�꫸���uלSI�[��K�78����N����b"��E�����Ơ�j�������t���AAA8���n��4###Cp�sE�w��l��uq{����B�	��X�m߾������v'ۇ]��4��Gf��0q"ʯݐ�okiEKSܩ��&��1�5[�fq����4��<�D�?zT.��x���͵��K�m644��4��|�g�4v�i��~����3�rV�]�;���ifx��Xݎ;�>��[[P����P������T�]���R~2��	�'��{S$��;����<�8��6�����
8p �ׯ����d�e����3���&�Ҳ�Қ�1-w4�Փ1V" �{1������;1��L��N����O��6m�,�osɊU�.<��d���L@&s{���ԯ3���	*�%�Ac<�t+��>5�Dh*$�i"n7��s� :���Mq���Vw�7a��?��瓈��`1�1��Iqa��E�}�&v��$��{�9t�*�_}�ܮ�R�\$�,EģO3�{�/���Wo1M,#�1��ݷƚ�=�|V�޺�<o��V�������{���p��y�f!�9sFh���:&�{�4�����KQ�>h%�vP��nɍA��94�4V#5e<z��AAA���Dg�[�p��
S�s��� �1�T������3;�Jc��z�~�8C�8��n��=^�O�5��3]_[Y������D�Dg�gL��l6�5����h�-��y�(��{W.]��ڻ�t�����3���ȑ�8es&�����V�ف������9ոq�l)����.��ܳ���3fL���w��K�b��I�{��*���~�3�d�!6��$�g3?�߸U��>�w���<���~��P��c����+�`ݺ�ɜ��
�j��ۧ����PhCs�� ���ݸVO�X���I¤Qn�6�#==���nű�X�F�D&n�[=��������r�3y�<Nx���)�=q�\�9�z��X�D`�龅]*�D���bLԥs�v��㔉����cހ�\vi��ۅ㑉�}*���2M�|�Q�"x��S�-��m.�8x@��G�K�9�,���{<�Au�����~m]hni�-���
u��N���h]ۥi����NQ}�U�j�/��v �jM�n�������ǟ~o����~+l�(&pק%C�i�if��N���v~@w�@�U7���N����AAA�M�KAwc�|��žC3w�8@�_���~5�L�-���E��δ������� �EFf&�-Y�H4cF�a���8��C�g�$"����eTUV����ȩhhjA$��%KQ[U��8B8�ӧO�ĉX�|�c��`�e6[Y8��@{��kzݾ�Z���y�?10H��$,݋�:]P*Dp�J��̉!.�$D�JcS'���{ �R�_��Dܮ`K~�qrm��A|-�[��Na-���]����]�%�Y^��H�k�pm�y�ߍ�vݱI��Ӯ��� �ǍǖM�b2z� ��s������j�j�E��Z�z���%I���桄�j�GL���2���ֈ�h���Cɵ=��k�(/]��G��ڕ� �Ç~��/bΜ9Ip�E�Q�΋��-fA*��g�C��f�AAA�ݬ.b3M��΀�����͍���ji�~B
d��x���~Cso'����K���
�H$�3faTV6�o��=� B�钶mي+W���W��� Ezz�:H���c ��f������������\�.���ٞ��nf��|\*�T�7K�P��IBJ�]�&��Q�n����T���
��B�mذ ����epkA*7s���#{ ��vA���Z�ih����vIݣum���`]�ײ�}���@�>_p���>\�(�7�$����\80q�@(�v�iάY�i�P�A������<y2V�Y�k�7}�$��u���|r�k����5�_�/_�I>������i�{?�;O�?~�o4h�Ah�����4������~��+�w��]����	�].�Ck}-r2������ � � �%/��n����)�����b}���/�HD�]�ģNgΜ��#G@8���0y"Q��a�e��s��AD����Çav�l�[�9Dg��1e�tܾqwjjA8��{��ҥK(..4"v�iF�����Bd�������R��f�I_H����FG{+�32MU�L5ȏH��Z1Tm���n��� �E^~>�&M�}�\�}zf�]�_�lTm��
�u�"qm7���#K�ב������-��k����r�:Q���������]۽N�%K���Ө��AD<�y�&������|w��3�.(n�!�4E�����O�f���{�m�H�v}M���g��ĵ=q{l�o-���Xǌ�Ǻ�Ǟ��@8�;v�;������ޗ�(�N?�����V)-����]?���G��B��� � � �6Fe����RS�B��[�7�������/�^�$ 2� ����/uz���Il�0�oq�rD��H���Ukp����׃ "�|r�����u`����>C��'�J�aצ�����4c�������#b��1���=E���$��@ߡ?�����&���ڃ��I���.t�����*E�2so���߅�N�����q��m΁����,��ٿpm�8���wm���q���Ţc�ڮ�3J�����9��#�Ӎ	�m���\�M>	'^	Vǣ�m8�
Ffgc��b�ٵ��� ��'l��o���yX�n���	��Y�^]#����,�ڵ=�zE ��k�l��z '�CsS3g��Յw�y���w#N�`L~�`A*�~��D�M?�;����r�6��`����ټ�@AAa%����+!�ۭ�bE��]��=\o^_����fR�\	g1k�1���Â�s�k�N��� "444`��]Xw�z\��	�6�sFb�외z�΁c=��(,,�z_N�So��~
c̱,c�wpWB��9w�Ѕ}�zA��;����m���B�a��~$�o��26��Ȳ�i��{��Y�(���#�ߴ���xKP]C&lק�E��nاt�M�k;/$GB]�E�;`��n̄�\ۃ�����w#C�+�<a�rr�y�&rc!"a��۶nò��1y�ܮ�����z�x�
��|��O�f��鶃׵]��t���f��|rzz}��x�A8����<���|�j'�dt��"bB�4q�<X�;1(�*]��d�\�Y9�n�AAA�d�5�C20W�X5��-���u}���ZbE�8��/Vi6l@o/��İ��1kn1",�7nO
�n�� �xÄ�l0Ͳeː7:�/] Aě9���-t�w�p���x��w�G�G��+LL��Q���3�c��!ۺ��o�+��{^
3�"~����,�Fwk���	"�
A��봗�D1���U��
�$`�C(�-�ĉ8s�琑��}����.�A�@[�݊�vٶ����������Q_m(�/DV)-��k�I^K��(]�ż&�<�|�pm�pi��d���}�i��-�� ��U�}|'� ����㨮����vu%����tc���$-J�vY��|�qm7����<a���&N���!�-X�G�Ƶ�2΀Mm�e�|�_t\*�ei�Q�7-`�}6����~]�"P�:1D�.,��AAA	�0+-�u� u���P�wy�v����B��=`��`\G�o(�?tj�_,Қ���y�f�bQ�R��$� ��G�)Y�[�n�֭[ �H$L�4e�<�v=�<��>2c!�Gjj*�.Z����pl��o~�៵h����iA�?}�>����2w��tHM.7����FeNECG?��@�;�31��.�(�S/H+����a��d	DE[>sM$�fg�`�b�ݩ��o���BP5�/kU����ص]1�D���z�u ]^�ŵ]�7�`�����vC>Swx;\۵<BZ8�vv�,]�gN�DMM� 줲��>؈G{Uwj���T֠SG*s�0+���۵=�ےk{D"z]��������/<����O�Yg���o�駟���������ZV��$�̂mU�J��n^��$.�������_�{꽥� � � "�,ۏ�:]Ǻـݐ}��6��s� r�(��͈W���B��7����s�/,��	E �x2|�0�[����C[[� ��ƍ������PE�]� �x1y�T�,��{w�p��߾};�z�)�	���W)1���C���������ٟ��]���Bۯ��$pw0�n��� �`�5q�1 ֽ="�&Ó,��pTTT`׮] �Cn�hL�2% (7���=��Y'h6�KU<bz(�v�X^�.��È��b��.�ˋ�aP�&l7n�H�D�Ll� �v���ŐU_���4�,Z��{����,:	�p,`�����㏣������
��v+�vc>���\ۍ�����s)��[���[�ApA������;v,V޷� ������GaݺuI+b�4���B� ��o����e��pmg��-l��؀)��p����'� � "��uԡ�dj����B{�Z�ڦB��P3��	
���x�/��������ouq�2D<�;K�������1� �inn��m���C���3�oh AċE%K�{�v2�u6l�O<�����Kop�����Xs,����9��)���K�AM���.����7D| ���)�B_s��P��.sq{�O��nezAх!<��
�ƂT��� ��=.YQ���=2I��k���a�w��b�mF�/QShG�ڮ�7�B�(]�un�>�˫ ����+�ε]_a�����o��������9رu]�A8���wՀ���l457��Z���t� n��]ۣ���A�e�Ć�Y]"��E��ȇ�k�,�C?�S�O����3x�{�3����b�2���*+K�`�b�2L9�sF�?�7��� � � �2-׍֖fddd����/������Z?���e��ϲ��ݫ:��az�,d�$Q	?&M���c�c׎�$�#�1�>Ý�w`՚�(����JD<���Ŕ�p�Jgp��%>|�W�vP�^|�7��ͱB���K��6��̌��Q42Md�H��`ƺZ��rK;�C_\���Aޱ/����H�D�CɅ���]�f�p��OC����tm��D���)��R�9/�W�A����!/X7�S&�WT��KC\�=��uTI1$j��g�1�T0[6m� A��ݟv�܅+W �`,���	n��5sa�>M��]�%"x�h���/76��Q;�'�k��,9�6���g��[@8����˘5kV������1���Bwq�A޽P	��9#���zK� � � �D1?�]u.i�z$�X�@`����~	�dcoE����>�1�8���L/����f��I��?A��`�$|�%˖"k�\�r�.^��7��C&���w�Q�N��ބKb����+ |7�*��B���ںE�}�hH��P��S��xGuo�M�n�� t҇R�tr��t�v��_��i�&ܻw�3`��y狢,�k��z���#����k�V�G�B����J@6nH7��<"���n���W.�W,����%"x�x��E��n؋�OwP��L�2q�S\عc� ��#���x�̙7�5�j�(E�&n'l��(6@��؍��sm�ZD��H��$�v>���R50z����h�K��_�����B�߯�@k}�5L�J�&6�.�ܬj�m���_�wȍ� � � ���(��ܕ�b�3P	��|��8ت��8(Y���<'^��.��ѣ �ü����
��%�����]�]%�Z� �ͩ'1s�L��u��ID�IOOǜ�p��)΀c���a����ǲ|�1���o �X�L�MM�t�r--���[r.��Cw��b�OL]�M7�@�Tq�J�q� =�/��F;��s�=.2�3&F��.�������#qm�jl\%����k�>���ntO룉�c��.�'�{N�bH�;s6���� �H&.]���&ܷn-�S�tm����ѻ�G�w�G&X��W�/ŕ��>�(^��@86 ���1j�(�{����W~�aA*�t�)r�>ՠ,`%k��\n�ٍwR@AAo�MCg{��Tm�K��z p(3�@���=�dxe�o�������IӦ� b�w�_u.�;�ښA$W._���qx`�Z�=x��ND̙6{&�]��֖���۫c������.��vc�V���X6Ɗ��P�����{��8�3��IV� ���pW�"EQe[�eK��ܖ����ǎ��wt�an��|�ϳ����;�s��ZIJ�7p�DQ�DQ�	� �}���UY����D-�
x~VU'��s������y��@?��7��i��B�{�R�>���0�,_2��=� UR��,'��|�g��ӧO�ƍ �Ał
�۴�,��n��$~�r���VXk����v�~��'�>�l��;���?ˈk��,)�t�x�ܶ�?����!�"<��={�֏���A���z��L&X�������N�S=�k�;*{��N֯_����p㫯A�3<<������ T07��L���|����=]�%+�M<��9~L!�B!Yd��Q�N�FX�ܡ�jT�A��/�c	�9��Y��fk��ʺ���o�>��a�s�CM�'$e�exu�wp��qR�G)0>x��a����q��Q�ID_b��m8u�8H~����#jjj����K�M�c��{cY�"w���xl���7��d
��ڊ"�<Ei��TЅA3��I4�A*/��$R[Q(
ͅ��M�pFc����m(.N\��"k�k��Ĺ��w-�v�X�v��=^h�3Z*qI�5{�Ե]��.wmr���<��%΃];v���sx��B)d������g��ס��$�����v[��vؚ�ڇ�4O]�����+6ۮ���'�����?����>~��_'�w*l��OM��:1X_�'��I�w�[&"��ť��9	B!�B��X_fb�I�O�N��.�nu������������e�C�y�l�W�}���Z�-ES�b�I�V�坻pp�LLL�B
���~>p���uܺq�d������Ԅ�O���GL�۳g~��_�+�1��ϸʴdް(�7�\-M"rǰН5�d
��-�/J��l�%�T��|V�T��*�� ��H~d�彳�G����b�Xb0-�v�l��N�X>�퉢�]�����rm�	��2��n����Ů�xa���8~B�B�\`||W._���;046���Iq{�\۝������]۽�0�]۝hiY��/<�s�ς���͛�jS�w�V*b�����qA?%����čA��En�Bcx�%%"�H�k��j�ΒB!�B��֖bL������8�Cw��ļ5Q?�|��4�>���<`��;==�c��@���=��LR]U��݁O�����!��9Cq=k[����?0 B2Ŷ�w����h�'������/�"k䣁Uf�+��*�5�r���4k�9`�����#�ho,�W]S ���<dQ�����9H%��bj�'*���� f7�����[wn���E�u@�v�ص��ێ�%��$��rc��n��m��䳬���bb��w���Z`G�2�ɶ���կ�=Ч`������l�\�ni�k�Ҡ"r��,����D�
�vg��o���/c��Ey�����
'�L��M��C�����P9�!t�D�U��=:�$�����PB!�B�m�c+N�I�}�T�C�1���s)vY�I�:�X��m�l^�����q����`պ5�^TB2E]m�oڂ��|J�!d� r��~�-��?��^Fo?��HfXTW��m��{�6�z���K�={/��6�2���Xz�=(�1���.���ҕ���X���5S��$�P��gT�i��BII�+q�=@��`�A*�c�ʌI�nՃS�n���>��#��`��%hji������ۨ����w�M�vc�A\ۍMA\�ѹ���y<�c��y��%�w��5����Zk��D��a�vC/���w���O?���!d."�e���?�'o���؅|tl̼�ˊk��|�\�>w]���e޵=���=�������k����O@�s��A��?��.]��σP�߯�QC`'�>�L����>:2������$!�B!$�hZ�]Rw8,w�l��_Ja��r>�J0H]�m�1E�yBII	6<��d���&<Ӿ�����2��5q}{�W��W����B2������}LOѭ:ػw�.p7���XF�0�1�S�n7��qsw��c�Ǟ�Z� �9(p�3�o)�4���P�z}ø��h�G��2��L���ѣ�{�.H~�L��-����P�����̵=)7�#ub�	�-�s׮�qzRk��K�f����vS�n�gݵ=/�2  ��IDAT---��gw`Wh ����������?}[�L���H���_Uۏ��>L�%l7��&=�so�u����h��M/�et?���a�LLL�U��[��PA�<]�
��]wX�d����*M��v�2����XW=�/��B!�B2��R������B�']�J�$�5������=_h�/y�l��?x� ǎ��mڀ�
�	Z���m�n�E!sq�s��a�������o��q'I����}-��vD=���׍����=ch��'tw���9El����A��[��=���)(p�3�!�H\�|�}�f?H�ωA�C{�\�{;gg���VbQm��$=�v�Kz�]�e��x�Tl�oʞk�T(���P��rѺ}q���-vm�|q�Z�⎝طg/���A!�q?��{�����? RY�!�(���^��Y�g��=��h�c�/-+�k?�>>z���������~�;�	
*5��Tc�*j�ud0���_���%nw82�Vڈp�i!�B!�d�5U���H�^}�1�f3ƒ���r��	B���y@?��/~�ᇘ���]�@Yy�lh!�`Ų�h]�G!��u�=͡����zN��}�~��ٰenݸ�ɉ	���={�����=����D�n�c�'��$b�'�����X��uS���!(p�#*J�0�߅�H�+a�-lפ_*���U�@�C��08eE8��<yD=�ܸuK�U�_���m{�)nw�G]�n �k�mC q��Mqx]۝��Ko����Ч��n;�D�s�\���w���p��45c�Gs�2��>}�!^}�UT-����`V\�eq�˹��&��]۝�عk�9���~��'N��W^)�A�p���V�_��A�V��g�'�˖tNH����{�B!��QF��+�%� �C�Y�f�%��r�����wOI��g��S���A��lIN�'$U�`I}#�suB�<���I�|~�~_x���%��X�q=�]�D=��~��ߢ�8.	Η�_:�M�3\�/��0��rs���M�D߼t�7ւZ��@�{���с��gwxT�]��.)��v�`$�UKi&��P�� �>��LMq��|`պ5���,��I��-�"l���K���\ۓU�Ɋk�Dt�ˢk�=�������nۃ-N���sm7��[7nƉ�G���B��>|���z\�><�ؚ�k���eB"V�HGܮֵ=��`=�>�܋$��o����
���"�ֲB�
��Ml��<��]�O6����-�XE��Gk��M7!�B!$c�o,���0���m�mgc����4��rq�b�s��B[���}<x>Qς�J=wHH��_��zp��iB�|���s�ȽdU	����k7��ͯ�����Z��oGG����#c,�5��Yc�'�k�m����K���C���1V&��=�h*�H�ؖ,���v�s�ҥ��b�l�w�C���a�����G��G����v��z(�vȄ�]�!�D2O\�M�e�RѺE��Ի���q9\��KK�u��۳'�u�B�"�[o���bhH��WSq��h�8?q{�D�����`�v���׵m�v=tO��@�"��ݻ�+Vx�� T�A6s�f~�����1X����1�	u{=!�B!$S�/���ӈ�D�$ͽ�vc,-i��7��O��웙�.w?�I�s���#L~Q��_�6nۢ�߄�C���(ӊ���#cB�5B���Xݶ7o�!�E���߲	��^ Qχ~���1���c� @9!l׵��9Ck���_�\7�;} ��<�4�/1���5He=�]�T.�T�]9�dKt��:��C8�vQ���%l**�ύ�&���E�����um�}�o�og���]�>�vm���\��m�曻�ř��D�L,���q�2�vY�]����f����`����d�^LOsV!��]���[XPQ��1�L�L���q����44���{���gB�t���G�"�����?�D-b��}����ì��E��=�~Խ]��`sd�LO%rO�1`e]3n�p50B!�BHf(��������B#?(q�2Ɗ�t��š=S.�n�3g@�#V|^��������*���s�A!�x�v����Q|{�6�-�֭�7׿����Z�;�G�����3f.�N��F�c,�O6����&�֮������D�[6�k�"����=O��R��i���H�4�#��Y\,N�A�t$U&q!��l�<8e��O?�C ��6mt���X��r������>����ԉ=L,�Y�vY=��>�"Ϋ��W��h"NK�h���g~��6{��G��%��-).Ƌ�=�=}���@!�ξ����O��/ޣ��zY:��a��abú��#nόk{��l��{�fGp�q�&,^҂G;A�"���o�F����B����hbl�N���ܯ�l,3�pc�<#�n��q��B!��6+�1<4�����vc��e�9��W��&��`���՞�e{�졁N��y�V����Xֲ͵8}�!���9}/��&�&q��2�}��-�q��4�Z&&&t�;�7,dw�p�����x-�/Ku�!W��EKU:g@҃�<aI�F�	���%x��̹�)�U�]�.�n�C�_Ygg'�?���½��L����yn-2��<�mv#^�(� �(ϴk�m��`�q�qm��M���.�w�m�pmכ)qm\e��8��ك��"�b�ھ{?ޣ߸Bq#���}���w03����������26[�����;c�9�7�������Z<x�;��޽� �f�s���;:����67-�CR�n�2���u{-!�B!$]��Mc�ے7tN��zXr����9�@&l��������K+�}��' ꩭ����A�lYҼ+Z����	Bqs��i|��W099�GO���кz%����@�"&���w�����|vgϥ1���]�W�����a��#�� t��	�y@$�����r��E����C��.�Q܁���/*�r�̰o�>:=��%�X�a}�\�MSp�!��#^����G%���}Kc��v��ZM��]�ĵ]K~�
r�ڞ�b��]�vK�%�6Y}��Y� n*^��8��5	!�x#�����?�+���X��q���.ͥk��~YdỶ;i�ݷ	� ��X�J܃�矻B�:mw��*xRe̍�)2�=��RՀ�A��B!�Bңd�ӎɵ�>�<�|�g���*�M���0�r�'N�����AԳq�2[�zy+���!��q����꫘��BwO7	��;lxf3�� Q�͛7q��y<���y)JOEƌ����c��E�r��Wfh�`�/րj����=�����8��+�K��]���\�Y%.��@�I\��R����s�0��6l@Y½=�E؞�v�����#�����k�`]�k�{��$�qn��S�!�k{B�8�t]�ݓ����]/���C!�������������������Wn/�����\���2lW|z��0��vmڀl	����o�����<x��O���ڸ�x!�+������ʍ��/�����F�1B!�B�cqUC��(++��z���'��V}����̱�h�G�y�l��d��� �YTW��eKA�l�]��׮�Ⴧ@!$5G���?�.|~=�� $,��Z��g�cr|D-�?#�A���X�|�o_ؑ+4��F�:���e�gC���ۍE��762{(p�V.���x$� U½]���s`���w��"��M�th�C�_�x7n� QKqqܽ��"nw���\�m�rm���]��h��k����|a�S��vmw�W=�x�-��v�:a{�˙^3���o��-��k��j�x�{��8q���!��azz�������:�cj:�<�k�v��P���ꚳ����� �{��^__���u���������^��
�vc��RirQ�ǀU$��Ë���P�/ !�B!�̖����POQ����?��#j�ի�} �����3�Y�~��B�%Z���ѣGAԳi���쨩���m;���} �q?t���x�7�q�,��B�a��v�"�Z����ӟP]w�1�\�n��W�,y���q٪k[k8z$(p��F{��x������q~�|E�H|�-���6k.	a�9�%�,ȝ�*�PAii���%%%���&<�wI��TP�%u�6�
m)�c�����zLQ�Ġ=4N�xow/����T���񑆛��+~@�O���_&�����>�"�(��2��m������K��S���e�[��������./���q��m�`rrR��/�ѿ���e����X�;��ק�~�Ǯ�~q���K�7G*�]|߆��155�����!���a�O��B��v�j����]>p!o�$���gltT?��]O=#�n��0����8~��_d�}�W%��ݻ8qԲ�n�z�4��`4�����A��2�os�!p7�WQz���0�֍�.�X��VC�OQV܊��|�!�B!s��� FB���XEvc,�������6�!��Bth��Ǿ}�011��o�1�'��U}N����n�8�d�W�T���ÃCY�{|l%#��Ψ�ǋ�Q6�Ϸ��9>1>���,�����,�_�۟=��;>�hEh���:�s���+\[e�����8�t��'ר<�D�Je��n��R5���;/�=U���;���^x�E\������W�[#�.^o�@��|]C��[��F���!�Vy-מC�����y./�ȶ1�������n��}�g���9A]��"B'�&>W��]1-UE�/3½�>;$�R��A*����pHN}�g?R�C�D���\���1!��'U������t�/>�m;w���~��n�� ���t��(�m�W����_c��u�*�@MZ��vm7�o|�%�n\����-ǝ2�2Q �޻u���(���tm��/�V���K���M�b����X���[�n���*�!�ljjRR�ݻw�b�
�B��U}�B�.�����J�Wy������;�⚯��.+?~�e˖)������G����w���\\��:�=t�}��@�ziڮ�w��t>|�M[6��cϳum+�����r=7��ux7˄����}''���؇��Q��{��T ���O��;w_}�����X���:g��`���1h�����ݱܠ�������~�f�!�B!��)/������D��J�;��~�v��A�-V�<��5,�6a��KA�!pW��?@+�Z1����q��+�
���*���~����ֱ�s�}�j:p333�qB�j<Oh�k�
��]|�)���B�y'�s*E�Fݪ�*?{q�&p� [�y��E����l�T8�j41�B����c��PW]c}rB�
T��}4�w�0�w�|sg����ጱ�&��D�F�:����?6Ѕ�e���etޣ��4��ڄ�2��e
">_������.���> �@�ҽ�(4�z�xq1W��KL�nܠ��uٵD`����v�J�����qM��܆���&M+5Z���g)lO��%���q21z��v�g� q��l��D;����L^p��W���T:dB�\B��p(vo$Dڏ��$��A�".Ll�B��;̽�l�~�*D�A�J]^o��y�N�m;��'�Q��^|��'��]�-�P�^fPF7���=a�pn7��81H��,��6n!�B!���ٖ�D��Y��4�r&�5ۄ��#E��#Ih��kN�B.�/���+W|����XS�˪@���Ps�8�d�/����M�^���4��`�"�!:k\ܬ�n���Z��?�.Χ7^����h}}����ʌ��6A����FI�Kձ�C�.��T��؅�Y�Ω����1��ÙB�g/�7�~q�*H��{{z�׿�5>=zh֓��d��%���������v���U�����\��.�+�㩼�����re�[9u����[�Z�������{c�İ�ޚZ�)�1i���=���cc��\�K�j&���qU�A�El�o���e��Vw���$�A���`�Buf���O?Q�����L<&s�tm��{	���b��y�<�k{ a��<}�voa�۝��{q�g�f�u�y�����I�v���764�~�4|~�*!�d�����K���ft��J"��{��ҵ�u�y� ���f��v[Que��˗�@cS��<Q�޽{�����U
�]!l��:��Ӊ�շN
݋��UIa��/?=$V�R�&�B!�6K�F0	�7�c��v3�n��Y��*v�2�rR(����b��\�ۉ��۶���|�;����S2!����s���/����N�����+׮��s@�!�5B�w�w�m��?̶1���՟5ӈ���]��(k���%���
�RQR���2�^��R7� �u�t���]�m_z��P봐�%;;;q��Y��n_���2Gi�\�=��β<um��~Y=q��+.*�ˑk����5�,��;
��.X�`!�5/֗�"��y���+�TWc���l	�d86#����9֜��=�^p�#�(�|�U�����@�����>}/��r^*eӍ������4.�w�va0����`]C1�~:B!�B	��E19�n�g�t�sf5�r����Y�B7�J/�e��hD-�eu��e $/>�<���s��N!�������?�g/Q�L��x�,��+��cϞ=����\A#�g�����c,��"3��9C��>&��@f�
��R��Xf0���I.��� �]�F�p��}�߿SS�D��½�JP��x,���p��ZC&\��(�ڎD�!������k���\��C7����f�����,�i��̵]<+-)��͛���BH�8w�ެ�ח���J�޵ݽ�t�Ac�µ=��ƥ�y�3ؿ���2��
�]9t�.p�m�ww�ٴѹI܃�rN�^9ͳ�.l}��M�� �B!����o(���(�+*��&��Z;S^	��&w?��\�%?~O��3���MAH6�mG��.}uRB!����{���ĺ�k���o@HD?E��.�9���y�]�vt>0��X����ٵ�=�%:ࡁA�.jƝ�i��Pஐť�-�va0g�_"����V�T�`mV��6>� ׁtVM��UX�pa╗k{\�l=Où���]�����;��C�ni�G=2���k�����<]��u��k�f��n-a�Kvn{��������c�����&'019�,O[��]�%�ȵk{Z��4�P�Ov����@�q��A��?�3����ׅ�0�x� �n��rR%WK�V���K�M�I5 �B!�������d����qc9�8V����X��Su�
E�tG�	��Y**`Y�
�K�cay�]�
B!����_⹝;�t�<x�	E$+׬��Ϯ�y�D�F�s��]�m^c!�9��h���֒���+?���ƺ(��nVP������S��s��t`p|Y���2w�A*#�Z���f���_�ڵk jY�q���ߵ]s��;���;c��칶�c5�vm���]�ʹk{"�ϵ�-�w���m~�s8r�0&&&@!$����{�����/���}rQ�"�,��{�!㱅��&v�Ǻ}��� Fu�����!�u�ʫA��1x\/��E��;����Ace����@!�B	F�D��\�<��˾J���;�I~Y�P0�L��e�/}��Q��vq���:�-]�cG��%��\p��9����12:��~*5IjDf��u�v�
�:��?��?���B=o����X��Bg�ڜL���=$��3�Z���wEll,��ؘ{�A�A����t���ͅ�21s����Q�4^RхA-KW,â�Z_�v�.�*���)�����-�gߵ�v<2��,=��(2��E��f��C�[\�5��C���m�l۴ϝ��� !����i|��x���
�:H"�k{�D��(�WZV�_~I�5�����{�x�B��ۼ���s#R��܍�4�
j^KFl�֋��	8t�B!������zQ^^.u}�2�*J���X���·�ub�Y>1Z��A�xя"w��Ҳ2��YB�P�^�|f>��	!�䎃���;�ctl��bM�Z|}�:&id����nttt��^��|`&���]��c�&���]���7������nT�Uax�ZհPஈ��S����`r ��E�����Rŷy�[�(g������C�@�Ҿy�[ܞ����8��947]�e_o�{S��[l��"H��u�A��pme�˗���C<~��Br���0؏��*:�'JC܋e���c��X��gBp,������8~��r��1������N]��
�ۼ�L��Í�ZH䞘\��
����U�@!�B!����o�_5ʚ\�c��� �v/�, ��ݗ|�E��Fc,��Y��Ŕ/�Ԉ��+/}��}��-!��q�=��~|���c�ჼ�����b������uu9rD�!�=��X�P�1��c���c꠫?M�d�����;�Q:9`.3t��s����U��KǺ%N!@�&�ҥK�w��:����d/̩k�=6�k�D�n��<��қE�b��2�hx��)��k��m�]�5��XX^�Kg΃B�:?z������U�����ڞ��wx�y���4ڔ�Xk[+T`���q�����t��������2��׍!�|���KZ����*�{��c��m)�9�O!�BIA-�0�BT0c�p�v�>�$���ܝ*�e����ٳ �����ׁ� q�w���@�BT011��'O���_��3 $k7�Ǎ/����4�>��XUUU���v~/�>f�=q�縴�2�;�*r7&�['�k�O��џ��R����a�'���RC}=�%�	�\�ܽt��=.{����P�'���h��`�̳a�f�E�\��%9��v[,��z�f���p�>$��QH�y�㊛�k����0>W��Ƀ���������lZ��!�����+XҲ�e�7����ӵ]��`��ڕ���v���';033�C�n��B�t�e�T5��A]�+�I=�*mcc�X���.&[	!�B!�Db}�сni<�1��oc�1�2����Jn�/~������Q�ʵkPV�U�Hj6�߀�7�E?!��C� ���lX��o|B�(�����m���M5����y����yot�~�Q�>4��Ț�-[�����[����Oc�/	�
x�9���vG|��3@2�̠U��{?���L������-˗�_�Ե�^&��pmw��5i��k��===�v-�k�~8~���2�k���W��$â�k���۞�����!������/~�K<z����场��>�>s-"�G�}�X���E���a�F\��9�.^��G�����3�0���m��'OZ:��Wߺȱܠu����{����)\�!�B!�x����c(/����c���T^��u�w�0W��lݝc,���� 456�<R��oRG!���7����P_���� ďu�S��?:v�.p���*l�s�3��˱��]���l%hy�ݥ�D02<���b��1V(pW@K�(Ɔ�]\IrKR}��:g��禘� �l�O�>��<*++A�P�ؠ�ӆ��tޔU���k��c�ص]���U�+.�k��=�gQ��|����[����ܵ��n�v�ٖq������BH� ��}�!���?��G�΍.iN]���fKD8��]ۃ��˻)pW�p�?p� ~����B�}Iz�A*�>���]��`W�����ޫ@!�B!^�����D�՟c�e&��}'�ܡC�n�c!۹���=��ܿ�.]�{�B�j���j!�C|G�m،O�}B!�C�ɓx�7q��1LpE�C��4/i�㇝ j����n444����dB�1b��4�C����G��n]�9�)�E��������N/H(pW�h_ a������J��
�}���/���l
��l$��Hq����>�ʵ��!���v���õ]"D����\̵ۡ��䱻]���/�P� >|B!����0:N���v��ӄ5q���{�ҵ=xl����+�t�2<�wDN��_�>�x۽���`��Z��>w_[�ܠ�@�1X5�׃���Nz�xA!�B���M`&�Z?c,�jSAͱle-�3r�~�����W��]�� �q�z���qh?Wi'��|C�O>x�|�U|z��c��v
�bc�򗿜�X�9VPc,_m�Ĩ:̣ñ�+@�C�{�i��`hp@_fй�� ����b�nq��!vW׌���Ln��3�P�� �ѣGAԱz�Z]���Kݿ��黶;��Brdյ������kΥU4���ˆk�����ϊ��c.�DS]=��B!��ݻw��e1�����u\ܞ�k��a>���Up,6�}�5���/��������>�<��e�<c�I��N����^6� �נU�������>���B!�⦢�C��()-�:�K��i�e:��_��+Ih��v^�sn04�Rˢ�Z,��$�w�¹�g111B!����8._���}g/�!^�,[��j��������=����O���g���K��}w��l��OQ\�SL����1v�ȗ�%œ_���{�A+.�v� U|[�6�%g��g���ӧ ���>~�?ϕk{�ܚ:6���{���µ]3�����0˲��.��uo�������A!$�9{�,����(-)��d<���{�{�l���!n/t��0�Yrmw�nܼ�,܃��!��3==�O�����uW�M�u !��l�)t*n7K��j-!�B!�8��T��B8�iǸ�+<sp�jݥZnЯ�Ν;�v��:�lh!~�]�O=Aww7!��/O?Fcc#V�\���n�/V�_�Kg8B�ΝÓ'O��ܬ�V�Ξ�Xn�e_1ͽ�Zʼ�E�.&lnj*ƕGS ���=�,҆0������E�*�[\7� �񭵖ƙ���P�:::B�d�e�+P]S��s��.���n��=���"K���z��K��N�x@�v�_nѺ,\ۍ?a]�m���69�q�3�pp�~]�E!�0������/~�{��k�G�<.����\���⋋#x��p`ߧ j8q�.p7(�z����������?@�\%���d�z�1�k@=!�B!�ɒ��ޑ 9C�r��֜��,K�3�kn0SBw�^(V&j(+/����.�QW[��E��8q�B�k��W_{O�{�?�Bd��^�k��bb|$�LNN���w�y�`��Y1�
l�%�oK܃�#����)\	
�9DӢ��1O� K&� EfR=���R��z�,No�ʏ|qf0��:�nhϝk�ԉ�ܷT��ڵc�Q��Fyn\۽�SV����ڪص�_ ,_��n���� !�"	x��|��W���q�<}��0�9�ӵ]���۟{Gb�X�ϟǣG�����3W��M��3He�c;����=���@��&<�$NB!�B���w"�#ghwp���}����G��DC����|�;�����k�~4!2�ul׶طg/!�G��o��}GҀ�H��m�*|}�:�N�<�܃�_B�pu���ːǵ��7���&�Nw��jAVf+��j@�A�{io(���8��+R8�[Ov#����z�⽐j��B��2��T�/^�ÇA�P]S���by���ڦ	�ø���oE����rm�8�;�i���k�Ȳ?� =�����)��ĕ���aQ-��2D�R��e�:�?@u}��z>���E��*���=h\��JlںW.\�=bb�Hڿ��#T�Lݚ~�'�t�}�[�0�,+�M<O��`�R���A��!B!�BH�����QVVp�gs�&]�ٹU�U��]�]1�|������K�P�8wW�[B���/���GBH�133�S';����p��9"c��u��ŗ��W��ӧ��ۋ��:�u&rx*�~8M��ew���}hw?�����j�&YC���.[��q��A��=�����Lw$� ��%.�R�V��ևI��T93ttt��Q!k6��N�"�B\@�n�C���":w�:�k��#9$qR�vg=鸶'�е��[k+��eµ�-�w�E۷o�BB)p�����ܣC�;�vyd���g�����+6���θ�v��]!'N���A(�A+w�#����C���=�du�r����X�e �B!��-���I_Мab��)Μ|kN�5^��P���C;s!7�W��cǸҜB��.GyE9����]��100 B!�G__�c��K����� �ɂ�J,^�D7P#�gllL7���O~�W9����]F���Ksk�s�&X����tpO�7L����M��7	�
�sH�t?F-.n���.^KZ$���vr��`&�4^<?z�(����u�J���� �+�vHE���.�;�|��]o�!��ˤk�S�n��̵]r�b���M��q��ELN�B
���AUe��$Ǯ�i�3�ڞ��|D��k�]۝��[W���	]����3g�d܍�U�V2'���@U��O�.{]�����{����c�Z��B!�B�QW<���9CS�n:�Y'�5��rp�c��O!�S!&�u�n�{;�SQ^��e+ph�B)\�~v?|��<~������C��	�{
��ܖ�1�s�碤s�!rO��S�bELc얲QP�~J9����Eq�8��e�*Ѐ����r&�-��Q9`�ξ�^��;w�u�*��%�
�k{n���횵6��Y��[ږ����k;q�����`z|
���!���gddCCCh���Ӟ����rmϥ�<h�k�W쮗^�G��H��'����?�K�z&�vbݬE����N���{����B�>:�����; !�B!$���S߾�s2m2i�tp/
էI�$��jnЯ����ϟQCuM5��@��ﾰ�!������#X�d)�!�+�bxp$�����WUU��=�7�}e���p�����eyC�?o����� �
�s�Ʀb̌Π��18�y/Q`�������Dŷks>,3��}	��c$s�.6ѵq����:��}HE��x���6y��]���tc���5�µ�8f� �&n�����n;N�k�f��~F��C\�6�]��� �B�O�>���8JKKuA�A�\ۥ��tmV��}�XU��N�l݂O�����8H��UB��d�Z��`5��TԼ���`��U���A��bU������B!�B�ʺb������ܞ�Ni���ܽ]�:��E�2
-7���۸�-��ׁ[6l��W>���B�����ʲ�_�.���+�d��5�z�2H��uBO��of5痩��i��m�wHc,i[��Z����� W5���4�?����1=.wr�<�mU^.>�p�X���� ���u��15,��E}�1��*�������d��0��y��n��S��)"O�3+�vs_.Q|"*�<.�k;$e���'j����[���|B!s�O?����]��|�s����У�tE����#nψk{��\��[��l}vΝ>�{:::R�1�Q(�V�y�T�8�/7C��+s����]]U��Jm$��2B!�B�� [�#7��7�2�$a�mX�D���`.���E���������@��ښE�,-��@!d���ߏ��ZTWUc`p �Xi[��.�����#�����I�c��.��Ԙ�m�7�c�9B��7�)�9�=���AR@�{����d��r�0��b|1S�.h	;+se����۷q��5�oڐxfum���S0���2d�v�ݽO?�[���C��9��"xM�ڮ7��ڞ����d��ɏ�T�k�H�qI��n�}<,�k���˖,��{���!������4<����u=ql.X.�ϥ�����
�}�
�1::�S�N�?�AN��a�3Y���A��uҨ�=���D/q�&���ղ�B!�R��`4	�3�����Ͻ�.2dY��PyC��3���g�p\B+V�����Xמ�?�}{��B����x�7���A �ki�rܻu$��`�҂XYLP8+8�ۗ��6�[֟���l��L�|]�#ԗ�������-���}�̅A���pg�8ù��E�:�/���{|���=I��r�d�pa��J�J���-����]��h�9�'��b�]����Ԯ��mq]ۭm���g��n���n������ڞ���w�]�%m/))AK}#��� !��e�<y���Ge���$J�����YsmO������_�k�3nqK�._��������w'��
ZO<D3�UK�X�p���)n���	�Ep���B!�2ߙ�N���c9Bc�碐��3yo4w�$�s�~�¥p$9VErͪuk@����z	�;N1�O!s��}���z�9��x�XY�n-��E�p���91�R�t*c,3.x?;��u�߃���1��E�?����%��Fyy�t�JvBk���e������_ZǈT|����R̞�z�ЅA+V�BIi	��v���H{��C&X���!n��_�OO�6�B�`��k9pm7��rm7���gp��AB���8~����1<2,�N���vmO'��];)pW�����/��/(.���@Sf���[���T�����ܽ�����X@$A�"��@!�B�ǈ��b�p��3�c%�&�W{v��*�xy�6Zn�/� j�k�Ǣ:
8��%--���Eoo/!��]����r|M�x��467�zQ��Ar��3wٶ�d���򑜈�9�~�S7<<8�������Z=�h�D��7k�"dO&ӋBX���`b��O�X�����9��S��u�������ȵ�C�̵]V��8�vmw��)���,�����cȺk�}kC]�߹��B���ߎÇ�ŗw�Q�cK�4�c�H�wV���;VO����k���6���155�[?~��W�b۶m3�4�}şG��W��#��WK�#nQ��2������.!�B!d��^��:D�~Y�m�e`�Zͳd9�B��m����܉�֬!Vĵh��t�>B��\8?|�M|z�W� 6ZW��Ջ�Arϱc��?�)�G��z&����XN�v-�O��׋\ۼ������K������!�XE��*���<�U����Uk�)��~�j6��:u
��� �G̮Nq,bl�k���{yP�v#6��=jJ���ܸ��"x�{=�eڵ�������5mi�btp�B��=�`� ������y���.���-��xY�oYy6=�W.^�-��ELwٶ�hJ���V6P%��8��_7��[��2p5=,�Ț@!�B�����c���_��fX����/J�nM
��;9�V����v��e}������� �ʋ�=���N�B��@w�>s;�ن�W�"&��W����03C�o��}�6nܸ�u��e,��9�P�X��C����Z��L�n�6�	]k�7�gM�bt���}A>c#!b��C�-�cWI�u�j6��g��am{{�Ea�ʵ=�I���x�>�wm��%q�rm��އ�]���{���z�ҥ8�!d^r��A������%_E��(�^���;��m�N��"�[������|h�|=�{_�r����T�"��D���[c�V#��h���sp�B!�����H�+��3�:¹����=˰�]I�Թ�B��m;�<�X�b9JJ��1������8���@!d���ݍ�PS]���~"(�(G�t� �[D��̙3��]�mn�M�Mf����n�O�7L�����T����qq���,����(/��]n��k.3h[rPsX��pc�q��Q=���z�2�B�.�Be{n�6¥@<T՟�c�[Uu�>yj�O222���N��s�%n�z�L�n)��NNOIE�1��6!�k/��^624��;��l�v�L.��3<8��%mu�[�ڃ~L��va�B<�|�z������1���(�[8��ttT�(����$*�]\o�o�����cW]�������������=�8�T�?�֊��|�޾����m�J�x�9M��� z�{PV�>'��<�]$cn}�m����*�^������r��鍝�S!������p�z�.*���~/��%��c]KK��{�a�)�z\�[�U����U������c����� �B!��C�F�~�5o�y�ܭ��d�<�Ù3ķ��W��T��
��h[��XY������B�#';�Ə���C�A�AۚU�+B�����-��?�k�2�rN47��~�`K����C�}XTр�QcyA�{�YU3�'bqy3OV�lk�������ݍ�ĺ�d�X�m�}�?~��K��U���'�u7-nƂ��1V\�]\��{;��Qص]v������������!�����.DF���f=�����r�����>���Y%�~� Y��&����U�m_���_�^����*e�Kq�UU���MNN*=���Re"o�B[Q�8n����[u��^���.�s��{�$���_v�b���M1�N��.¸�K�SS�(-+Eł
�}z�7���Op켏{y�wVK�k����Ů���y�]f�����$�������o��u�x�<2��eg�t�DY�DYGG~�����@S��1�J�C��#����S������'�p!�B!����B��_�sr��d;ۜ��o���(�ܠ_�Çq��]=O!C����VF��&�g�Y]�dp��&�|���U6�2<8������q������7��=59��ё�c,�u/nlҍ:��ef���~ܾ}[I��H�����J�Wy���D��7*�]\g��OLL(�0v�u�2dS�ً���
�*��w�?�_����x�+ku�����]���*��W�;/Py�1:<���^�����5���Q&Ӯ_�cT!�s��W��������?׍�jk�N�\\�����ͱfk�e����iIM�|���=���Р��=�Q�2U��8��35\�Q�e�
ݓX��HY�K!X	N�>��$za�D�@t�Ŀ����V6�^վN��01��ş�']��]�8��K�l]��5�ㄫ��F�Q6��Bq��\��.u9�J��g]�aQ]]��Q�8��sm7%�	�{R]g6�ɣN��׹c�a�}[�dmw���m�ܾ׮|��VVV*�����j%u��1h��~q#�5h�����c����PU��cW]��]�`���W��c����^U�b�l�ʖ����q?��_�����2�ۼ�"tKaoy�~�ײdI8��4���?�޼��-�������o��������Bs�~/�!l7b��\͋'�<�m�v��"Μ<�tQyo��{��.�� �N�a�)��r��������;���N�n�JtT,�� B!�B��CLx�&��	r�6I�<p�0Er0��-^�"�s�~�'N��E�^�qLU�3Ch�Jt��c߸u����ݛ��b�J��񃇨ZT��Ʊ��L�����z���x�Ҝ�+ηm�7�??�D[[T!Ė��y;qݭ��QR��cW]��'O����_�@屋q⮮.,�<x� �/VfΤ���B/��ب��|�ο��k8s�FFG�Rw_w�~��'������z���z�0�=��_��ŗi��{{чƧ�{���>q_"V���<�r�nc���n6�X���9C����yC���e"��"�
ܳ��`�Խ�s	s�����BPQ�\�:u*}�	���^��:�I����wmפ��Q�X-h=n7v��^����z��}?�D�.�vg�E�u�%�bN���N��\��|_ض/�\���	��L!��$��_ÊUm��띕�<e��� 6��ݷ� qY�ͦ`=�8y�<VL�\�f5n}���b�"&��H��B�8Д�z�ĸT4�@���Ⱦܠ��]��><4��M��O�B!�BH�����܋�},Μ����;,�ܠ_��s�@� �	1���.�t?!��Ǐ�{���Ǐ�A��U����>��/	��l[>�g�����:������qq���JͰ$⢉�Xj&��g�5�%������C�e}q�J����Q=���z������ ��u�J��m
��o�3x����2C�n)����p��sm�Ǝ�8M��!Z���[��ʵ�^��,�|n�}�ڮ�o�����Ï@!��%�֮[��/D�vqgnE�qmOI�]�5!M�z�XQT�n�{f�3�+@�4q��E���y*F�]=n��M�9K��ܓ+���|���o(�ɻ�B!�2��[P����x�P�<s�.c��
R�՞���,S����2E�� �o1ћ���&,T��,�/6�[�_~�\q�B��F�,p��-�[�_�n���u����-�=Zqq\N��9�L�!�R3����shC�+?'�;����Pʋal
D�Ydբ�I�/wl�T9��!�L>�vb�#�g2�Μ9Î�"V�l�!w��hy�LH���n��B��[�?�]�݂}{���n�h]�ׯ}��
w!��9�?~�֛���P��v��s��&�����u���˒��=���K�.�wٶB���4�%�V�GX���:�K�� !�B!�����nmZ�|��_�|�9C��$�z���_.�Ο?�����C�vbPZR���&��!��o��?xㇸy��DDg��6
���ݭ�mݺu����+���Y�cYs������ ���b\��]�Y��dc�6o����J]�Iz�,��P��\��{�CCS��8���^�v[��k����r���K�s��no�۵�k�(?�Mu�p�!�'������Eii)�'��Y�g޵=�"�|um��՝��7��W�����J�/)t��x,�U��y��k�s��r�ց*�C��Pl�t�#�B!d>�T>��ሴ� �����v+�����&��B��m�3i�E�!��+���K;w�tG!�'�;N��gw���� dy[+�^��{�1����]��Ps�nc������Jهv��f{��;��2�H�KL��
ܳH�Đԩ�ӅAs;1���\N��`���2`%ܢϞ�M�
Z׬��k�'S�n-s�г���ƻ��̵]Ҿl����ݽ��q��ז��8s�!�/�>�����yx߾a.��k�<�����^�鸶;c7?��
N]]]hjj�_���l��S�b�A�q�=&0<Ћ������B!�B�ҩAL}�ܡf�1�ΤyC,g�О�O�;�d�/��iC�	�$s,^��ee dQMF���!�)�+������@�9��T,�@��f<�|�[.\�������b3Ghbl2Ӆ�P9C�������E��h��r7�g���';��봗z�/�fhXN����^N�r��5W�u?�Ն�������=m�e}\�!�K�M.q:��\�]ù.x.\ۭ�5�E��fM�%������j���q���ѩi��p� B!ވe��q-��Ȉ�y:�����gA�J��`�����d՚�(+/����џd���)�;w?�я�&e��!yg%���x�V`���pf���������r��B!���9��@_�?q���cY��󆎜a�r#�|���c����|�� �g��V"xa�N|�w!�/Nu�����*�8B��;�G�ń���j����zߵ��1V���]9D��}r�7Vy�
ܳD{c	�#Q�I�� y��~�ۉ��%;�ˀ�ŋ�L��բfѢ�+�v] n/�J��p�>$�A]ۍz\��ʵ=�xoB nۋ-�.lw��;�O��R��������8�̆Mؿ�B!��t���Ż��pm+8�� q!bϵ}��vQOqq16lބ��/��+W��w'�ࠐo���l�xͶ
��@Ź��ʚ(nt�B!�2XU_���)����'����2ł{2��4P�s������½]L�&����K�-!+W����o�U�	!�/�1�4/_����t���m.�9���366��.�����Dp�6hW:���������`[���߱�Q�TE�98b��,��2v��Ig\H�\�8������Iy��|��ԀեK�@rOۚU0��LK�ε]*��	̽�c�,=�v�@�g��]e鸶Ǐ=*�<0���)i����zt>x���	B!A8u�$v<���v%����е]�����U���k�m~f�
8u�m@'_2�c��r���@�UE.w���dc��b5��B!�2�YU5�����_�����p�~���}$���!���l�|�2H�Y�b"Ŕ"�w�5fM�*����X�BR�����7ߠ���%/]���x.��w'����˷����2ǒ<���]���kk4t�8`�2KTFG0*I`���w�v��yXќ�����$se�J�jϝ;�{ZW�
��.uI7�,����0^'y�%�V���no��Y(��d�A�C /ڑ�v�h�C ��>��F�ڕ+����B	�Ç�\��$�'����H΄�<G��h����cκ���,VVϊ�V,�����0H�x��n޼��k�zƨv`�4�];�۵�����AE��1�zE=!�B!s���8�Nm��;��^1*�Ê�@+{yðd;?)��={$�,ok!�m}�/�ЂBHp�^��-6���/@�7�W�R� g���A�[��⢽�%Ϋ��1	]�
[S,�(��2a&[b��,19�﹤�|v��������(��.^drPʏlX	��������܄+%�s�v�gܵ]&��/��������m��ݝm7۰�u%>�u6ru!�2w8|�~�֛���1HA�v���ѵ�3>����Ѧg6�ܩ3 �C�{\�pk֬	5��O��t��V9�����f�8��P]ր�q�?B!�2��w%�}��\��R��&��K��-&t߿OQL�)+/CSK3������e���!��G�aӖ�().�����e��e�����$H��ꫯ��ى%K�x�D$G��Ѩ��;�<ٯw�}L�l������P��j;�g���FGFP^^�q!�;Nr���\7��\�_0Gi�ǕO�R\f0�X��*����Q�`�.�v��#����)�w����
o�h����*,w9�[��µ=�'x�]����{e�8}�6!������)*�+0:6RD�I<[��;;�]۝�o�@����������<�
���s�sP֗��rls8*9\ܭ�T�ފ��P�s88K!�B�\��T����.�t�<��\}�"W�$P��P�k�|��}���������cff$�,Y�\?g������ �B�r�dv�܁�s��g"������� �C��Ν;����'s&G�M�?5��)������?/��&�;���PRT�IvamP�����N�Ay�k6�yr�N�K�n�,����By�����%Δ�t���3SHn"sI769bø�����%����_�m�;��um�	ĳ��G�� �umO)6�o��S �Bf��c��w���{�\�º�;��vm[���rii�8��`�Z޺��I����)�	C��K
�d�A��h{$6�'��.�^��ec��B!�2�i�� �n�&Ib{cy=��/I;`� ��s�o�����I�Yֺd~S_W�������B	���f&�P]U�����˲+(pW�0w'��#̬1���,s>��ۖ��L��\��=��=> &�k(Ƶ'\��
�Y��l�E�U�GQ�/DJ���,��]'��چ��a\�z$���ա�:�<��k��L��̸�����k����n�k_Q�W\\������B�l�����;����C��:��rm��l9�#Lh�\ۣ��p�*�E�7n���@rG__�_��-[�d\؞��Z�*�se�U��i��KZ�b��i1�c!�B!s�%�Ә�;����˛����K�74���>N��a.ȶ�^�5�+���󍋛A�7�nڂ���!�2[Ν=�W���8
2iY���źI�b%,k.���A1�pu1�NsJc,٣Ȧ�i��V~��U3����Y�dz�K	x;1���6H���ra�Ǩ�R� /\���@rK�6��":w�!� 1��Z��5�2����"/���M׵QwY�\�]mפm����v��'=�c�mj_�3'��N!$}Μ9�w���.p���*�k{�����7�r9�|_pI&sߗʬ����Z�ny�d�J�H�{�Όg������qΝ��z�c[[�e��k�U][֒�U������ 	 � ��׍" &H"���'�tm�~��5�#���l�0���.)-���/���rJ2���4 �
Ύ�	w      ����1���5��V��M�:h��U�1w��Y��1�{�.�����s�[�1H/K��fk+2�<   �	�x��O�ss��{�Ԓ��h��*m>A :677icc��\����냜#���[}m]w���ۨ��ܡ�C�1�sQc����@������U�Q���l	�v�>f�>�A)պ������KmW�ڵ]��*;�ѹ���&��� ]����+*�v[K��;��j;K�>��S�Z��CL  �ش[Ϟn���4�W&յ�G�(�^���l�.]�L����1w�ܑ�G��FpA+G�C�������fpS��˥�Nfi�N      ��||�pm7�*c,�����Gq���+�'(�$�8���m��_�@ �|��w���v   ��՗_ҟ����/��������G�Gݼy�._�I�0�w����Cr�j��q#���ꬹk�ża����X@�0��Y�T�T,[�R;���g8�B�H��I��=(nܸA Z�f�i�����ۅ�B�p�!����vm']R�g8��k�u�<)�y)��y�qm�{um��W�;�$kV���H���   ��y���&p�,�n��X�k����۱}J]��=f�Yz���t�k��G	�n�M�Ȧg$#�,�)/ Q\��@��O/�d��'�2���      ����,��J4:Zt$�U}��M����e��Z�k�E�9�۷o��\>GK�+����2m�x��%   �c�m����"���&�NV��Z��FFAQ���_���<�y@�(��4�9����{۴��:��쏢������tR����si�y��GX�.Z�"f��w�Q�JA����7�|C Z.u�"	Ƶ]":���ڮS��=��i�]��:yI[����yj\�9�]j�ݶo�?�+P��L���   ��{��1�./���������P(������U�wo�����>��=b޽{G�=�k׮%F�V�L��*��W^|"�ZP�����2?R#      �p��\��(��ɸ�5r�FR�0���24�A��$c��^�ӗ_~I ZV��Q6�%�^>��1����/   ��믿�?��O�ۿ$�N�1���
m��$�?���t}�s��:1_��yV�vŜ�)v��3y��7���W�tc�C�f~�JՌ<P�tbp�0xsb0�ZeE�>+6-D�ѳva݇k�f^�6�v���*yK/�!���]��W���A�]�ڮwD�_�N����&    hX�����v�U���	�}?J���z���{<�k�ȅK)�˵�A4��ͭ[�Z���*��~�ٮ���pI�J�+�7� �����B���W�       ��b�F��1�,�����U��|��ܡ>@�A7>|Ho߾%-k�H/���i��S��  �����--/-ӛ�o�����!p������ܤ��{�Ǐ[��uC���=����}za�L;�g[Z���56p��H�jB�Ze�}qI���*I�J��GPJ�ݻw�Y�����.�;�����E��e�Q2\�e��"u��c?y���:ϐ\���s�����@Ф0Z���	�J%   ���~{�-�����~�LRO%BA���p�U~(�FFF�ҕ���ۇ��M����׎�8�I�c��Z*!X%�J!&(�A�����j� p     `8m���HfK��Rc,�C�z��Y�ۇ	��d�[���]������������-   As��M��_�������3Y_������7n���z�s}��ݍ~ukQ*'���w� v��]�f~.j����@�0�#����R�2�/r�p�NE��̆��B��F�i���ٵ�YF���\�me�g=;�S��pm���2�M�m�=���F��?�F���N   @X�������;ؗ�O�k;��cG>q�ޗ�ݷk��Vytm���!p��/��"�v��U��_��{�s�i�fF3��       �p���f}V.ҙ��ܡڵ���\�3L��U���D�����a���.ғ��   vϷ����VVi����Q���y��~G :�ܹC?����>�9B�u6%��KiPM.}|!_��)
����qs��@� sc:+��h��ف!�u��]�.e?��>�A)q]�Z�o���@�8���]\�5aC�p�������*�����$�#���|�rm7�U�ݵ���k� ʷ�ۤvm7ʊ�︣�C*��   ������\�cgo�,É�O��wmo��X7Z�v��W�#-�_���O��{�E��G��`�)���U2�H�@����$���{��rw      ����zB�¨ÙM9Vҷ�'o��k�Н=���	D��:�����KW����   �oݦ����{�a.��G�W_}e{�=�u�:�*a}k]w���-������?g�e�h�R>;G�:f,`@� Wg��9�8�nIm� �07��'�qu�Ş�$`Ÿ{�.��l6KK++�
a�Ñ�t����\��V��n�������by]&�'��ڮ�+]۹6���ѹ����k�y>
Q����ý  @$0���_3�tm�P��ޠ���u���iii�޾}K ����͛t�ʕH�I����x��,Xe����Un�*����^/!n     `�x>Kک&up�������=��:.yC~�0���A/_�$-��k���WޣG�%    l^>{N�����&������5���M�������n�k�>W���i�
v�/	�y>7���b��N������*�e�X�Fə�vso�.NE��!z�P�0xN��$v����s$�ϭ��T���2޵ݢ}�J���µ](s��5ތ���9���e}��;�Ѝ6��ٗk��}��]!�'�����n�`���U*   ��i��<5?G�GF�v����x��k�X��G� p��H��wPo+�]��N��_�q�nY �E��pp/��
      ��u�7�Upp���(� ��"�ża��C�0IW��c��7����)���$�N.�������   6L����'�����Y�ӓ�P���o��������煵�!
��~6׷�b���g�����l}�A�1aA�dT?��$Q-
�m�3� T�d�QO�r����u���'-�/�/��\�;bj��;�vN�m�͵]s��ޮ \��gb�Z}~�^]ۭ���O����   D�7_C�����]���%X�k�����{٣���W�_��	Dǭ[�(�z$�>v���Ry]d+1f�(�      �tF%n�qޙ���[����Y�Bخ@���u�~'�Y=�N ��.����  D���-��ӻ��ce�=y�@4�>3�bwٺ�ԃ�a�!t7���n�<��<�`�=�eƳY�J�t$�f�pJ�R�Y�r�n���V���۷	D��yn�A_���69�����K��5-b�v�y���.�]��&n玧rm7^��ۚu]    D�m�~C���+�P�pm��\��W�x�v��s�T���)�h`B���=���k����P���s�5��K��:	�UN��`389:�b~�J�      ��r$��w5����pM��T���FEzn'���s���^�{;  �H�q���c��_�+�����{԰��gnQP?}k�i���.�k���xs�
��`� �11��ӓc*FM�����S��r���wb�+j���y��-={��@tL�����D[�ΐ���l[�]�ퟑN�(]��N�s��vᵣ��;�g�n��F���W蛯�&    j~����O���>n+��*vI\�{�M�������X����W�֍���M7x�����X���un�8.K!X%۷l`����F��,k>gw���e���     FrDǇGT(ly@/b�L��rڵ��'�u=�upp�����/.H�SS����V   @�`�X��3��#�����f��\���7oR�T���g���i~嶎=o���2M�}lo�ϼ�d����!e�i��^��xo.KT��=N-(���e|��QGZ�	}�V̽?ZѲva�ŵ].��<#�3Q�-sm�
�%��g��zv%�Y�k��L�^(�.o=������vvsm��>96Ao޼!    j*�
��:y��E���6�*��v�{����@�!�o���Ö�}���y��b�ʪ�ra0�WR���%n���x�0?      ���y�3�&�e}ǒQ�=�tI��7�8�l�6�#��X^]i]� }��w?���&    j������1�귿!�.X�xay�޼�"����Ağ~�ib�a�i.�w������7�H���x��7�ժ�>��g{5J;���X�2�tDE7�v?Ir��~�,1�������V��ѣG�eem͗��.��	މ����J�tm��9�w����@�z+]ۅ���ڮ��a�����.�ӟk�f+�����[�tne��}��   ���կ~E�ӟ��W/�|ֽօk��vY�J��W��%�r��}iy�
a�k�3�|�{\���qc(f��=g	      0���5(Sq�ޔ�����_��;��<�@�0z��&H###T=�P�Z%    j؀ƑL��Uk�v�	�{t�>߃Z���h�Xe�v��\��]�k<�a�ͱZK�.N=ۣ��{@Ld*t&qa�%��1�~8$+Is]�e���w��&�XZ^�ܿ�?
�t�Y�k���BpI� \��7W`�uum'�c�ǵ���� ^�v�h��v���)v7��|X[^����s   �����z�)BUjأqm�R�&�v�drj�5����;�p�֭�4��	��z8p���-�l��A+bv٣����t��      |&�:�2Μ!g�e�7��)�~��.�c�^��"���U�T�Ax@��N~��ߡ����   �����/���|����5�t���J����=J(Q��?2�����_��g|�b���23�<�"[?��
����H%���
�8V�Z���0>>N��F���bb�������'&'���'����J��tG%�{�C��s:����U\��muy[�˩T*�
w����r@��c��
��޿}۶�׶��)_q鈴�fѻ�o���[.�9-�كG����ȓ���b�����666b96��b.l�8`�ξ?�r�988��/��f� �s����z���%�<w�Y;>>n}�����,Bq��0������WZ];GG'���k�}描�iow������n�����׿QU��Wi�����?��g�������I�c��7[��ޱl���y:;-)����>	�W�k�؀��ϟ��˗)i�j�i���d�'���O_���)�n��     �a [/9��]��r�^ך9C����X$�u�Dސ=�m˿����������*d�   ,9;5Cc,0�L��Pq�H%��!f�œ��q�W������wM�y�.�XBܠ�3�S����Ѳ�MuQ��xa�]��p\�$O��q
�ezA&nBp�\�%�k��㡗s��;��kJt�V/w���V��ާ>�f�S��˅��3݋�{�N�޶��KK�!� ��`~�\\��2����ߺM׿�qOm'�L�vѵ�lS�՝�7��O?q�ǥ��ɧ���?�ҥK��_����Y*���}��i���+L���K캋&P�p���������~�صq�{����ަ������K�����y����c9>�?ZXX�mpA����~�3z��R�noo�^o��k]�
CpmW����~M���O?��������G]��i�W�v&l�V*�~�|׺�{��i���}{��wR�$�I�^�u�Ν�g9)
a˸X�|�K�"v�"���׬83����      ���5�����`�s�B�6!��H�~��I���/_����݁4�byC�������Y�}��㾎ͮՃݽ�qB��������&���~{�^��%�Jg��[YZ�������cai6bF-����ۋ��)7gb�`�{7�<w�=�οR��r|f�=��L�0����!�g���o��Fǋ���#]_f�`���	g���;ψ�>�trJ#{�{�p�og��}�}��8������O�Ȼ����X_������ܢ���JX�[��i�`s�7$י�������ww�`���~�����$�[��Ī�lSߑI
t�u���#-���)��v��&�G-q��K���n����le�<�.�_gs�vv�8'ׅ�:�t��T}������u+����O�5�+��A�N����v�$/�s�0BǇG�   ������u�۷�*��Wq{�"�~�*E�rex_u�ܫ+{��Q0/����Y`X�D÷�~�P"2h���d�2����.V���7�%x��_�����     d&F2tvvJ�¨ҽ��b�7��V%һ%=T	�8�l�v����%<3�&q����'�&1;����O��{�)�l��əi�˨��c���{��\:���ZY_�ݿ�����������l�̙�w���t,�O�{���[���h4�A��L̜��|����&����6�{��=��e�(�~o�ʰ����~�/�$]���ۺg&Jq��|���~������D8�X�����k����Y�gtt��IX�����7oҏ���ԃF���tx.��_�_��N�(���Z�ӆ����,ig�R�pbp��_�H7q|p������K�?�o�[aB���y���S�����z|G���ќ\�����\ŵ��;��~��׵����l�̶K���������+   ���{�飏�c
�u��]R�k{�����O��݇`ݯk;O~$Ok����]F������_�����+c`hkQ��O����sA�\Ly�
     �!��l���j�;���`$���E�~���$�(o���>|H :ص���L ]\X[��O7   H
L伲�L�߾!��ϭ���{��QK����:��|?�S(7�r���>�[�0c�
�FC��39z�[�4�{ ,�5/����&f'م�t��	����v'ɑ�<x@ :V��Z�uQ4�ݵ�+ٵ�*K�k;;�����ǵ��.��C|O���v�l����	   H
�w��`���lkZGgYQ�\�Uu�ڮ��ӕ�߃�=B���9�
�� B
�q�;��K+X�}��՟��� ��]��ևP      ���8Q�"IP�^�}M����n%)��Z�@m����<�;�� =\����?��   ��p��]�џ��)c�Xl9�����N3IWA�=���m����1@��K<7I�x�R��0��RY��V&�� �p!���F�I}A���?B����g]�\��=b�W��7K�lI�V�ڶ�%�Bpm�I�F.1D���;��Ѻ]D�>��@�o��smw�ݕ�S�ŅEz��	   I㷟��~��?��/�BkĚ����zw�v���k����k�6��ɓ't���X�M`�.�.x������28��\�����Ϛ��       ��2��PYq��g��D�����[�H� ��	·�~K :�ޞ:
#*��7{  �t�~��F��Uk�v9N�~��`���Z6�m�N���������};�ny���"���s�|�l�Ni� ��N�#)$�v��])d�vl�[�j����8������trrB :�W�h�Kx̮���	bpI��W��ծ�z]ۮq��}����v�\Ϗ�~���/��   ��qxxh��k{�mRW���G����γ���
�����G��0���k�"�{[4�0n�>ޏ��[_����      6�z��.�X�����FWlyC�[�3�<�<{��vvvD����t��w>��7n   �4n~s�>����~���}t�Q���+z��5������仺�v�A�.�Zy?�_�_�=.3�*P���= �g�����<\�F��{8J�`�8�c�A&�����)���ܜ]��~D�my�].��zе]V�һ;����.�D)��e�trt��  ���f�_^���ǺH]���'\ۻ�����rt��:��xF X�KF\�a��bǥ�!`%�M���1 	T�J%�-fh��       �`R-[����ۭ���!u��G�7t#���G�D��-.H�ctttD   @���ۣߙ�&�.0�2RX���Çt�ܹ�ЃA<.{.�{�}n���=oH�~~/9�F�� p}1Y�P�D�¨�sV��y��6�뼻�>ѮX�"��
~����A :Vέ��iF��R��,P��N;,wQ��vm�� �k��
ܵ��&��^x����+��W�}N   @R�}�����M�K������z���um燐W�vq�/]��=Bz$�]�?�н�W���u��ޏ7�I�������Y�     P&FX��7s�lI�]s�N����`�����SD�0Zf��(��H�VWi��   �ʻ�oiq~��w�H�B��f��p��@4����&�ܢ����j��7���F<���r�y��8m�{�\���r�(!9-wR�3�C�ca�1_G0�%)�~���cyu���S୓�ƞl�vN
�ѵ��_O��ƶѹ��$>�4� ���x�
����'    ��{ȓ�c�f�T��S�ڮ��k;+����.k�������ݻ�h4Z�3F�"t���e����b]Y�ݳ�]�b��X��T      8g2De�֌���<�=oh�5��$�y���pp��e��kWާ��/   H*�oݦ��G�����})�����ci���_u۷���~�V|Q=@]�74���z��w�昵��L����(�@��'�E�2g��v���.X�*X%�u��v'9����9+t;.��	��ݻG :�W�5�F�\�ۓP�k��пk�D��E��j�Y�h�M��l�_�v���ֱ����E��    ������O~����զ�<M��A�߫�=.�v�peu���g�k>;;;���I.\�k?�����[�N�ʵo�$-��/V	q�n4Si�3K      ��ce�(S�8���.$�ct�
K�,¼ar��9��cai�@z`n��r9��;   ��7�4c,������A�k���
^�.�{;�{�*�L&#5��d4Z� z�K��>��T�"��������*��#2%����W^�xA��)��FL.��مYA�ݫk�U.�׵�o[��X i{�v*]ۉ���v��wm7�.�[�����A   @���ۣ������ۄk���ǣ��������iu�m�xI |�ߍ͞u�����н�M�ݶU��ߺ؏Q#���מ�,��=�(7�5F      ��c*[��b@�J�Nʁ�Z��!��G��k{_�~�Z@4�����ӏ>��7n   �tn5�>��ݺw�@:�}i�lll���>���v�;�W���uD��(u���r}xO�wS�������3 p�|�LUc$���5�\�|��;N��8�$�.�Ӧ`�x�,�,S6c�j�rmw:����g쇀<:���.i�]��k�M��9�n�;��rm'��]�vM5�|�u���c�Ѭ��\Q  /�=�əI:<:�L��R[���z~�&յ�������\�t�y��i(�MJ��ؕ�R5{�]��|^pue�/��)A�     �`�m�)���Ͱ��9��P���t�vٺ���#o!ӳ3-Go��'�����   ���f�����.��P+�����Z��2���?��XD�n�[��c��˻�;�󆤈���eTg3?�PZ���OՒ}zq�E�-P�p�a߾{8*�	�?N :VVW�c�M�]ۉT"x�_�f:�;���.m�\��ݵ�lm��K�v�#��dmĵ]����6���:��_�[7n   0(ܼy����˖��Q��֕{�]a��˵�����[�[[#�=��'E��q�q)#`��������������ͥtrBYm��z�@      @4*%3O�O+޵O��d}�ֳ.yCUB�%��W�� ��d����Ez��   {;;4=5M�������G3�b�^��"{.�j�E�ۋ}z����z�+��~F���9+��ܭ�M3h\��Hp;.lV%?�Z�낌�����E��ڮ~�t-b�vG[a{H��r��؆(\�ݏe������m   6R�Z�t��k�TD�"�v��vym��v~�������ȎW�ʀױ���µ(���7���q�%.� yv��S9zyP'      �`qvzB�\�S�Ж7�&�53?��uI��7L�@y�hYX\$��]��~��&   `P�}�6��������������x�@4<y"��"P�|�P�R�W���k�@6`�R:i�a��
�}�8��Z�J�Q��*Ub[��e!��[$!������-�bj��D���QF�z�M��Y*Z���{pm��%�]�]�n����9�˵]R��&����G������  O����"���I�õ]Z�����˵��M585=E����ٳgtxxH��ӭ׃���q���f�4e}�â]��݉�-���     0Zy�Z����G�vU�[���@uސl���&!o�P�<�ava�@z�6�H�u�'   �J�
�<��0��@ :�`���"C���l�?+���\�^��۫��,�X*�hb$CǕ�����d�����R�0��2:"�.�p���u���Ar]�� �gfh�P��ӵ�#��T��=��i�߮�܏k�ޏk������pm���{-m�b�3��-sls��y�s�6   �ƽ���?~�!m<۰�G���,�O�]���jT��Ы��v����t�&�[���3�������	��lɷ7��;/5s����jv
���zݝ2�e���       ���T�޾d�����������$�����ڦ��c��� ��Q�'������-   ���=������]����4�G�T�T	��Ç�I:z�$
ԃ6�jI���˩���5s��$[a���hm:C�ә;�������T2��u���]b�cX�)�gA�j?HQ���Lm15	�i"C���:��pkm�Yd���(k�`�����W�����g�͵����\�e?{��G�i{{�   �A��՚i�0��pm�ϵ]��z�����˖�]�p��ۅ�f��gQ6���B*T�eX�7C      ��a���k�9��'�ż�8x�y�a��&�7,���a~�i����_��   w�ܡ?����	f�I�4;?Oo�^6��W�����}�g�r�����������zM��*N�q�2�4F��	�}0��SU�𸋋�T�t������#`�6>D͠9�3��".��4����ݵ]�Փ��w�	e��U�����f\!���m�S .�Ώk�c_Q��P{Y��]�$�A�|�N��   T?~BS�S�z�u߂u�u�9���ۧ��c�umW�Ӈ��Gq���*����܌��Q��)�\X��b���su:Z�K��E      �\��}�gQ�������C�P�7�Ǡ�ٺ/^ o!s��҃��l1c   `�`���,$�ibn��0�/]�40�ޏk7�2��BT�o����>�y��\z���m�#T����5P%�P�\�m���"�@,Kb����D��Ғ��[��nWP��|n�K�ڮs۵7�����,>���\��O�ц~]�e�v�����t�"���   ��������O<�ǵ�O��]��{�7"<�v���>���K��f�d���O�J��]��x����_��/��Te2��^)�      #�2�$��]�>�<�yC��}��q�N3s������s��%>_   ��w�hzj�a��
0�P���KNnQ�S''���I5��ݖ;���k��_
��9�R�t�uPT����`�i���%�ݮ�pe���3<H�l��l.G3�ӝWy����������ؕ�f=��Ei��Vc���)����k��NB�*v��� �:�NSܮ�������drtu�e��f�+����   �J�ѠZ�ҵ^8��5�µ=�=�W]ZY�-$�#�ɓ'�׃��}{��]Ӭ��B=Мwb 3P%� �.g����Y��       H<z��I��o�ж�|��yP��ٳg��]s������G���?   0�ܻ{�Ο;Gw�}@`�a� :�LZ2�#P�︖�O��X���m�~��]>P��.[;k�e���}P*7/$�*2.T�]��}v�@)�Q�6KZ��WDa�ťE�d�d(�"o�;��������!��J�v�#ng�I����v�\�.��mm��i����k�}��Nz��3v*w���I���#tt�Q�   ��_����r}8������ܫ+{��k�������k�G��ũ���u����2T�:�A��]�H� d{6;��D�^a�      6P��U"�9C�AL�LS~$O %4���   0�T�U�e!�L��Q�����cᣚ��W��[�4Iʚ�+���)� x7����R9;!܁/f�Y��+T,���[�@V��^7�sJ�#���	�#d~a��$0�v��,�ε�cۉ�#k;�//��f�mD�fەu�cyqm�vJ���x�\�H_}�9   �Kj����r��+w�nR\�E��	D�`�'�|K)L�v�:1.Վ5��!�Px!�!T1�+|}���d��dw      ��b�*�*�9�#:���i��
�ffn�@:8���2   ���=����:�w�
��m�hx��!�j5���`�(P���jQ�7S,��-. ۟�C,�JT�iT�����Y�ʐv�=0e<��0
C6bC�����0	�^a�v&� �0�0'\_N9Q���Q �	�Cqm��k;/.w�������~;E�����   0�{�Z��(󺭼\Z걞�nH���� ����b3��x��yK�"����1�gF�����oT��,b@,����     ���>�E��Ǿ�8.�m�\.���y����K�闿�G   ��Ϟ�'��)mla6�4037K/6����C��ڢ.���A�-�D�$�[u�}{��\�E�.�X���n���=2W�)S񗜶9�u�#��1/R늷���oP(��,P�񁝹���3��g�v�5qs�L�-���xsm'y�I��h�F1��s;��ڮُ���d2tV:%   `X��ݥ+^��f��+pm�����%n�Qp???O�l��u8\G��f8�d97؅�f_��������pE�C��H�       ���(�f���#o��q�@l���	�@:�kj40�  ���~ϲZ�@:��jt���Y����!Pb߬���4��A隽o���d2�L=ޥ��{�L�4;u�G�g���Q�ū�h8V�� ��#��ׯ	D=O�L�J�ݛk���[7kr"m�����zDζk��л�m����7A�v���u��A�_�?���
=z��   �a�իW��s��C�����[�
���˫�>������}��@���a�+D���L��bԕ��{�X�ZG�"��:��l�       �g"_��Ϝ!����˗�czf���3?7G��m   0,���hrb����7�GK?�X��[��c�}p�/���u��@w2��~̱24�O� T�{�@U�h������ �vq�#5��L�;6p��
F��o6��6�`&��z�2�s�3��,�L� ����ڮn�L��ŵ�!n��.���bqm����߾�7   ��Z�Fz���jx����um�S7�v�zn���������{D-H�s�$����|��׉{.]2����+�;      ������n}�v!�}웙�h�����H���������g�   0,<�ؠ��O�_n
��4Z,�Y�D |T:�$��z۷ l�N�]��K��{��O��N�7��V'�p�?�@��#9�JU��$�@[�����~����i��aN+�����K��Ե]!�����Z��&'�õ��v��v�ޝoCԮ���=Q����Q�Z��   ���c�f�T���ٵ]�PO��@\�����[,���-�A |666�ڼwi��]���R����vW��U������~�/0��V=k�N       �d����GbyC op�L����e   ��R�D�㈳����Y�z	�{�2�8.�{/������~"��u��]�.�sČ�
�6 p��vfKB��u��dImQȫ�0�D��}��������?N ��;�:Rn�k�W�s�ۮ�s/�k�ŵ�&��ӵ�s��bq�2�v"i�bwj��]������ŵ]<�񾍏��λ   ��{w��ǿ�)m�~m+ϵ]R
�vO�Tu��KK��������imm����s��$,�H�Vq��`�����rvz�|��f�      $�z��U��=oh�)�7�o6�ߋ/D������T+   ��ѠL&C��#nff��3=E�q�y�$�_�z\�X��5�����(h7�|���Yy�D��x�rVrMD3D76���l�N<�2!`�g�F]���-1��v�*`�vC�M�2޵�] ޏk�&�N�v��P~��]۹#+�Wtm�&n�ʺ����[�_�˿   0l�)��h����~]��ԍڵ�K=U]u[=��#���-�3A0w�s��%^�ľm"waq��U��X�ʥ���h_X�}����S�     H:,o�D3*�5����߼yC ����^�B�>"   `�x�t�ί�ӳ0Vvf0032؀㓓����Z7I��^���%�vu��9K�)tw���K��f~����{����T�tq���m\r^�<bB��gs���g_�̍D���\(��ium7��RGP�+�k�̧k�Cl���L�f   F*g�t�um�ֶ�\�=�S���v�C=U�z0R(����ku����n�0���7+s\���<���o܌��z� >C+�     �t�G4�T*T,�[�7v�,o��ؙ���=�..Ӄ�w   6�={F?�� pO�s3��Z�ҫW��>��_/�64�|ܾ����f=���%�����N)��TO�������d���P]`D$<�A*�%�y��2IN����ׄ0�̈́A����&�㻝���8e�j�"!���7�v���7�"uQ��pm�0���ŵ�^o��j��m_���|t��S��"u[�I��aS��5�p���"��õ��@V���4O����~D'k�ݛǋ���{��繳ABq}���޳c�}�����ٱ�����7��\�� ���8���Ϩ01FG��B�d[*�E}����תUr#�v�_s�۷k����F�}��Jɵ]dna�޽y�}�2�nWX�x�sn�"͊^�ZdbT�D)�h�[��x>;
�      I�L���{��yC!�����}�~��@4
-�H4  `Ha��ls8 x�'&(��6
X�mss�%pw����_��҄��κ�Z���-oHB<������4����t���Kc�N��g��"�E<��'��������靤����[�A���ߧW��,���&�q;���)�x��V&
��m�ʚ�b޵�x���KOُ!ݝD�-)pEl��Q[�vx�O�9��q<�Q�|!�M�T��٥G�;���qzF�ǖH�0M�λzx�MNNѷ7����E�������v3y||�=L�W.�[#��������M��={�Y�5��
�<�����󑑑�oN�y��c�yq�γc��I��e�io߾�>��v�w�+}|�~J����1o߼�k�~���������޾�K0���.��P�^�}vo�g����U�0R��ޞ��U�.��}xTΎ��'����bF?߶�>�.��[&�po      �����'ޝ��{�yCqP,�ۭ�c���E���J\1T�s�������Ўͮ���i��p����;0f�����Yl�^�T�����O�OЍ������Ȏ��QO��,�:�qǔ%��]��}��g�+���B�y�,R*�b;�ql����8�{v���q�ާ�3��޹}�ʧ���#*���g���]L�g�,�7����ǚ���z�;/�{{C�������e�2x�E�9��p�����{i+�Ms,� yQ�̖���;Ӆi�.��´��N��ET�*��
�`#~NOO)H�{�>��~0��k�7N<n�~僫�އ��]������j�k�y����������ݵ�VOӅO��l������7��+�폓ҵ�ٮ^]��:�&����9��e?���w����d��O>��^�����������`�*���-��8`�����c96�������R,�g����u���{�:���gc�B5�s����3366F���?�sg�Y�4�����-,,�(��g�VL�o|�����������D쾕����~�S��]۝��r���;��t|՞�U��o��X��_[_�p�n��W/��������3��[�t��4�~�kj�^P��5aiו��+�kj�I�3u��      �b���c��x]��&R���8o��_AC��@�"��{lb��Lx�R�2-P��p=����1;�i����_:�=�6R���!?~�����q��yO�{o�"�y�����q�Ń����W��t��z��atǏ�w>����x��&��p� �{k�1I��Pͬf�/�ܢ�ҳ�4iRѩ�������|�;_G�O�I�u6���D�Au��nIj#H�����N*����X���^����K�0;;�zE�2���f�Qfsm7�qmS�-�1���gB"�fu5�Q&k��Z���m��u"idBr��$�Y?r�:��M���&n����6�T�Vy3   I�%��N,<
��"x?������'"�z����ա���Odn~�@40�;�b�ȓdw�^�W���uDq�:X�P�{�ә�T<D      ��ԩ&����H�'����F$�y��ϟ>c*s2�kV�o����}va��C6�9���*�NK4>5Ic1��ۍ��˥��߽�:���ޣ�Ϟ���hd�g�LOOOS\�y|#n�����3'if ��� �sg��l悸���দ�bsp��g�t&r�g>z����׮���w�?������L�����D��X3�s�s����pp���n���E�9X�E�Π�_�؇mˆ�~��O1���_�s�rog@��y�R���X�$`e<e�"w�rIoQ���[T���LZ0�m_/^� 3�3�6��mN���B�Q�M �ߵݱ/�k���l(߆ \�u������k;9��Vh�����)��@�N�=    ��g�ra�vv����wmW�k���Q�����������{�U vvvZ����Ůu��+E�
GgN��)��Ur���(����A�     @�ayC�K��Wn�ٶ��^��8 ֶV� (&cāh`�-�L�   ?�z���3=3C �6,NZn�-%���mP;_�ꟛ��5C�u����R�� �tI��u��mT�#%��f	Te�vˉ���`]�n��Nr0�딅'''�)-@�L�~�;�o-@�v~?*�� Ж���rm7��6D�ڮ�ֱ�o��������'   ;t���t�>\ˣ��k{߂����Gh�Ph�@�4z��-,,�*0�mZI��c��y��S���.�Z�	�!&       �d�e���q��.T�۝yC�����2��г��B[�^   0����������^p�lf-6;�1�[�.�����w�+G����r�bސ�+����y�d�4�\�����2Ή�(�/ޮ(V!}nM�0e�۷o9m�02>1N��QS	޹Z�x�[_��ߵ��Cǵ]"ZW�Br�%&��m7?NѸ�������sg�ѵ�:?vv����,}��o   ;�����U�ݟ�]V?R�v����}
��
A�.��=ө�������AP�0�V�l]s����ɬmV�b���x����D��c=D
      �?j���^�\��'�|����v黤8o�^�j5��F��������W���   �a���'t��З��^�&�)���R����o�O�C�s���]b��=�\K�to��g��3?)M@����Y�Q�R%��N�=�2����R%!��7oބz`137�k;9�um�H�.�!:�v~ �p�����	�H�o_���{�	��k���&   ��Պ�u�]ەM0�v���1Ѱ��@} ��blJ&t��Z�{�ʸ�w��f��K�0�]�E�vO�'      �T�ʔ�f��Xƣ����;�ud3@�����O���D���/�@!7�r�   �6�Dq��p��Hl�&�?��ڢ���ĘW���/�$�vY���
�X��!�4~`>
��r����'���:x##���,H�)pqb\�T*n���IF����G ���;�'w���~]��u����~��{um'�ߢ�]-R�	�[?|����nP�P��]�   3o߼���q:>9	ŵ]I�޿�<�v���꺝�1��w�ޅ�_=���΍��ҊHkk�6|__��2��]Öٱ,�b�*      I���Z3�es9ǀU�Y��A�D|��ڷל��_� o�095E �h  @���^*)���n�XI�����m"w5�Fg�n�%�%�W�~�r�[f�Ŗ�1%@�Ѭyqے������X�2هA���`�;;;�����	�Crm��J���۵��J��N!��q^-�]�Y����+�H�]?��d��G����   i��Ç��?�1�H�µ�뱒��η`��`S�� U��S+�]�Rv����A�|�S��;1�g
�     �T�3ds]ScY�B�@�7�	�S�7k�5p295I`�-����   i�tF��Q*���9M��A$�9�s��r�gc;�L�k��8Ck��B����c���O�Ƴ�ո�3ɓ�ݝ:��qg��F|�(C�*:����t��Џk{�����n����$
�em̵�l�µ]*��m��������O	   HGGG��e�R��{��_]?݁ \�yFG���7o���f�T���:}s׬];���*��C���w"�;      Ief�y�^�;�1�I�N��3���ʺ8����Z�5o�T����F�����fq~��>yB   @Z`�{�_���%0�����=*T������Ͼ�9D��z���ܡ3o���"�͏e pj���j���]l*�6��V�2+JV��ۭ���{P�ޘ���
ăpm�]��P�յ��/��֕�v��i��������.��rm��'������4�R�D   @���+�+��{=�/�}߂u�u�ۏ�(��P����|\lmm�?IP��Jˮ�x��0Es��֮',/)�B�     @R�.4��+vc,�l�g���]���l�לagI0Ȋ#o���[�0��������O   @Z`��^��;�9#ܣ����`�-e��&M*�f~��yC�v6S,��,���j@��ɑ��̛��rY���27epJ���3X��=h p���q�Eꌨ\�u����T�n4�^f\ޢ�]���\����|��J�е��#�Q��  @�`.��|��ժc]�N�pm����{=���~���4����ׯ_������u�w����U"ws��H�&FL�z��`U;� �!��n�#Z��CU      I����IgA�.KP��^������ڍ1s��5q���;�~)���q8�?��    a��v��I�u&u���kn����|��*����iw����ĳč����mIl�A*պ������-�@>c��Ϗ�ir��rm�������2lr���vq_����gLW��]�p���n�K����N�յݠX��Y�F�  �.=|H}ﻴ�%@Csm��=���	˵]�:;7�{�����ŋcmG��y�S"?�]��q����(s}�iu��     �dR�4�ݱ�bsI�� ��;�<�ob�l��fz��$����o[�RA�0"F�E��!%f�߷V�   �6�:fr����y���?c��l6�z��U��Vi�5��7�����yC��\�n7��Z��4�^�O
Z���+tuq�'�5�zc���8��b���u���c���!>3�3���k��˵ݱ/_��6xi�b_��b{Tۅ��n�Y^\���}ZZZ"    M���4�}2ҟC�ڮ�
�l�nR\��z3�D�	D �L]�pa�T"Ҁ�!l������j����}68n]�%��      Hy�F�1���>��K�����.��+�����Ak�319I`�Y?�FO�?���Q   ���˗���J/67	/�0Ɗ �3<99�����u�,~w�[j���f~V�myCu��܂���V��� p�I��wS�ncOb��m�|e�m�R��~�{{�f����𙞙�<��~\�u�k;_��=7����Ե�YG(s��7��A4�}�]���Um�~�&�ƨT*   �6�=J�Vϵ]V�g]��{?W��lzz�@������n�:����$�+Y�S:�T�-��J��H      ��mԬ{x�'��O��i��yC��;�K_�[7J��!����	����<}s��   Rǋ/�~���9�S�G�u2����q��m�*rW���{���e��|�8���[�ȥG���3�L���w�ywpo?'�l2+I�4԰/��G��sb��q����� �m�k;2��3O��d���N⾽����	ǳ�K�-��V�'z�Q    LjoS��k{?�p�v]�g�aӏ[^�T"FL��C��enD���w+>``�͛�h��2      ��Vo���!���6��u�o���sW�O�,7��C0�:�����a&�e�y  �J��*�s�L;��(���w���ի�0������7�q�g+o(����F9�`q��|���L�9�yubhc�L5�B�j�7G��i_���m���#���a7��2�v���pm���\�M�w���2�z˵]�_IYK�b���"rm7D�e�j�   ��rvV�\6G����P�S��^(��Q���'n����31g������TB��:i�]��k�d�pbw.PU)�       �Ԫe�}�Ù]��n�l��=j�~�chk��i���7��h��'0�@�   ��gp���lTt��m~6-�µݹ�\+l���3?ט�==3?C��Z��z4�N.�v�4��Yg�����~?�I���@Ut�@�Z�.X�tm'��Q�v[|��K��:���n	Qt�v$�G�MR�z�v/m�(��R��   ��勗t��y�~�α��A�۽���\u�;>�{d�)�t�;@V�Kf��:�*Peݫk�x���ئSΦw/htRF�     ��Q��)#1�j?�r�\��&n�d��F��a�0Ɗ�����%�ɴ�   @Z��|f3^p?���_�����>le�6U�L�7Eiw��@s~�"n�<��Vr�O�*����񉎮H�S"�ٵ]D�"tm'��D$�۵]�˶�ͭ�"/��q{�6q��F���9���$    ��|������]A��k{�'��f��RE]YMi�Iq�H�\��5�Z6������V�n��[E�蕲/	TA*2��f]{�J6c{�0���2�m      �D.CT���PuTU��I�X�^��=g����-b�^���7�cp�f�����6   ie�y_9;3C�
C0����=2���"������� ��Frl���s��kYB�x4���"$R����ו�-�@UX�#P�v�@|8\۹�+�X�
޵��Nׄ2_��n�v��r�=�n�o~�   i�\.S&c����ڮn� ���+��ӵ]R455�
J�p�KM��6ʴ�RפS:gg��a�1�%,�p�1@��S`��#      H��l�Q�p6����mV*\ڇ���=Y&a����	��^�� ^έ��7���   ���js��]\��}����=*T���ͯ�B�*T�5g��ߙ�k�:��htRI�������Ӆ�=���`�9�ɦp��T%�m����86F�\�+q
����D�2�k;WOx���zw[���+�N�筝���nַ]���n�x�~\��c����k    R��ݏ�յ�_q� ���u�g�!p� 6�*��
~{~�h�D��b2��!l�����=p�\�x      ���"�p��y�}�tJq3�o����	Ⱥ6��v��ä�_�c�h-�R&�!0�������   ����+���'��|>O��<U+U႙���g~��ڟ�f~feS��T� p��T�y�4�y�t�:�)��T���QQ<r4�����!>����gN�z(��2q{d��rq�%V���+qmo�R&@?�����;�C}���u��   i���=���õ=q{���:Wsbj�@�looS�R���QFTZv�=q�8���8����o��o�:      ��D�y�^�f^����,��|���O�$��V*r����������#�    ݴĭ�v_[�����A��R�&{��Y��r����#�����c��Q�'��`�#A�]��
D��TVY��d���'�h�� �������=��KD�Ra;_dkC8���l������zsm'�����)\�%mj��1j   p�9{��tZ*�^�k��v�k;�����9::���cO��u`P�]�ޮ�8�,�z�`�,�0�m       Y������Q�ԃZ;6m�}�#�y��8��35}����̸`�H(�C�>�@�   �$
��0ּ�=܇�=l���R7��-��ʌ����KA���^�5�@�x��J@��u�A[�N��O��:ʰ���#�۷o	����d��h�qg������/�v�p}�]���"���   �v^�xA}�ݖ��_��JDޏ��o�vV��0���`�� |�����#� W������*:U�p���`�Hw      ��h��4�o����f�0�U��6� ��Y�)c��W������16>N`xay�ӓS   �N�Z�|.G�Z��pR�}m0}g�f~v�˶w��1 �-�`�5h��iw�欋̼H�ܕm��t�J������+ ��	É!��ο�z���+µ���ί'nwݦ�v���PG��nqqv���{�   ���:�86ޟ�9\��u��tmW�B)�o.�p�
э��pW�N�n��+��m�K�U�s.֐3�J      ��P�ڍ�x��^����/h�P'���+��!�� >�&��˹�U�z��   ���zk������M��f&�6����i*g~�*t��r]�|68Q�\�@�$ZS�{wpo��4��*[R��s��~��wmפ�r��y!���Nr'ٵݾ�ו����Nܱ'���ݻw   ��F��ZlD*"���o���������"������!P)]ܻٻ�����\p�Mܮpp�Q��      Y�5���;?PULL�5;�~K�P� ZM�7�q�����7b?�;�1�W���E��G   ����-��{߅�}�-��xa�m���Ѱ�w�g�Z�Ϯ�tup��XȦ�o��F2�K���GY��ic3�kk�H^�0������TED�8&��ڮqE6�v�흝��u܅��xum��-��k;�_�T�U    Q�w��k{���u#vm(���!*،[i��� n競�VĪ�`=��� f��@�     @��i������J�sי���FS$�%�H�	�888 5�l�!    M����(�{���(�Q��kI��9��I�X��ֿ���0�$17���=�?� ;�߁*S|��bN�U����T*�6b�6tC"v�����yumׅ��(�䡻��N'���tmw�����n߮3�E�7G��
b{r�Q*��|�4�u   @�z���\!y��KǊԉ�O�x\��6a
��`��^�=��+q���BA�.	�����      $��^wܿ��V���0�}�[ZPQ)�.R̯��
�Q(��	   ����h*��=:�`��:�b�(rW�����G��{�X�0Ki wd�nsTk?���@����TE�hK�����.��kB-R�	�ܵ����ڮ�_���   ��ĝ(�vy��tm��"*�v~E6����U��2ȁ*�y#&e���U��*���+b	�:n����      H�������A�>�~)5�B�0:�1b0�:    R�����8n��̳|�����f��-o��4��l}&E�s p�T1����c�M�#
�)`�v��]������]�S/��O�MH�y�;���(t�H���7I��]�5�u�9�   ��κؼ�)��;��ȣsm�'��n���"��T)����ciybL�j�s��vmK���&�Y�������      HZ�2���߭�b�Ј�;M�4IA܏t���ӏy�I
� ��F��>�@�   X�wq�����HKͦg�,nw��+o(�se|��=6X�0��t�ePp�ii	T����{40��\>'�����*n�^�Jq���.n���������}��!�wm7���l�Qr   @�x��]�z�N�$��pm�Y7^�vU���c���{�Q	K`/ƨ�AT���
w��=�`�����
�      $�F�b&�����;$�:�DY�Q�c��ݹ�7���h!��A�
*��	    m�ad&��FƑ�H.�k-�f��~�kq�g���l٬���5����{,�����sMC���^��"e���&�m��|>�������l6� ��b��>|Dַ� �v<S`)Ĺ}��v�wg�=xh+SȦ��o��f/h�tpЪw����M%��\��vک���C��3�m�tyc\\�e������Sz��M��9m�z������*�J��1�<�j�J�r9��f&@���q��� ��z�y�q���e��q�;���8�o��z+I����١��#�q����U��w��t��ݞ�W�%O0a���;�>õ�g��tg���q�k���ޛ�I��g�/�̳���>���[rK�|���w����iw�[�ǲ{,�#�j��ե�+���Ȍ�8�	F�@�#H�A>_);3 @F1"��}����,�fξ̺�C6���?��;��q�˹Ee��p8����7���_���!d<�"      @��N;?��Hu��zᬼ�3���W%Ņ��6�.�9����}�\֙۷>�Ã   ���#���G�׿A=a.�,�	�E��s�M��r��`]U;4���y�:oȷ�O�� p��lqc��tO������lR��	2�M0��+Q뛉M\��oa�7n�ѣ?�@)$+�=I���I)��W,l��Z<���ӧ	Gt��\�SOc���x�v?(�{�����,�'T�	�}���z����Ŷu���O?�E_�{������Y td0���۷�L�y��M��zN�g�~��'}����z���յ��	}ٽ�w=)ux��wg�|ϳq[D�~\��ڙ�����}��[6�p�������w~�w���p%�����OON��gOu���]W��>�}r|LO�>�4VwxW�����^��w���������>|�������M\�-�(�Y���s�A>eL�=E�p��x���q����!�j�!      �g:+���aX/��In9g��t6�ڥ�,�-6���ަ�p��`0c ��������ܟ������~rx��5����N΂ݮ]prtl���8:��� ����췫��-=��\��7c���#1e�_�И����kg�yv�̐�,���}W�L._{��3�&W��������>o߿O������q������a�����X�~������k���%ɇˇ�﫸+R�s���z�͎���%�������������9�2A����$vpWݘ��hɁ*�q2i7?�_�@[�Sf0���*X���us�?�����7�)Ru�//)���_L�B<�/�:m���H�õ����:e{f/��P�u/��긄�]!$_���r��m�;�Qt�{A�׈kG�K�/=�����ݻ���AD8Ha"'���� �\����U�L��^{W������\�&\����fT�=����>o\�ۇ}�
к|����H���q������g[�� ������L������h{G���3f7��y��������8H4����:�n�z��Hro]����.�i�y^�v�p�Fܾj�e���i����;�]���6]M���      @�_σ�\<L2�b~���9!d7�&ʪ��(&L*[�Jx��]��p�.=���V�~��7��ӏ�o_��ݛ{Q\�6Lxe����?�3����qGe�����ٳg�
�����̙��������Ύ��8]^;X�{��=z���/_�7,����}���ݻw��������l�����~�?����|���W��{�����1��o����}k}3����F�"e�y��d��]ܣ2}���q�_�/�^�+����)@���ٌ%��7�|S����nX��+8A�l�%q�Gf��B=^����~�X/\��~j�X�n���ɣ����~��Jr�K�Ƶ��P�N*�����}e������"   �'ؙiIyZm���
���3�V�r�pm��s���I�@g�E5�
���E�"w�=�y^��k.D/��      P������O�$s��NɹAZ:\�$t7�ra����\����Ϯ�a   �,��>�?�yC;,3_�onQDm�ū�9=�p��7 �'cw��m��h&,yߞ�db�Y�̎��*��-*U�����ȹ@*/ZH��tmO
Г�<��~FQ���Ke)���9������]��O�S^����F�ΘM�   d����x����YaѮ�i��ڞU�l�v�n�7Uv`w��
�]SN�L�?�i�A�n0���ۅ����vgM      4��`�<?1v�I��_��>g('���椬ݙ�yC;�;!�����}   �t��Xk:=7��7�u����[��u�U��0�=e�7d����kN52�k �!��)u;�L7~�E,�M:1��?
vbX�@���9��	@���.�M�;b�Q�k� $�����.���J��Q����e��     �o���U]۵*v��+������ʇ�ט����&Փd`�K�'��xu�8fO�x^<A��;pp     �:lt��x^��3�5�k/>�����DE��?ߟL&��:]�    �0�PS��Ev`�X�`|]�՗Co��7Ê��۹8���6o�S��Ѱ�@�G�[$�c��7eRԮz.�L	N� �b[�_\\(�n�oϵ�Br&�D
A�\پ�k��<Ȟk{$�����?�6�   @����;� 9*�v�k�%X/ŵ]����H�ڀ�3����e֭���g����v��EU�굪�       �K�෗H2�P�?V/xU�N������bwg,�srrB�|  �9�   I<���L�V`�ټ���Dus�zq�X��;�tbɰ'��{�+z��m�pR] �lrND��v"��H\�V��H�^d��	�///	�O�� ��I��um���]���Ūk���^)R/��]#�O�rm��-|�gT   2�g��ߠ�I�cP1���������um��E�[P&��`8�:�L+ͬ=�<17��uΎ^\!��P���=      Ua�s=J�qIgE�O���H=P��0w��H��vC�� �w    	�kM���6`F���6fչE3q{��n�z��>�ƹ�TS,.o����,W p7d�+�����I�%��X
TUiBw{���e���D�Zq�,l�D�NH.���ޑ���vŻE8G���z=�um��^��t�   ����)���s�;\��ߵ����5F�Q���mbr���R�*���)�G���     @e�D�U�<�y݋�s������3�VӘ ���!(��k���/�ì    ���z��n�1ެ)�>Ʒ6`:O��s}�'n�ŪDQ/�����yCw �n��n��	Qn-�V)+,<$�e��n�^#sGB��/O+�V��5BvI�>���ubm{�풐��wm[ԞS���b�D	q���f�O���     28?�~�W�k�����!nw�ڮ�[����E"�E8�7C ���"����>/�;��,J     �����bWpE̞C��x����ԨJ3([�Y벃X@\��lmmqQ    �紵�Ig���%�ځi=�1���nf�Us�U�-�z��Q��;G�!��\��7�8Yn���W���� �i;t��V�� ;͵�����'���'�*A|)��A=Q��[v$�]ң�u���5��	�u��^'�7tm�w/
�766���   @�- S�Q��ڮm���i3�C>�����m�)3�e��ֽ칽b�<��'��ږv��x��      @�t[�|	{ ��Lɼ�j��dy6i՗�Uiw�4 p��*�eg{�X   �������{M���ln����2�E]�д��a��X<F�7\����^��i.p/̉�<�T�[�V�+����\����RYȭwmOuW'o!���u��1���K��<��|��E�9Iu���K*���    l��^��/���Zy\�]����"Z�����x<��#��x I���"��%��bt!p     �2������S������ �����t!�+ۛ��pL    �h{o�@=�$r ,��䪸��$�T���H��z�"q����3���k/V?�&N)��e���U�`_� ��E�E���Y$��k;�k.�v�pޞk�X�ͯ��������+L  ��ٌ�er2���4'q��pm״��k͒���O��{�X!Y��E�	���q��      *���RZΐ�G���&S�u�]��d��%ǹ�;���Lc,    	�~���>�z��4D\��yk]s�&g�(D���ý�v3�Ș�����
O�
Ik� ��{���:mYQ�L%�����.<��vw��i��������ڞ&��w�T   �@�n�ڮy��9�!n׾�>u:]�e�%p_�����\��
��EnR��b�ߦ      �A��Gۂ�����k�������zTU��=�1lW<PO666
   u��j���ԓv�X[TA��2�-c��?�_����o?tz�T8�Z$x�խ��ڎ\s���!L���	�x�v����r������4��I�{��|)�v�r��/?�������e�vA_   @���]du�v��]ە��uqm����VSq;N]l�m���5�b)4��H3 �a4c�����g[��6�      T��������T�+}�b*nϢ
�U�B��
,�T��`%��e>   ��a�u;]��wk�aޖ�[̓3̚Wy�~�/���e܁��݆�����|ERz�w�V��/O,�0>�E�����]�)w�um���ʶ]۽�v�sZ��]�P�k{t��%�)   >'po�k���������"�^�@�4z�f�J���C$�)�W?�      @shyB�c����K����z�1�
�%+�p���:po�7�%    @u��dmas�V��4?ły[Z.��M�5=e� y���t�f�������)�X��� [ʧ91Į��{i�v�q�F�v�@�N����v�S7wm׋�m�e
���/����u���ή0�v�3   @�l6�^ݵݼ��uӺ�]ۍ�I�f���<�]�@� P���y~R���!�     @eh]�ϧ�'t;?{&s�7�C�    4��:�ƹ3�J'k�V��˕G09Ts��ɝ�cu�TCZ|rY�h���Q�د��.Uv�;[.��j��\���R#���+�����q��k��J��TG8�?!\OI�b/��׵=!�   ��l%q;\�+�ڮ?�N[I�`�y�Z���A8?@�0�+��Қ      �CN<��{��9A��Oe�#�����    @��\�sǘR�N��u�-Ff׺���_�V�924�?�Ғo�7KB�jt�z���\;���c��ڵ]U��k{F�+��/Z�����t�,���ڮoW>&�k{���3    �!}O�ھ����v3q{���Δ��qm���nl�hNr�Aq���K�{�'     P!�8��:�񥌄�v�d}�����`�e�N�Z�#�    h��d�ic�k��tJu'�+� ��(M�/ĩF�D���]x�d��E�J�g,� )`�f+M�!+P��z�^t����5b�Rn��*��+�W���/�s"�\�iQ0_�k;�<a�   ���k�ڮ��޵}!!��Rq�cVp���� ģr��k��{y�      �J8���a����~�7���>w    -�'�ƹv���ݕ�ܧ���7��e ��	X���w����j�Jsm�R\�%��R��j���T�k;Ie�Ӣ�w����    J��ܕ��S�6=CL��󺪚帶�z�E���u=�E�|0o�F��NiE�Ųi�      nH찔7�'��6�n��ua��3    @�x��`�g;4:ohl�%�I�F�����.6�s�^C��D[GJ<����5H�H�A(a���=�H]S��?���I�r������uumW֡�\���|�#   @�j���k{ �^cq{^�vS������|����y�V�K��-6ҭ��U�     P�Ni��ZVN�@f���ÝYoW      �y[:iW�Д���⑿|��3.�nv xv`�Y���]��e��(��M]ۓ���,�v/���sm׉�^x�b_�k{R�ηS�k{�>bT   @*�Ʉ:�6M[�5Ƶ]�ĺ���k�O�>��Eշ�>��f'�dm�     �
��3P3V1�B����f     P?`�e�ۊE4�V����Z��!ѭ�%�j���s��}��m��l^�k;�(-�۹���%%w(l�_µ�����>�ye;庶׎�   �e6��_%��!�^]����B��d�qx�\�yZm�l�T��^-�[�r��     P��s���OJ'���m��Z<X`m�C<     �c�a�{�r��"h�!p<e"�zcV]@�@���\�M��Q�%�v�NX�.��-3���   �c:����pm�q^���pmO�� �0o��JK�1�     �2���sO)c���1p      ,&_Vh�-���I�����E�B+͸�!p7f�L2�U��C�k�v�-:��ھ����	�b�L�v�ڎoE�B����*��2���c?�b���+�����Q[r!    x�[p���k�Yai���4oXQw5�v�Nvhb���;˰!���      T�<��RWc6�����    @�h�0#��m��l/�O�F��8�t>�X�t�h��]�c��\�.�U�k{|J
���?}��k]�=�A!��T�k{,n'",   ��0���祮盾�e���`Km+ PU,�;`|     @u�R�˴c���6S�.ͩ0��vī9�+    z�=Yk<���y�Er�Ư/���]��g�V�]�k�T��ڞ��k{xNĻ�S�Kqm�����pm�1�   ��f>��#Sq{u]��륹��XP�k;_	Y;`a2      ��x� �M0���)��2    |O�*���F�O����!p7��Ce���̵Ԛk�,Ҷ���I='*��]�vV�+޵=)�O;'    Ȱ	���1Wwm/���L�^�v����R����VN6@�*/�     P��(�>Vh�ٲ��Z-�M�   �`�Yg�X����H���Mi��P��b���^�k{R�mѵ]�/�'i���Zյ]QV�k;��   ����攛d�µ}q{����r\�źH�١�n�      ��G$�&JX�uma�3    ��xX�l���Ҕ�� p7��Cu����ϾX��V�n��NI�5'$W���"ɑ<�k{xNJ�}R .��+�'յ],Ksm_�it�j���<n	�v��    5��۟LVvm�S��庶���w      @S�@?(�?� �����F��G   ��k��v���.M��A�n��1��}�@�n���ݡE��=N���k{�%=͵=)�����	ι:B_�t�'�NQ��r����.~�,��>_}�8   ��m�<�%��k�ھB�"\�5��>�"��g>U6���X2ߓ�     P0>�
柖@
��9a��    =��,��m���M wc��!$�*>/��v����[z�>X������y��>�L�g?���I-����5(R�ˇzRm���{�O��O?=�w��,J�K.8?;~�y�J(O��g��� ]כWo���cv[�z�L��.���c�bg��?.<}rr�(��`0���sg���驳k�����Ņ��ٵO�Sg�.����ap��\���]���w�}�~\�����}�M&'����{�._{�Y7��>oٿ�p|Eak�<��d���7�����r͕��s���o���n��n����k�����zZ�Z����ѿ��E��NNi{{�l������}^U��2)lJoؐX��*      ��vI�ņ�V`�&W���*;���wO_[���f`�ߘ��8�w'z���b�;��*�\����.�	�]���!� ���3����.m�m��!e}�5u�b��B�\L���.`_&����t�x�[;������k�S���#��k��~���;�ߨ��r����K\��/����E�U�um��?|N�'̟�b逮��}����}��	����+Ta��gϞ�޼yC�nݢ~���o���ٵ3�%�޻w�I�/^���O��+\�w����{��{.py����mmmY��v����۷���'��~���ܹ�lq��מ��������������Q��U�k;����~F��\�Y���wS����~�&�	=x�P8'�V����?��E��g����Ee����`n|��A�     ��0�rɘK�Źʎ3�\��n���C��l<�_��j���prt��%np>�������k��}����q` 2?.`F),�
f���5wi���w�?�ײ�+C6�A,�r�WWWN�g�;뻉�L���\��l��L��=wtt�Y��+�~��B�gc��_~M�p�����NzG�q6��ݟά��=�Ɩ^M�=�p����$�?9�Cl�fC򆸫�ܝ�d::M�R�Tܦ�+<�o@��7���䲰]/$_Ԏ=�>��ۓ�m�2~�\�u(QG8'��Rl??���^)$׉֥2_ѷ����e\;-\�)�^���	ۅ��#   @K��"6+L�nV�L����fuu��!n״iz^�^�vq���-(�C�ơ��K��f��      Tѥ'��;C��ĥ1V(4q%:�}��}��O�����o���޾|\��+��/�������S��_�u����������&v�裏��s�U�̜�����������w����>���M.pm�Ča=z���/_�7�.۸|��w,[\p��]'�7ِ-���_������������3c�*����[�f��;��X����湵�>˝mll�8v5?��9�HB�n�J+|�B����S�����^3um7�k\�=R	瓎��]�9��\'l���B�%��'������r���:    H��ti<��]]���*X7����Nʺ�\�՗5/�A%`WɈ��X��0P��0�     �:,3>��0]]
�m�     ��Hl�U�mkm�U���6���5�	��7�p3�Q��(�P)����lʜ-�tmWG��k�(�(ߵ]<�pݒk�J�_�k{�1    ��Zfߓ�\����uum'��*˵�o����n�u���?V��xF�#� ��=      �A;3Α�NoI����V�-b��f���Y     ����Z�{�'�b���!z�����ԃ<;�/pY���k�(ZW���K��S�Ϊ���1wm�w�+���'������4�   � �{����f�;��\ۥ�q0ٲ�m�ķ�/�J������       G�q\C���������   �L���09�D
0�>�#T���		��e�q~Z-����7R�l�0�*;��W���wm���C�rٍ0�I~i�vE^Y��+]�5.��)��
��
���9)�Ay    (��E�smW>������0\Wעk���ނk;_w2(��*gcނ���Z���      �Qχ����G�ik[A��0�aG�Z��!    ��q�=o3��/gl������k�,g��Sz|K'�?Y�B�k��xBŹ�3�O��.	�=OZ@dٵ]hWю�k��^�k;	�H|���Ν7�G   �������3���ZŻ�ӏ����ڮ(]O�q.(���������ߓ�Bz��     ����}2�:$���`�,�;�0�N	Ԙ&�   �e�x��L1εB��������7v����=��C�n�LvL�U�N���:eͳ���@��%P>㫫x�fŵ}Ѩ�	[��Ȯ�|��]�e�k{� >Y�_.��k{Z���Z�y    Ĵ��I��++j���}�z��tuM��Tw2�������z��{�틇p�^��Gm�k��     P3���9���s��C�R��"����?5a    4���\T]�^Dnr�i�<���9uÜa�c������!�@���UR&7xx��Y�ދ� p�T�>۟�e&$_ŵ=<�+[Ƶ�?Gc�v��X�k�HP��vR|�*�a�V�   Z<o�=��k��0���"\�M��Uwm���ʧ��0'{�/�3$����     �����)Ɣc)51X��!yC;La      j�t�q�ʞ�U�<+3�g�?�:������	���{���ү��Upi�P��Ɍ:�Va����K~�z��3]�I�Zn���yU_tK����*�rmO�7���۵�{�Ն�   ��j��yWum��4���k�I��u�]۵���w+4z�f���ew�<�YE}�<      T6>���YJ,�������ք�s�=��0��e��W    ��k�������%�̮3��ɔbv~q�"���!��;bSQ��Lb�&���mHuh=)"����	�a2�P�;�((׵=n[)nW�ծ�|l�ڞ!Z��ڞ���������2S����Uuf3?<\]]    DB�,�ھ>��|]l�m������`� ��ח��!�     @e�r��,S,��s����S�r�=%� gK     PG�7�Cּ������+�Қ�)v���x=	wc���@�N,��Z'���[�*r_�a���A������.ѵ]�6/���ڞ}>*��T���]ۃ�|^�"]ۥ@��j|E����   
�&�pm/I�_�k��x����T>Х�p��ȡ*��|��=!�0gF       �L���m� �fMZ�	�?&��f���Q�V�`�-   �D�Ŗ��l6~@��a޶jn2���Y9q�� g(�9n�m��!WS?vXX������aC�[���L&I!����	q���8��F���ڮ�K���Ο�ޑ��v��j<���:::"    ĴZ���Utmן�y�����L��A�|�U���H�[^�M�     `���@�sR��!���3����s��L�v�?Y�3��LgSj��p0   $677�rxI��`�c�*����M���l.��F>s�gn�;�5#��!���P�xnm���U
9�
�1�{n� ��ڞ&n�]ۥ::���̢Cu������w�X�F���FW#���%    ��NF��'pm_7�v�Jv��E��=D��{{҉!vl�)�=��=0�     ����z��H��}��C�_U��a�i��dB-�޵d0q���S   @�~\\�'l|�P��q3̳�x@"�(�T��L��UC���2��D�>����fl�q@h!6*�2�A0��t:4��b�LBqWp;%]�����e�UD6]��c�'�'�q�Lҵ]��ʮ���O��pD�;;    ����`!O1��\�>�$�v�C����9i��k{�Z]��ءW'���M��u�D)�Nʭ����X�     @e�L�s	>o�\�k�+ա�dU�<;�����d2����>(����   ����w+�y[hh�DLf�������������b��UC<� p7d8���Z܍��N��B���(����`aۣ�-` p/���0����>W���ι��r�G���um�(ص]����S�^�k��T�p�΍[    �����Ǧ�v���~�e�����0��E�:��߯+:1,2:      �>��z��������e�;�u��JN�����mnm�L��c,    ���6�9> PO`�e�:/LNK杧���9�d�����\2���~E�jՄ:q�6��&ĕ��P(S���-C���9kby����
pm'��[tm����v��{��=lgI��4q�*��]sN�y�um����]��C���y   @f�����^�k��/ee�s�4P�k���e\�yF�!;��!�N�N��      ������g��紂v�LSt�j�xeU)7�F8�\�s]w��ԓ����=�1    ���_� PO0������e��������]�Hx�=5j��P>r9aw����/�7��h�Mi(n�E�������0��KKvm����vmO��tm�}�:��=�k�\��j    Dvv����}�3��l�p�jӵ]Ӭ��}Eq���[�k����n5�,�*ωA�$��|��C��       4���F�.!�_�|��w�� U#Sh�|9C{\A T[���&    ��\�@�;?ۡ��Q��5����Y�A��H?��c�*�3F�������o���r����3(Q���R��5��bw�B��8 ����]�CL]�}Eٲ��$ճ����.ӵ]��Z    �^�O�	��Y76W���z�v�����
AH;��Ǚ�s�*9)��*N������Љ�!�*      ցaV�M�ļab���d7��	�,Fа"�3����3C TW��)u��3   �;��!찵��=���F�{�a�#w�q�V�{~4�F�LڝvꪈD����SyTx`j�����%P>���$�.ϵ=��%n���D*q��k�ԗ-����)�^q����!p   ���G�q���y����z�����k��ڮ�:�����N��P_r܃�za|�k�<�-vI���       � 3��[�D��.q�{���I��-wu0q;�(�1@     �F`|k6_�Rް�-e�_ۆ<�V���/��s��|!W�r<�& �{:�*����J,����Q�*��H\(A0��0�.�j�k����ȵ=^���c   �i�ظ�\��x��u���k��
w+���o5h�����Wn����S?*W�������܉aM      4�`���	��屾8�O�V�#|͜dM�ۋ�-���7 p���     4Ƒ��v`:O�d�N�;�d��wf��^�Njr�g�.���B��&���f	7��	q�3)\�(S⪘U�����!�ˮ�ĉ����\�#B�ԎPV�k�ܽ���r]���a�"]��Sl�[�0l�A    �i����"\�M��并��˴�uvm��k4���l��o5��@ռHw�'�+r3Z��Pџh       �`0���X�+�3٢{�A��oo���E��L��g2�1^�?/   �� �^o��nf����C�q�"g��B�Pz.nO�*3<�E1p��=�N����Ѝ!���Rߐ2�_���,k����m�s9^�
J�ȵ=ֶ�����]ۓm9pm���}U�v����3��͛p5   8d'���V74�6i�,�v�x4(�f-HNT��W�$�
2�+R��=4%R     �p5Y��Iqf���u�_�,n�jn0�]cY�5w   @�Ÿ��[;���X�ӭ���A�\_�����34�<b�Ӧ� �{ڭ�i���v⢛;&]���Q��]q�u�w�T���|?(ӵ]�N+��gԉ������=�'h��ӵ=,c�?�t���  �l��x�(µ]�@��4�vCq{IךO�nVw�v�����q᜷N��8F �����zb[r��m��4      ����t���ũ��w$lOI\7E\���yC;\�  �3�ш��~`�   ������@}����{5�j���>��BS��V�9���\ix���I�, �Lp����`X�f�����<��tmg(��M]�5�\�e}��	������U��Y�{�9ђ��a���~B�߻���/�K    �N��Ksm_Aܾ�k{�y���QWI�uu"�������gaA�U:Rcܯ�@��~��'      @���:4�ƻ0��ƄI~V�Z�<R��6�Z��`���C�Uj���}�����k    ��۷����@}]b�g�uA�.�)O�Mf�fX\/	�U9C.���w�)@��ߋ_.�M-�S\�n#�5!4ugpd��r�B��0�h:�R�n]a���9��u�B�k��8U�n�ھ8s�����g;��ג��.����8{<��hk�E   ��������i���sˮ��Z��s;�//n_յ������6��|�,�wU�*��'P��A*V3      �j�j�h:��%T#�D�����)V2��k|�����w+� ՙãCzt�.�   ���wn�/���@}�0����Ύ�����v̷�Kܕs{NG̻���1��a=��Vw��o��r�9*#�&����z���cQ��H�n���-v����,ѵ}�w��]�))_ڵ]rcOз�ڮ>��\ۅ㮋�|�   !7�nқ���B\�U�õݬ#�-�������ŀ@�T5Pe�2U±r���q�U      �-{q�u���0�����'����3dl��
W���r|rB����	    s�wvhpqA���9���@�4i��oڬ[�.�����4"�pݮp�s\��vs��͹�����V�-�M���X䮉L���C�������7Vwm�K�����v]��~Q ^�k���#�jv���L��G,�;�a   ��v�[8Z�v��sm_�����D�1��A��^����!P     @=�Z�x�N�|A7֟��#�	�'U"w]�`�4a�s�ilC�n��xL���I5e6�Q+��    ˏl�:���l��g��k�"ͷ��w?�a�-��-�'c~�9��\i����U���`��������Uڭ�d��`ss����\ t�vQ5N��m_����c�d�vm��z:Az�k�t���I~-�qm�w�   "�H�,��<a0cq{��<�V��4�����&�׉�//.	ء��*mP*�,�D�*u�
�*      ֈp���?�"Uݶ�QZ�����3�r�MI'���ሶw0�-M��      ��C��MY�,�[���LO9V#��UZ�לE����`<kQ�spo.U�j.ZO&��U��ʘ\�UYg����7o��0�2�n�L�vr����EQ�����}M\ۅ��?��n�   4���F�!���k��n�v]��6��_bIk42P�,�>����f�"wYC�	T     �.L�v<~'q�*I'��|nn �S�+A��U<�c,{0!��N3��    h8X�UkF�!;d�������yp<���#H���yY�<���7��=��6��U喃~�+�g�B7fC�}�6�Z���o�����u����}���'n��C�޵]|�tm��WWWt~z�i�'RI��\�Gz$��������Xj�\�������$k��/��d�J�~B}��P������)������jъ�kg�<�q��_^^�;`K��k��9W�O&g}3\�������嵳��3�a��5p���~4����s���ί�#��Za8��6��m'�6���Lo��?8;7vw��_D��˜���Ճ��̺M�<�y�d����ɉ���s�4�<�7n�>�� P�+�T�s������b�8f�;      �c�/v~&1�����7z^h%eq�^�����v��Ԙ�X    �0�LW��h�q�-�0_K���8�ǟ1��v�����%��3���=��G[�`=��O:�II��F\��0��L�/���C�j���_����*�^�\�^&4qտ����1���h�P<(Ҹ�����΄O�oފ7/'�W6�����UH)<9>&6���U��PInvN���oG.;=9���_��ӞuX�P�s'��B�������@�w*,.�����Q`��3�/�����J�����&^����=τήv�py��]���N'�q���[�}��oo����:8:�%�6Ջ_\��{�<|E�vS�{����mj�Z�P(e�zv�{-s�|u��	�ٜ������\��]�-�(�nݺ������t��.o��
�K�7k���     �c�Ue����Ry(1�,˺�ӎ���Juqg;�r���Z</_��j��{W�����7��㓹iE��\pq>�~��9������yS+�p.����>���\���f�k�r��_{����A`�����}�̙�!���Y�.M ]�w,o���������[&���O���_��]��{���kt9��S�c���C�c|vϹ�[�Q�yݹs����*�x��������y�0��MG��ae��Ϩ	@����أ��c���7�ue90�n�Ď����	1����ࠔ����	�\�g���U��O���{�&]�tm�cA�O?��X �s>7rm��3��Vp�Oo^��W�?|R�k��v�Ne�����(�De����O��a;Ͻ[w��l�p��=r�l6�P�M�l�������%��g�����+\�w�lQ�����{.py��g�Cl������l]^;���W�����MP]��g�$���G�Gt:���[7�-���svzJ}�qf]��\'"7;/V���?���Q]�����O��{���R��kN�v�{��)���d��rn�FY�
�h���gM�#:%UIq������0�G�@�/-x      8g<��E_�E��X���(U&�u(�ں�6ff�Pw+K�biL|�0���,D�vߟэ�{V�f���'g���a׽��C�H���֯����g?��~��/��]�.}e�⸮�f0����Y\jww�I߮_{����<�[�����w�q�?��{ޕ9����]3��7���u�i���}��:|W�w��ɩ�1��8#��7��햛�����K�c|��c����Ee�yX��h���D�8@Z��i�C���)�@��8��*e��H�jP)p��P��J%��UpP(��P4���_(�r�i�	ѶFHN�]�ħ	ă�^��=����[ �Nr9a����m露���{�>�ՑNU��|���5������Lq��^����  �n  ��IDAT �mn޼E��pX7��\�j�dX��t�G����<��4&�W;������	�A��`��V�U�/��x=�����_h@�� ���     `]�<�h�������:f;?'g���K�ܽ5�-�y($2�T0������U��3���b�n�k�?�^�G�����;]��>^����G�����v߻�����g�T쳯�������"3csտ�����L����5ؕ����.���{�>Y���>��^�S�wq��v6�`�g�t��X}�c��]�����|���>���<�p��}�a�0-�m:�Ͱ�T��D�0�1��.&5^�.�{�G3�;��q$�WM�6B=u�*!tc�(���^7�2�۷o(�p��u���(�k�P�8a{�@<�k{�?��{��G|���BJ^sY����(�8r�   �D�-n��KD^��� �vMFuWum��u'�??s��aӸ{�n��+��� U2P%
�S�}��Ѥ@      ��ńh;�r�TC�y��� n1��G�r��:��l��3��K�bpA��0��v2    ǃ��v� �s��Ma��2̧�b����
G�P�.�+���1�`ܜ�.�\rp<��A�9^Ȯup���bPkފ6q���=/�!�ځa���dsy��>�L������Z ��W�k��������\ї��]U��r�*   �-����d}�.\%�_M��Sߖ�ڞ�g*n��K��v`�4~���n��'�L��a�j�w�^�xI����@      ��E����M�d�g�^\!s��� �AV�w~f�X�|��r�    ���M�\`\k��H�J��Bm��X~.�#�����1�,�o
��`<����7C�=@|c�7b�����*�;Q�T<{{{�0\��M��.˵}�c��5��'�6qmW
�C!yѮ����Bv�q)�v�8Sa��n�Iާ��A��Ǐ�/�    ��0���l�x�v�)��ȍ�jO�������*ܺu��A"��^��R�┸������`�|�A      T���O���z�O䅯IS,mB\)lg��Bg��"��� ���3#e�   ��t�]��	�6�]	��2�4�"��P��I�C��}~���G��4���z��ጚ�9���4�L�`C�;�}.0��v@ws�V� p����|!p/ɵ������\�E�wm'ѵ���s��g�۽��?E�^�k;W���>��C   �
[�up|�|�a��Y�0��v��e����^�	�S��H�����a0W峎�����(;H�����0��ے��"~�?�      �Z�\^����1}�N讛7H	l�����v���e2��x<�_���;x�pxxH   @y��!�y�O��/.i6k��%��\-��u:�0q��D}Ew�;��	�$�������/��a;D�*������U"v��� �*��A�n������>.ϵ=C ԥ�]��sҜCQ����R��B�
�zX�Ե�/�N����E   @Sy��1�x�J,,A�n*l��5�W׵�Z�{l3h��`}E���9>+� �x\����]�ڼ(��n�`dW4      ��l4��v[X��'�u;?�[��u�V��s��7o�$`�������]W^�yM�<�/���   �&���#��_�;���]���N���<o�;^��*����)9v�K����e;׏O�1@���V�+��P���C�0��Jv���ba��+r��U<����K��������$\ۥ�b]۽ص]#W�{q���N����.p]���i  @s��ؠI��]��=�r��4�v���k�����	ء��4�@�i�J�DQ�8X���ɟE��      �I�z�.��&�I�[���5g��Ur����bp�{�9=;�O=%   ���7�4	�c�c��aY�Ue!��)=g��J���ۻEe��\����S���='�V/Le���8����3X�%+ڋ�W��[����$\�Sw��tAz$���/���mõ]�w��n��v   �(Z������j��F؝K�nV����U��������*����-��MԋHĸ@|�$P��:q�P�S�׬@      �D��[i��x~>gu��ynܸA��՟r�   �3��-�vp9Os�w4���*�h�;QjA6�nw��7��='�3�iHT�spO&��*�����"\<�c�N�����\�v�޲��~���W�߃E�����L]��g/��R��M]�úY"���(p�   ��>dcJJ�W���ʊzza�Q�"��D�Zq��9��+��>���w���|�Yg�>��p/����2~�O\�ɏn�Tq������      ��x����} &�s��崉d7v~����G����)��T#�   �߃�g��5���\���;&�s_Q+�.�R��a�0���R���='�Y�Z�ʈ�{��7n|��a���ʋ� ���N�⾿�O�\޽d��P쮪C���ĵ�Vvm7�Ǯ�gu��M��SM��tm�pՕ$Z_A����"��5�N�3�H   @�w���
e����z"[[�v���	ֳ:��\�u��߿OU�Ѷ�^4V��sٹ����}�֬լ@      �=^�r�X�<o8���pʡ1�r�34���"��t�o՟�hD�.b   �s�>Ů������6`�R]̯th��F"��D���q�K���d���g굩I@����E�aZ�Jn5 mC.܌�Q���~��/�*3�S���9m�A������&�1u�=#�����a��
�v��T�k�ԡҵ�TBrJ�G�'�������+��E�����l8���V��   4��}���j�m��t�
�vsq;��o�������(�~�Ow��u}ne
�{H����~tK��'�O�      �Ʉ�9�IIg"J���ɼ��9.����Y#l7ŵ;{0�{�ӡ1��AP����+�s���5   `�O>�����@��a�������V�l~�v|�pY����DjG��:_�I�1u�c� �99�"�$�@�p�rN!��[�����E�!uP�0w@`���3���m��8�v?�k{��<�_ڵ=!ʷ�ڞ�����ƹ��N��;  �Ʊ��M�W�\c\c�v�~5�:\��]+;�3$^�������0��ڭa��>*�ىRp�
R�Q�JC�Z���,t3#      @�Qgn-l%a</���$�ک-lU����)�e��s��ǳ��|��@�@T����^`�   4��7o��/��@}as����@�<~��z����\�U�st�X\Ԯ�K�ܵ���ߗ3f�5�� �{NNFD��@U�C��=,�׉�V'ǣ'Q)V/�o]T<�����(^UU�k�ؖ"��pm������T�v�8_�Vi��}��ڞ��V+p��F   4�v��kA��\]YQO�7�[	y������h6� ��6�U&�������mpA*��e^O!nWa.��z�       1���1�"�<�3e�ga~`��sx���"��(2��j��y)��3�L���6�6	�f�תЇ   `l�Z{&W�J���f���:oXt�Qg�g�3�����:=q2w�ZH?C�R8�����U�vn�|Ω��rM�*jK+lgTk�Y���m��prtLk��N��<�o���a`9���S���O֑]��kΉ�wm��m8����_��   �&���K�+��]Ʈ���fus֋���ԝ�ھ��}y���芀�Y��^[��G�dT�U\@��(�b��{>���      �����^�+����@7wH5��Y�Y睟a�Um�g�ל����-�q  �����G�1�z3�B��l���T���G}nҜU���9���ỳ�p���v��f-ހ�='��)�6Z�d4C�&:��n\��:煺�Bn߾M��G��U�k���^�k��ܗvm+Ku����\۹��hH>}
�;  ���駟ҫ�oR����\��޵]]���C�Z/�	�l\����6�;��7���0���G��     �t�x�N8�'�b�路�ȹC��Q��2�Z���ݻw	�apvNw�������>~���[   ��G�>�_�ｺ3�B����Eb�P7�����Xa���珇��|ߣn��L>+��~x��oF_���|�g.�ͷ��:�BnݺE���2]��B���@��Ĺ��˩A��B���666   h
��ߣ�����Wwm_M��^D��8�<�}�6!p�GY;lUm��u�J�0F�J.z˓1Y��~�.���       �F0^����$���8����a����'!n/~NT��"v~�����zsxtD���w   ������7���@�����h|�0(ʘǫ4�a�P#�Wc�e��7��}	���jx�8��*.�E��ŉoy����VyE�:��
�f+}����}��k��,Ӻ�+�J���N��|�]ۣs[\e���v�   ��n+˝���[��������.�������m����$W�+�8'�H��	P-:�T쇝��%��      T���)y=/�x'���b�M.T�iq�]���;7�z<v~����ug6�R��%   �)�q(�2�g|��-��7�I�7u��:-q��_H��uixJ��%hw��_^$VG���LZu�'��P:2'r�Q���������|J���4p����#q��k{RE�8.��µ])�V�#��'˔�v�/G��.)�m���\/�ѣG��w�   Pg�R7�L��1�kf��\��ԭ�k;������1�#���-�:�G�91h�T�"���M�C�     @Ua;?��}����j��=�.�͘K�c�~�;?��v��|�;��4L9�TZ%�   �
��	��&0b�g[d-@�s�0�|r����c��9.�����K0i��N�k^��)��!�O��M�
Ri��<iO�k��n{{�<x@/^� P>G�����]��d�U�v��yF�:���ѧ���   j�G}Do��G��ڮy
�/^�^+[�Űv`� ���u
F��p^.�wb�[Q�����\ݻ�M      T���&/.�c�Drz��b� �eeR1��]G�s�,g���������@}9<>�   Pg>|H���	ԛ�xwK�y�a�n���9��4��	ۉ���ߠ���\]�l�H�����Mɉ��χ����C������z��	�8<8��ˇ/\�\����k{X������텺�S���<
���v��N��{'   �χO?����7�ߥ����k�YG���u��tz|L�,�i�W�`T����]��W���NiB�c�q�yN      �^g�z ?H��DD��ryC?�F���w*��]~*m�S���Wm�޽{���Iʅ��g紻w�@}�Ջ��O>��  @�y��3�����@�9=9!`����ޞQݦ�u��E����$f'}!�ݼ�!�K0��i#�"��=d�7e��޼�*���љ��!@������w�R���?]��d[��v�k{���]�)�Ni�틺�\�墍�M8�   �=�~?XإB���L@���q�rD人Uܓ��������nG��9��hn��()~j<@���D���G      �j3]���/VM3Ǌۜȝ���d,�5H�/3%Z��b�ߧ�O��_|A�|N�O p�9���vo�   PwX�pt5"Po���y�X�K����v"}<@#j�bW�B�ǣ�W�ىH�
�����Nت:P%���.�g�&\� �n�a��b;��]�=y/�&����������kT	�UZ��:��A �׿�5   u����ԟ%���j����4��ԣկU>W8�ۃ�U$U۲0�-�������PȞ���~q��s9c��      �ː�ۥ1}�7#9�'M�PN|��yGy������]G�r��w;0��#����#   U��GgT�xT���SvX&o���[Ǽa\7+׭��B�.�-
��5-o������=R'��d5qu�d9���!l7�� �*mC�n��7o]�%7�EY �N���E�*�yY��:Y��j�������+(�n���}��� p  P[~��ҷ�^	ej]�f���`�y>a�j��r������><��ɶx�葲|��Q�m'�!�sX������E����lܼ@      ����M�)�z"��?,�&�bY>�m��e���s����?~L�p�lo�޽{���O   @a$�{��@������W�yC�����=��b��Q��K*?5/o���=��o�R���"ǅ0�-�[��T:�*�Vi�M�����hl��л�K����.	�%q{��z���b��
�e?{�w��   ��r��=��̝���j���P�^D�rD�UܯVW�Z�ˎ��ء����tI~�yT�ށ-�&�3F��Ǫ.a��j      T���G[|Z��V����C!�-΋usa��{��v�1�c,{��!�?_��+����=�  Ԗg�|L�?��@�������~)�V>o���6��#&M�@��~X�ܽ�@����F?3@�'�śS�s�4t�*��*�ȕ�"we���h��ӧ�j�h6k�
WЃ���sm'� ]�72���M��k;���d�2]ۅ��ybM�k{r��ڵ]�<���-��ڢ��   �F�3��uպ��f�u�k�a�e������ת�{�`VW�Z/*��c�����6���Zx��ɽ����X�\]���㓿��u��uq��9�      �ڰ���f�b��o�~� �+TDnqr���y�����J�w��%`���� ?�򴠾�[h~   ԑV��Y�N&t1��P�\�|.K�ބ��J�+�O�J�|{B\���=����o��r��3D�Vn��s���L�L
\��/C�W7o��o޼!P>�����#i{Gc���3�2�1A�^�k{�i/!�^Ƶ}�z��e����^�E������}���   P'����ٙ������8�X�.U<|@�l�ɶ���kB9m�/�$���?<��DN������.��.�      T�w�3j�l��}i~@~���8�ķ2������V��*��p~ZV��0!���ݸ�G��\M'������   �:��΃�%��sr|�9�%�|�ɓ'���a�����J�I�7�ڑ��t:t6j�Bܗ��'��<�bh�U���p�E�*����Si�*�Wm��nӇ~��%޼zE��{�;P�k���òk�\Y��S�k{��]����ڞ�X8��z ���C   ��g?�����X�����nMD��WQpO��f���@�n����Lw�5t	A*�Bt9������ƽ=�$����&��v      �Δ��76h2����� �7$
S��"D7៏r9E�:��[dw�6=	�������o���}����?�9   u������/	ԟ�Cv���-dg����c伡����c��!505���L��^Ȯ
4)n�P�>��!��<J�pZ�\�tW���ӧO����4m�7/_��(ҵݳ�ڮ8�[��]��'���.���܄�	  ����dI�I\��hµ]�Mq���oVq�*���裏���m+����{�q� %��k\?��      փv���3e"��NVS4_P9�e��ù��;(H䮣
�E�������+�s|xDO?~F���{G���o@�  �v0��_��?la&���L�n7z��a�w�$fW�de�۝>5ܗd�w��U���.q]~�Bw"i������Q������vx��5Mg3�[qኮ���`^hյ=������9�F��+�v��{=.//�����   �:�v���_�Za��`=�k�\\�����{}Fm�qm�K p�I�cQi.���=��H�ߩ��ǭ      քv�z�=�'._�����OL�E�T�iO�)PO�ȶY[l�g�� '����	   �l�8#���L`��Jސ���!p98�h;����ȍAvb��A+I�k�� �*�>z􈶷��(x�A۴Z�@|�~�����ǏL�[��[%$O�������뗯�����q᭑�^1��e������~f����Ǥ�ۗ<Y�껗����D&bt�/pš/_|G��W�n������ϩl�A���}���Z�N�Ex<��Ņ��ٵk�W,prr���F�9��嵻���l�.�j�&.�������Eq������eN�p��O��`{���_���kp�x>��<������w�����r�i�S�������ſ�<o��'r}c\W^^����ø0�)$*f�����9�˱=�u�:�</�஢Lׄ4�n�O�����n��M����: -�W��=7ߡ      ��L�^jr�T�)]�Ĺ��%�*2��T-����G�7������ݻ���;   � �^{��5����'�nt!M����@�0��R�0,���z7��`H�9�e�����/����▌D�eǶ��+��~��I����t�s�vEֵ߹���o�(���Έ�M�2&n��?����a�o_�~?y���v�����П�ş�'�<S7�����㿡?�˿�ˮ�{@����Qټy�nݺ]��7�гgϜ�̈́�Lpz��='�����>}J�`BWW����q����=��v��� 8�*���iypy�lA�۷o_�l��ׯ�Ν;��|����g����*E���A]&n�!?6�V��f��/~�o���=�v���� X�q��}�s��3�������5��ؾ*��(���Q�Z[�Ґh.�A<�W��x@�����l�      �>�~�<����'�ùH,lO1ÒY��9��P�W��?�E�1����U<��ڿ����~��89<��̍�����N�N��u#�8=:��_~�of2�����0*��W�������ߖ����9����ܸ̞4ܜ����]��v�9ˮ����I�gggA�M4g
��\�N�y��8_>����Ɖ��y��_.�wt=Ʋ7�G���H�?.���s���]}ޥQ��Rւc�S�S6~qc��ܗ��O����vn5��Ɛtb��ԫ?��w�殐&�b��Ѝ���7o�7�	�"�(�D�J�׉��zi"y�P���|,Y�D}EJv�8Sq��"xR��}�ci5q;�b��9�gp�w�E7o���   �:þC[���`]W/_�UE�y�_}^��ˮk*lW�8�{��=;����,�ܪ�Ӷ4��V��XM�Ȃ�<�����?      jN�Z�g8֏P$�żaXM�FXq�]���jn��Ç�P��ss%<�&�D���k��ݦ�O�c����o���޾|E�7�h˕Q˗_ӳ�����00�x�Dt��?��?��������l�r��3noo�I�M~����igg'0hr�ks&fN�j��/_&*�v{w�ڳ�X6faN�.x����?��?��_��pK���y���{���펽1֋_=ƴ����V�666��})�ua���;_g��V��yãQ3��/����;}����pÆh�]��@��-���>�&LT��W_(�W߽�(\������T�ĵ�O���*)�[�k�'��e���da��=x����o-��������ߧ��o��   �u�g����n�� xl*B_YOe��Wܛ�S��y�~�sUUֿT�g�c{l[�����,�dߑ!yK�v�"�%��]�/�$�g����98      �xޜ�0�'ʄ�v2o��[+���|ar|e����ǇG�	�A������[!   `
ә�_^hǇ�ڂ�?�����������z��W`cs����"w~F�ffdz»�0hR������=�-������Z$�Ƴ]�)ݑ=���]�3��&��K���(����28�r��'��Z�v�̣���H   �����'�������RW0�;�WUpoxR����vm�R��o���G}D���Fu����Ϲ�����#E񀤰E��a����f�      XG�;��g7��{�>o(��!)��3��<OS���U�-2�۷o�{��f&p��g��9��G�E���H   �:�����_��6w����r|tL�O�<1މ��y��Q&yì���=�P������Bo�f��vF� ����58>=*�7h�N�+&� v`� ����{�/7�4��)�hE':�I���TKݚ�3����={�������|؝�}f����}�Lw�{Q��#)�˰��@nP	��HD"��D����f!�EFJ ���c�f]&)�k;�qU�E�x���q�e�.��zX��\�3��������"���� �B���[U�cb��ax�"��	���>�U�~��{��$&������oDG�����`i�}F�\�9 �XEgklnEr�4cqB!�BH�YM	c�f$	��ȍ<�Vdm���e�gA	�n��-���R�|�+���E�hB!q���+��h��1�$�N��Q��P�mM^uC��uк�1Qy�v�XF������ ��,�;�~dn�X�H��AٳgHx�d�Epmr�g�G��X�c;�E�յ��~.J�ڮ�[��3����B)G�;����]�zQD�A����kwC��V<_��k���#���uX2Ѹ��_I+���9q���$Uډ���B!��򢮱���ܽ�kIqU�����X���)�b�{��A|��� �gyis�shmk���-ΧW󛝝!�R�l޼3ss ����4VWVA�a����yM��q[���u��a}�Nա�= s�48�S�*�+p'��Y\I+k����W{��-�;}�8u�L�\۫�O��yl�cP�\�e}����6hӵ���X?>f\"���m�A!��+��ǧ_}�k�!X�k{��Dܮ~�Աc#���d��e�1�T��!�$�u{�j=����RH�������B!��r#UӸv??�]����(n�#��8��P�>VQ�%r/������b�g
�+��~��'�՝; �Bʑ'O��R��p��0��uCE;���qܓܕc}eݰ�
�_�®��(�u��6{�*w���L��xg&J*F|�A�N���X]嬫0��ۭ��u]�AZ.煸������͸|��fl�]�n��һ�;��_۶m�r��B��$uU���݊��][:y�zq�XC��j��=��&c#� �JT��T�W��>�Ȏ��`O\YXYщՍQ[H�tW) �B!��X2괄�m�`/p�
��
�8����z+?�cmq��� �!V��{� ��gqqͭ� �Bʕچ:$	TUW�l|&�s
aP\(�Q7tO'׭fb��z/ݰV�0U���$*
��7���:�c{�vHUr7Y"G���м�ܒW�}b)4��ųg�@J���������T4�v�Ūr���p�XTZ�퐈��v[�W�����XY�[�������3����A!�����*z�}	�K""��)lW�W��u?�y�{�)l�+�SI8�	Ư��
�%FϿ�p#n�ds�H%&������';i^�1�m��5���B!���bj��ƺÚ֊�pL���J�#f�+�_��R\k���+?����8H�03?���LOO�B)'�n݊�	޷Tc���x���e"T/��!�1V��åVˬN,��:���/�P�������WQ���ȴ��擬N~E�P�z1��СC������o�oX�k�LHO�|�؎ߊ�sm�}8c��n�K$�ر�%B!�ƞ�/㇟��u���҉�K%�74�����U��}I��0?7b�������x�у�+��j ��{=^���HD9U)��e`��vB!�Bʍ�y�)]q����,l�'��H�s�)�¸
ԃ�Ӯ]��e��Sx
���ql5�P+���<Ĺ�'p��; �Bʉ�'����wA*�Օ�Nπ�Þ={�c06JMQZ7���t��Z�G�p=��� �U�n
���Ԃ��E��*8�t��Pb)
���0�����p$�1�ߏ��epm�]��pmw��+��um7?c��˞�k{���4Rx饗02BWTB!偘%^U-�7˵ݗ�<��� �T�ך��bGy�*�.i"�JT�,[��p_�j��[|b&� ����|B��w��T�v\$�B!�����$�HL��j��U���bY�V�b��`~�ul��0Ƣ�=�+��O`��m ���e4�4�B)7j�밚H�T½=
�c���M��o��ڻ�u��6W���̵���^E��)pHuCR���v�_��q��zJ�U����[�J8��������W�\��	��q�>Bwm��*׵��66>�3g���w�!�R�8q=�}���CB{P,D�q��ũb��)XW�l�ر�Q���*Q'��ݯ�r43W�Zلu�0E��r�\̤UcS+�����"�B!��YJc�f���ܽ�XN�sl�.r�c'�63X��ݤ�̯���o��$&��(p� �fg�y�fLNN�B)�����H����Hx���+�n��<U�P>�]�9�M--HNUnݐ����޽4�����u�1��:Kc�Ų�>S&N���t�رȒn�HwW��-v���s��[{4�J�ڮ)lõ=ݳC�n�K&ؼcgzyI!�!�B��������E-"�S�T��K���>�~���P2�W�����c�A�����%9n\]�rQ�]w>��K؎�y �7��#�66�B!�R��74aq~6��i�%7xM�d��'���C�r�-�j�J�ё�@*��~ƥ�g��g��B)^;�:>��5H� �IxD1��S�0���&�K��'�L��m��U�(p�\�u��K/aeMRy�ܰ84��.�jx35�Ll�ݻ[�l�r�!�������ع#�k{���q$�k/q��k�뜊����n�K�^����{�����Y����x��!��8#܃�bk�s��5��ب�ŏ5�o��`]q���+�LT����x�ȑ؈�u�wN����Ð��q'����
a��9�M�{���B!���$U״v_?��Ȫ]34��ng�Љ5�`X7�Y�p��&PzN����0Q+���467�|�BHY jյ5H&� ���?��i���JQ7����w��p���� �a���:Wzݐ���Wc�Y��tn�ۭ�n�� .#�/��lm������]��s���I���� ���v�ڙMf����Cr��ҵ�޴����vm��Q��k�����65=�#G�P�N!$��=����wD."W��Ϋt�� �T�����bĮ5��p�������8��r���m�hD9ݰ��'�K��<��7��*^�B!��#KhP��k���-��]�XV�AI	ͱ�Xw4W~nll���H�YZ\������A*�']�i!�ӧOA!�ę׏��_�>��&&��X$��� (i��E�ZU7��)�c�������k2��M�^`)���� ���;a�tb��JD)�W�$��=J�{��tu���鿳�vG]�m��q.q{	\��q��:E���������4!��8"~����HZD."����9��+���Ǫ�U[��8�Xk���0Hx���k�	�&��֞��4�ݞ��cv�DU6��pu]�(p'�B!�,�X�A�b�&]�,U�Њm�(Zk�V����k_KK:��������Do��y��Bbώ]���Jbt�u�0����겏�#Fף����p�=��=�w�a��T���Q��ܺ!��[I�ik#�	������"����3P�h7���<��]�U�\n0\:�>KO�p9�4]ۥbw��Z*l(��\�Q�+�k����s�+�k�3nxl.^��B!$�����\�cu�)L�|�v�� �T��A�P`�?���A����Rn�n��L��}�����yU�������&+7IE!�BH��b6�v�b��G��8�ǲ���!�e�B�z��b~�ū��J�{������� ����Rz2���<!��8"���fi�Xi���IxR7�"�5E[�б���FX.���~�k��B�t��E�����I�D�ډAqa˶�8�C���d����^y����NLL`۶m���]��b���n��\��P]��m��K$ص{Od�[!��|�;����y���pa����b��Vչ��F��w�1%��T�#� ᡚX\N�
��	���cҊʅ!7�ϵio��������S3�B!�R�N�prs��@��zM�������1��@��^XN�W^�X7
�*����gN��/��:!��xr��Y|��]��b|t$<��Y2�6��ۯﺡu��mR�ӭY2C,��]�7^o��o��te�)p/ɚ��jJZ��ve�� ��92gf���� �09K<\^t��������{��[���cG���cB!q���ˉU��܏�=��\%�5�)�rL��=�`
4������b�E������'����7�VM�n�q}�	�I�M\�B!��r&�v_��ڊ����_�,׸���6/�^��V�����	�ŵ�{~n-k�:�����m�BH���55XY]�������*c,ʡ����U��UՍ��j	�%�㦶v����(p/3�z�).8�ŘW����賛K�j�������}���8v����;�p��������æl*�k�zlY��{���mF�8�b�o����|<5=��^{�wB!�����x������\O�n(��/�XC?V%"�=���O�f�y^#C� �!&>�r��$�˶�b��5�Sg�w�,5��k!�B!����o�1?o���4��Z��qG��ݺ�ڇ��Xn�W����W_EMM���^�=LF�F�r���J�yowZ����B!$N[�|�����B�"��8.&V��V7�����{��S����z��KoW:��х*�r\h�|�s��q�ex3���D��
�NzQ�.O��Y�f/ĵ] �gv��<붧�]�]}����˄�A\������
���.�3��󿅁����@!$n467cee%�8L���]u^��������X�K-Lp?��b�c}}}�q98+�"�ב���8�O:����I*�C&a��|R��dB!�R�,��6�Uo�`�p��:k�Yr��b�u8c�(�[�lI��?NaSXAсï�T�{��浛�B�{^~|�	He!&\���X��}6�
�.e�u�mF�qzn��{�d��Y����V�
����)�l�̢(`�A��]'aeub��G��E!�+1+�����"FF��c�N=�v��Ј(����ID�"xw�����*�u���ΰP\۽D��F�}å˗�ч�B�G����P�q�"r�
[�S8�����P� M�z@��y���bl���_!p/&qOtY�Rִ�r�r/�K�]KY��B!��7�+5hi���A�Vl�Κ��swPW�"\�)p���A��c%�@SSS�nL!��a�8�0RY�����Hx#ⰈCMѡgϴ��9 ��N�2c,�6�$�����.�а��^��qq�n�<�r�t�0�C
��'W�|��-� ����Jܵ]��jC"�N����8���cU�v�!�k��+�gc)]ۭm��v����k7����?��BH�>zw�>��R��"��\�b�4�)�+}�
��/5��^$�x/.G�>k2�㞠G�sr&�I�J5�<7n�'P�&�L��E��3Mq;!�B!�Nߌ�W٪My�	ʱ�z2�5ga��k5ȉr�f�P.�򗿀����"f�g���R9|��G�>s_ݹB!$�=w�>��������MJO��q�)�8��_��~��Ms�B�T��ɣ��"��܊��i�������� �*���%�u�t��y�ɑ#G�i�&LMM����'Op����c?��6��C�]��*{c&�p�vg�/�v��8#Pl�:��6C����ə�A�Yܻ{�BH��ر�33J��4۟0\����4����y�Ā��u�8_��4�7 ��88$���0W"t��6��^cxuK����؈�N� �B!���N��M59a��K�f��*�U��F?y��q2�
��Ƶ��Q���_X@k{��!�Ă���6�ayy���{{��q�X1+���a��4ho+�k��f^`�����4Ƣ��X$j��2����)(�e�W�ʌg�K�I���Z�8q��9H8�<�J;z�/�R���+sm�v{<�P=W��r4�]�ak˵�u����#�6��:|��B"���s���GW{iD��*v��^� �c���u��c}��}	�s����Ƕm۰�~đb%�̱��M�y$�;2X������B!�BH��\��onk��kb���"�е��1ctd��k�AꇢfXWWG'���W��T?���O����B���gN��H�120---���͑��P����U��f(5�b�0�Eb>U���pc(l�_��Ȋ�s1*!kT"t?�
������H"�@_��]ǵ=���܏`]*:7�򸶫����~����킢����nH�W���'O�>!����XY���K�NDn脭7_�^
�ZDP����M�󘙚	�ӧO��OL��P|,��R��>�&��ݜ"�d]3!�B!����{Ø�Nn-�f�[^3��#菵�ʤ�h�'rG�U�~	�ѡ���V�y��adl�^}�wB!��y�V|����Bh��G�@���ɓ����>�Sݰ�5E��=7��z���]O�r� Ǻa
܋��Bv���B������a&�T1��C�b�N��K!ɫC�������Y�{9���D��vm�ƹ��7�T���ؠ��p�NNO���S�B��KW.�g����������avX�u?�y��*��yP_"x�dM�� �Zf��LV��s}�=L뻵R:I*�x>Y�vd.�M!�B�F`��q�^?��઻���laݲ�c�O��O\�pq��=<Lq��/�T��}8x� ���@!�D��c<���P%bN�$�!��@duC�x;����˚+X��bR�u
܋ĳ�$v6���0���$�&IV�b2��>�quW�O|��%iV)<}�o����]�a�Q�#X����8���*�A{T��n�W�����Z �{Umv�܉��!B!a"��������j��X=�u���"�b��W���C������=T���Xf�R�%����O��'�e�J{E�u��HT��|&�!�B�L�Ԡ-eX�d���@5��.n�aH�*��A��C�-	���!
�+�g]�x��-
�	!�D�������>�<��Y
�ÇK�����[�P�����uj�NSm��.���X7���H̯h�ֆ��{� ݋TZ,���N���!d-w�'Bl+f�?�$�����,��۳me���n�q.Ѻy���smwoxt/_��?A!����K���I�D�Je��)�=X��k����Ep�X_"x���k�߇��R[[��^{-6���gMPIw�k��=�3Q�˅��3H;���B!�����I'�r+?�c��-JͲ�cG�K'7��B�	'ϸ�47*��8~�H�11=�m۶all�BH��ڵÃ ���"�W�P7�����a�I61ݭ�Ͷ���m+�Y��'(nP�^Dj�Z��<f��dK
�Kz�`��q;A�~VK��+�ŝ�p�|։�����.�������j"l�vm�r}��pmw�� �D������bnn�BH�ߠ����������@�v���� ��<�`]3Nլ+lwƎ�`yi	$<��ݖ-[���\*�>�X��ĐW@R�ř3him��4U�B!�lg���RCV�n-T�����c˄���y&�
�!M~�С��vtt$&�'����ƦF��⧟�֥���Ï@!��ɉS�����T�󘙚	��{���_�FB���[k� $cv��]U3T����1ɺa
܋�bU�t6���ݙ����Y����P
]��P�}���3Hx<��g�;.�wV�g�vC!x)�k;����Nq{�]��{7<6�kׯ��w�!��N�Bw��5��\���4E-X�ӿ�|=���ՍU�u����~�p9y�$*���1v�gfC5d�:r5�m �B!�l,[ڱ8;��甬 n/������fX���=&z�XUU�W?���8q}D�mX��~� �RY�ﶕd---���!�����P�4�>/X7Q���Ƣ6�*�>7��a���;#�5򜑵s\�e��J����Y74����/Vc�5Ie��N)��.�[���YŴ�>�ŕ���_G[��u]]����}�D[}�}�}���OP]S�~\��������O?����&V����;3�����ӣy<�gD"(W���U�{�������̿r|��Z�~��)�����<Z�[��ۛ�.�p}[T�������#�{uu+++XXX���ړɤ���1�����_Zw����f���Td�]�u/�w�{#�(���W��.�HDҿ�[\�Q}�}݉����aK�Z���]������Y�}��>�G�����ޡ;�:���8�������Z(�?��%�����<�W5�w��7�"Y>���%Q�����:v옴����V�}�q�z�{R�鞨?�ݖ�&�ֶ4��PB!�BH�HԴ��&�c �)��v���	��M�����n3���Cq�c�X����>�_jjj"�_���k��� }����=�
z�xݢ�����(X]Y���rd5�d"�k_^{������ĩ������~��[-E�r���Gտ��ﰨ���������BT��(�;�]������wͺ�$l����5�{��>�gΝ�W�~�D26�}�om���D��X+���k��}+��t�[���7�O��ߋB�a<,����k��}�nN��g<��v�4�r�E�ruH��}�ʘΉ������Y�nVq��b7����*k��mSUU�$���]�+�T~�r6�����ňn$���w�ٍ�G��$��P�����_����q��vm7����϶�rmw���$���I}�ɧ�q�Vd��}�	n���3%�g���~�ڽr��o���!l޼�!�<p�@$}����,v��I�bB¾}�Q��B`.~CĵQ����� 777k	SKA��]$����#[�kpp0�sT�����mC[+6@��\�Ų�{��)�Ւ��}� ���N�W���"�z�O��#���k�`jb2�����v�yyT�^������Ͽ�.Q;E��ԩ��y�pp/��Ai	z��P:��Dn�U����R��|�{J21~lI�gVA!�B�8L�֡�HI��~W�2�2I��	��5i/��Za�r����bbLU>M�M#�(��E^H/r���\ZX����`a~>�y�J�%���'VX���os[�&�~bGQÉ
!8�����{V,�~��_�3Ң����Q�k7E�Q�����wET�u�yT�]�-��Q���|�b^��~���c##Z�������B��'#��[Z��q�!�wĵ_,R�f�g��[���7��Q]w^��[�P�ɟ���&����.���6�,�;�n(����L.�м�	Ʉ{v���E�R^��͒���L��M�t���=}�tAn�p�>~��+D׆D8-�{�U�3q��*��<��nt!�W��V�~w$q�;���+����m�v�s��)l��󾯬���={�B����B*��������0�X=�u���"�����s��С@7��?]a�:6�6�$\�d�W^)|I����y��ڱ�S&�MHώٝ��+���f���d4MB!�BH����]�ِ��c���:�q���Xq���w��ق�4B��1��[1@~(�k����K�v�\����=�qʹm�@sDF-bUĨ^��Zߵu���O�V���ĝ/��z�<��Y�5S���znڴ)��+���w���i��(��s&��!�0�پ}{d"o�;�k&4bb�x�Q�k7�/�u�7������$����}��h�o��cwa�ܔ{����E|߶����Ezr�n�Q�ۛ��,F�ޯ���"��
Y�pV/�>�k��f��ayk�5��֟�5�	QA�{��oj��̤ˑ���>�%������rbv�s6�-�*iu��)
�C�������븶kŭ�۵]W܎*�Ъ
���^q�P\W؞nUL p�i�3{���;�F&�p��M|��� �BJ�,��y��v�����S���k���\�׵�J_��p9��kr��r�gx\��M��Rmv1Jʐ��S)�s��[�'��"�B!d��;��k�k������]�.���1F2��������ҫ?��� �1��_����7B����Bc,B!%���		#K�0	����p9w�\�Ϥ��<k�^�r�l9֚!�f������������c�P�^d����.�q��
��w�Ju�g?$�f�ʗ���*��
s��������Ȉm�����.(o�v�ݩ'�'Z׉�OѦ-n��2�v�+E�.�7	�=;v2YE!�d�;x ��p���GX�+l�4_�4��q���v?�������9���'I����WɈ��zq�J�a[�{�aMd�T��Ĺ����B!���Gr�~����s9C,Պ�V�6e��^X7q	��Ͱc�{q���N�{���σT&_}�-�_��/���BH)�|�
��p�r��=l��pe`�f���(Y�ݡ��S�S^� ��X�H
܋��J-�,�jg�ZZ�NɒUގq&2�9��t>=A���A��>}:=[O,�C��ɣ�i�����ϵ=�l�s�R��pm�ŕ�k�3ntr��x��!��br��I���ݻ�����}��Op���U�k`���1}	�5�T}A�~���L$<��މ'B�/�}����=�?^�u`0ۗ��Y�B!��-H�����]1nH�
้��L�l�w3���se�6q��s�pp�1V����afz�� ��pӭk�Gcc#���@!����,'Wi�X�L��c����#�U2�P�+�>Ǆr��Z��~��c�o���d��DMH
܋���NVIfWH�U�6庸��*+�6I�*��7��y(N�J��Ϝ9�/��$<���#nܾ�%:7��m"s3n������ڵ��~��u���θ��U��s���9��BH��Q{����g\���w�avp���ؠ"�u�8U�Z�����{��A�e���8v��\
�O༗7]�w�:I*��==q�>�����ZOT���@�B!����L��)y�0�����2�aH�t�C�^�z�}�fXSS�D�c�0|ч���A*�o�����.�O?!�RL.]��/�}R���L.b�0���*�ڠΊ��ڡ�nh(�#����87����.�N�ցu�����.lopϮ��#Y%��B]ˇ�p:0YA�I�M�B,�A�{���crr[�l�4d�rq���B]ۑ��µ]7�0T�b�����[��_�B!��>s�=]�u��X��ZҤ/�Kخ�U��
�u��Kp�>p��/�K�bYk*/^Dmm.E��RP��v�N�q����*^�&�$B1Q�B!��1y1W�����c���X�%z��q��l8��ȭ[��'q?|�$<�zzq������jkh�E!�����bae	+�� �K��p�����$�_�P�;|�y�v���=>�������v,�NggZ����\�:2�Uָx
�K�� 	��??��פ�s�k{�ܹf���l,�k���һ���S�i���z�`]ߵ���.�Ov�܅��6��΂B	���ڵg7����"B&���g����µ]}�c}	�5c5�Bܾ��De�qHJO4!sa�?&�wU�� �y����Q�N!�B�F�s"��Ȏ�u�|�g�c�<c�9��YV\j}A�99{�,�!39>���9�X�0�������|�">��B!��ҕ����; ����4f����ӧO�8q2�r���G��5C�����sʜ��m������Jd��I������ֵn2���ǒ�̝�D��!����KKK ����?���ktm��C66��w��K��nA�ܮ���������_�
B!$�ϟǳu�v;*�^A�P>_�W�X��\S��)"Wӗ�^3N՗</�z@�E�?~����>kj
J�v_����w��{s�`�B!���j�@s{V�uC���ڡ�.���Y����ns�8	�i��1������_�L�W���ʸ���́B	B{{;f��Ƌ�r���y�U�=}UU�����j���f(�*r�MH���朼�Y;\ۚ�:����@T
�����:tH
�Ra{�����]X�aKT�	��pI��9���'p��]��x�ۋ�il�ؔ~l
�]��R����������W�c7�k{����õ�~@2�D��m������4!��B����܁�.�v�[!��\�+U��Y�v�SRח`]3֧�^���_􁄋H���	���t�槠vbp?G1.�LTW
U��z�ru�}�	!�B!eGCR�sҺ�z�g��!nי��^ ȞBf��ĝ 5L��.�M��A£����
��{���K���A!�A��t�s�ʦ��H���ק�Sq�񕂜P�ږgܭ��j���1V����%��x�kSҋP~�z�܀��aG���Ǥ��,���r��=|���8}c�ϵ�&{+��u�ܮ����.:w����,�k;4��;��z��@!���k���E!�V��]M��K[5�J�\����c�����..\@]]]�q9'���!+j7���*���Dx"�ԮJT-���*!�B!��d��˙-��������1VX�Z�c�ر�'O@�cblK��hlj�LV	�$Wӆ
333 �B
a�֭����d�
gnv�SS �"�Ž�IX��(�κavlI��f��S�񾗸]l�+�k=r�
+����Zv� ��p]��V}q;g|T�wy���q�e���jߙ3gBs�'9��.]�\|�v��Mi%���%lW�mD�vY�vmw�'D=5u�8p� ���A!������M��<�:�h
ƃ�K#���+Ϡ y��Ԃ{�� ����>�Ν��3a��{�1�u,m}N^��c/[�-;���֘�!�B!���*u��X��.zOIk�^�XY�B��1�}w\j}A�9�)p�ߦ���z�r���{x��u|�� �B
���Kx�A*���^��9��vl���B�9��.� U�;_��Hyc)Vx{:Iͫ
�KDMSV�G�3.d"w�s{Jq�{$��[VPk(��a�$xQ�����mmm���,Hxt>}��5�ڶ�L�!�ѐ�����;�%n�ĕڵ��f������v��\�u����;cG'�p�����p�	!�_�z�6����"r��Z�d���ǪE䚂��"x_�{?�����h����Muuuz�W�u�Iw�ò�]��6s�nNBw����Đ�����nY?M��}�B!���N��*�o��Z�9;�P��������X�:FPs�BS�~��i����	�ߡ����i}�C�`?z�ihA!�G�����ԝ���n6bl%�U������k��K��9��ݜ�w�1��f(�mni�� �N(p/�h#7���\��}9��L�?G��)�r�~���>-����A�嗇?���˱wm]�q��������g��ݻ �Btعk��f����ڧ��������XC#������=b}	�5c�7SZOW����A,--��ˮ�ϠH{Q~I)�~2������`D�[*�R�k�T7v�B!���1�*4�n��씭^�9vȎ5�.�	�y�f��H�ެ����F���]�t	����7���������R�<�|�߾�z{z)P$���0�9x����G ����&�'@�E��~��ٲ���ϡǵ��}O6W������ؼ��%��\5�(�!�.;`���R��UI)�D���6��e�&�T��Ν��=�~�-.]��h���+��ݍ�8�g�v�k�@��θ��9=v��	+++ �B�q��E|q�kW���Ї0�8�u�8�X��{��vu���իWm��qHX����r�݉�֖w�+���8r3)Q�!�B!��rM��X`B��Tܞ�j����9\�ӕI�PF�k�^X���с�'O��o�	��������@*�����3g���߃B��¥���ӏ �EW7H����M�Y����vh�*�堮%Z5�*lU�P�/Cmg\�����D<M`oG���t^�v'����r�qHh�x1���O_����a�m��qrm�	��Bt��%�vq���|�����]�!�+��oxl�n����B!ċ��N��}�Z彟�`����u�0E�rm� ��^36��[c���zzA§���X�ڧ�^��&��x�D�غg�q� �B!�D��r6)��ұ�ȇ�P�\�Y>f�b�w2[��Xs��,��p���w���7:���^K��Nc,B!�hjjBcs3&&��M��'�{@�G��k�^X���v�p�to�ku��T�5k�K�ء��D����v,/�ۖ�9�e/h�,_��DUF�.v�~�A���^{�5�޽ �������mM7���{����3t�
tm��IK������ۛ�smwƮ��b�Νزe&&8� �"���/�ۋ����m���f�J�.��F��US��WDD�P���ɮ�Z�_�!��{؈�����c���8���xں��8���.�[��ּ@MM5:�WQ�	�B!��x�h,������%�mL�{�|�Y\�X���`���\#T�;}�4H����anv�mm �͝{����+��OA!�xq��5|~�k259���i��Qǳ���L��V�j���������N-�@��
�K��Ў�ܬbօ�蝛ɑ���)��־d�*�{��R�S]]�^.��#H�|��7����6�h�p���@۷k�K`noL��Qe_� ��|m�4N!�7�?����~b�q�øy�6����B!D���7���/鿕�����RN�
[I����
=�] �s��q�ر�3&�	+���'���8���U�b���}3��B!�R)L-&Ѽ��+�9�+����v����w�=��y�2�	.l/A�hlڴ	SSS �"\�_;u��Y\\�J2Ac,B!�l߾�s�\��}�>�v�±c�bQ�Y��RS,���*c,������S�ˠ�����ԣ�Zȶ�eEoC� ��eq%�r�&��qHh��@�{����ap`�v��
�%�k�F�[�^t��u7vC3�}<�bvmw�K' �vmw��NJ���j�iU:���NB!V���Q[_���y�}�R��`=�of��ͥrm�=Cf �����~��˴[٨	+�3'%sb�?�˽]�(�Kr��- �B!�T5M�XYQ.I.K����O�0�a��uuu�x�"�{�=�p�������������[x�wA!��8����C"���	�+W��W6���U�}&�ڡ�fX��۩�U��,�4p�+����)�uñ��b�A�����5�U�{��z�~�K����˨��E"� 	��~�	;w�;E�R�q��=�k{�/k\Vd�+X�'lw����\���a;�1��A��;&&'q��%tuue�S!�B�o\���?h���ڮ��{��]������j������B�.v�}^�+d_X���=�[-�U�Jm�I�#�k=��B!�R9���v��b]c
����cK�gѻ�R�>��3���Ħ-�A*��=�Gc,B!R�;�_:�M�Fʛ����̓�ϙ3g��q��AZ;t�3M^cn�~���i��z��;��D�Z�Թʠ����M'p��iA[v[gpd.�TZ�.�px�JTY�K��`1����;w��ѣ���A�廻w�߾��˵��h��rm�;.�k��|1��a�yč��.k�����7��'��B9z��H&��J��߬�߂�f����q��k;�b���ݝ�A§���ϟ/k�=8��ck��)�ߪD�s»�:�I�B!�T���ؗJ���e+>\�Y 3�rcdk&q�r�����_D��=��4O;���7ޤ1!�b��}����>!q�H�G8�_�t�,�����ܣ�@5Ô�_�8����p��9����ж�S�v�l����B�������ڵk�G���4�?��GC��.C%n�=���[�@�n	v�����
�!�X��%�)�o��Kس{�mۆ��!B�l���q��Q|�ݷ���������O�k���Bjo������0H�\�z�����~I喰�`q1���%�rb��t�dv�+csk+F�� �B!�TO�8���=!VR���+?��1N\m���n.�o��E��A�F�ݻ��� ����'Ξ.�$zR�|u�[\�v_|�9!������o@�@����y����*v�����❃E]�z���\+?Kk����\��P�U�9f�A�{��C�R�YQ{\��~w���]�*����%Ո>���G�	���j
�ڮ�]�.��G̸����ѵ�y���!��7��ÇA!�����m����\�R�]�߬�ڮ/�WtԵ�G�����g � �K2���P�c9�R��3�N��D��q�,Q�MR������M �B!�T��ܱ�3�Rw���l�m����i�%0�@:ò�8����7o�w��H�,.,bx`;��!3��X1رs'���A!��ٽg&g���� B�}XY^	�7n�ǽ����Cg���果�Q3����Ա�(��*(p/1�S�x%�t�u��-c������nXE��$��+��rHZ�9s&�=::
.�����G����R�q�v���a��[cumw?W!�7J��.i*����ﶉ�)<x��� �R��y�e�,�aii)Ӡ)��-B��TDnh�>�+4���⸶ku�!6���>b�A��U�L��G��\P�-HU�})k�,a�tfL%1���tp'�B!�Y�i[Lz���&�X�9����Z3��I�_C���/\��������!š��9�$����۷��7_B!���g;y����bҽv�H�G|/^�����<����O��v�f�|�ܭz_��˹��|U�Z�)9���g�xu[�2Q����3:���[��������|���U�sP(V?����~�:���?��K2����p���k��ն\۝q��yqum�[��mn~[�oC"����
!�T���8s�Lf�A���L\�3�
q{�#��5�_k9����a~n$|�?�ݻw{Ɣ��]�a��[�{���g�9(����<@2���q�0B!�R�����%�[�9�P��5C���j���1�#[�0�[��".��+W����333 �������hhh !�s�݃�k'=BH%s��U|��=b�Y�g$|�oߎS�Nž��2�Eǘ�! ��VTKY��)�ڡ� �g�������F�:�8=�JT�_�ܾl�5a�w�A��;2�X3��ﳾ�D��O�SђpD�����KW���umO���t����� �v�u&��Xw�8���>sS�Ӹ~�>��CB�,nܼ���vu�V1\�u�TD�K����
���E��N�h��V6��=_�E�a<T����2��}.Y��҂��!�B!�Ƀ�$~�^%��*~K���J�n��r�X&z����uㅸZ���}�]�p�q_w;
B�cc���CGG���A!��زe�U&��@�I�����E�͛7�F�&~kva����׏EU�f#��z�1�}R�uºs|�to����ӱUHœ$�!�Pպvq��MRً�)�Ca��+cm�&���FLZ	�HX---��K_?���c���cma{���[��pmw�\۝�b��rr�O�Ə?�B!��֭[�Z�ᚙu;u�Ƶ�_���Jqm�s^��p���++����1X����p���f؝�������e]K:Vqkh�B!�BH岚4�ھ��Z�v��ʶ�y�C�9��V(#��C?�/^��="��>����x1Џ����x�o�BHeq��U����A����.�h(�n�7>NuFk��Y3���녩u�j���c��6�oEr��v/(p���Z���Đ�[���%�Rz$[�ʐ�z���(��զM�p��y|�� ����������Eumϴ���~�9�D�n����#��ڮ�ƾ\�3�rq����,N�8�G����$����cW�_×�~mk7J��U&��~b�	�5�T}iƩb��p
��=G2�	�;v��2�A����ջ�d�-9eMbI�S�Ñam�2��z��;!�B!��r]���`���f8����s?"�,ֱ��6��ʵ~(��jjj������	LON�c3'~������c�8y��!����ܹs���O�����gld��3 ���؈K�.EZ,E�Q����=w荵���c{���U-��#��=������2J�7ð'�d����55;U�����F��^�~���)p��o�|����ۨ��˶�@\n��\���vC�\����hS��u��>���;��zWKP�OA�^$�?4��׮�?��?�B��F�={b�E(�k{i�tm�3�Z��=��A��\�,N?�e�$��{tD�V�H6����u`�nI<�`��B!��Jgp�[�IW�Pe���:W~N��-�-�1��0݉�
΅k׮]8y�$~�����~��/�!&��8z�&�;���� B!���4��a��b��Y'H4�U�6oޜ}\��A=�5�t�Ϛ�l�m�S��貚�������sB�Kc,/(p��Q��-X��T^�r�7�C��ڮ��.ITم��s�HI��W��~=�8�D�p�3��T��Va��;�urW��%m
a���zn�q���nm���Rk/��S���O ��1ٶ};[�1�ە~L�v"r_�u�8U_�q�X?��f���xz#�Pi�
�q�fқ�c�9+���Z���M��K !�B!�΃�q��*i�P9�VQ4wn�X�B�cE��^�c	w
ܣ��yN�;�jO7Ri|��W�}��{�]B��ܸ}��1�������^�h�|��vlj��9�e�l'{���:&�kcFzu�ǣ����X�nY�8��I*���ʍ!�pf���	,G��I&�.��ڀI�W^yǎCWW�������%������Ghjj��MMN���3WlZ�G�n����&q�����]]Y���:mq;4�MNL�ɣG�P�y�N���_����S5��u��&#C����M͙�aۖ�X\\͑aii	��ш�V֮7�:�n�a"�+�򽟟����F��ƣz�(����9�����!
�|�b����Ey�WWWG��#����I:|���ct>���E���	�ڃ��/�/`d`H+�Ϗ���}a�����K�a�����|<��q��E����C�*��U__�.����7�����Q�13����)t���M�Ei�ʑ��6mںvSB!�BH����Bk�&,�Ϲ��b��]�9e]�\��ܬ�X�T$�1S�!W���6���?��?�����e�����W����U<�|�S�O�i�E!�s����_�uTB��vu!�J�o��ѕ+Wʪ6����Cg�����83^wX��ElK�f�N����虯�n�l����� b��'�����������^Du�7n��Ӿ��� ���³������[�nͶ��ա���'��m����U�׺\����l��D|
۝m��%�F!*��ԑ7.=�U�q:�?ѿx�U�����֖Ʀ&4�����5�g%��_��&>x��P�QN*�OM����;*�{�ｘ\ ��('4E)x��q�E=�,���D�������x���������GCs�4F{▲����g^�[�N�R>[[D��x}�ucSc�X?��oU�����ٿ�`��u��j�
�T������U�^4�{�8���y^b�������R'��Z�0so�qiQ��wmw�mIT+�I�YC|7��:!�B!��O��}m�0#]�YV7�������k�"5�Xg[k
�8��\h���ɓ8p�@��D�ӢB�R�9G���w=y��E�&�{MOLF�W������,j뢑MLON��i'�@����I������ً���qP(�OO���Q &{���"�?��u�hff&2��(_�����f���龣�WG�ދ��0UQ�ϼ����o�78j��KKi��dD�
G�;u��l�~r�+��mog7ZZZ������{N��G�}��}ٿ�8؋r�z�ˌ�UR7�cV����I�)k��CО[�-�x��$?���/ëػ�Z����ڐ�1�OPْU�$U&�S��:]���V¥����m�ė����s�AT����;�=ë�_�����'himŎ�;��Tn�ra;l���vK��z�f�]���wm�~����Giq���һ�[�����?{z���!l߱��}ss3�������_�ԈH��+LĄ�(����Ć�6DE��H��6��>��Q��"	->�����k��bBUT��$��;��؎;��ц��zt4�ɺ�m����Ԧ�o�7m���� �����Ɔ��;Ա��k5|(��؆�����v�4O@�ZU���d
ɵ�����yU��_�de�(���п
�y]�~]��qpf~��o�xٺ��_g'�����	�2���9U
�	!�B!���:t��d�>����+J��C[�P���a�%����V��K�-ꆿ���\qQ	�L�IT�CAX�]�s��lڲ9���م}�"
��ж�#m�Btv�ȡH�^^\���8v��'����]|6������o��_������NOv�Sؾ)���(_{��������UD��E�xtt�w���~�ܹ3mQ���OL.ؾ}{$�G��������_�/���q�5�߼��	TUW�csD߷��G����pZ����}�5>:�񱱒�CT��B��ؘ�����"�EV6FmP���U/��f�w��f��f�����༐ns��|P���ܾ��S��v�f�ܽ�� O����_G�&�N�>��_~/^� 	���|�����.'[�v�8/a{�5�Nw�_a���=q�?|����	������/`�� zϞ=�A-!��򦩩	5uux��ܵ����ԋU��5���}	�5�T}iƩb�ܛ{�>�$D��֭[%wS�S��:�0Q�:�e.=�tWt����B���d��9vB!�B���X7!�����e��k��TW{�����Zfxe����ʋ���~��߇"�%n��>���A��y�s�\�r_ݹB!�}���o��}����S��qㆴ�k�������s��V�,E��1����h$?���bM��:�d�-I%)��
����$��%���P�Ф����7����˿���X���O?���\�*s������jm����S�i��%q�#g�İl�R���
����ڮ�?4��7o���?�g�B)_~�֛����E۶�Bq�ր���rm�o�!��:��ˏ�}?�5�V024�^�D��˗�u����%���������/nwO@WNZ_���&��6m�1Jq;!�B!$��������0/]J9�Eu���=~mrg��~�������uD��s��u��El۶-�dK§�yN�=���hV�$�ejz�+Kطoz{{A!��9x� ��3�fg@����e����}T�ݻ'O����|�j��14T�y�8����LB��z�]۷�M[�<ŉ?:P�"�ӵ؟JJT��;���0h��q:��?�z��R;5���n�G��|���~���Ɋ��^<a{fO�v�c��vm׋�o�~��_A!�<�p���v#�v�j��-�����#��=�N,]�����ڱ�̠;�LP鎩�"vU��S�nYfp"%�=�dNB!�BH����fg��C��f���E�.�D|��nh��+�������o������I�&��;B����!޾�&������B!�X���#���矢eKq���y�,�DÛo������i��ceƀcP��W��2>�2�2Rr��bm���������k�ASخv���l��s�����V.\��]�088>�}�x����ۛm�k���@��|�����*�X]]EuK+^�u���� �R^lݶ�mx��'�8L�zԮ�b}	�5c�
��k߷��--.��.�QWW��7o%U�u���+D��ڲD���������B!����xI6�+B��6���E�O����X^��KL��=::?���(����՟?��CB)On޾���|BTt=}*c�����;g�e#[�����5��
k��W��{Zȶ ���=D�
�[�05�Y�v?^OT9f|�$�,�KTb�������I�1���+H4|��g����o�um��!�ǵ=ۮ-l��	��.?����m���x{���$N�>��1;;B!偸Ǻv�>��N�!��[>b�ڮ��^�O�(Z�,��$\Μ9����E�$��ߩe������ͱy.Qe��&�Z��0�GB!�B���ë���5Jw�����nuz/h��y�s\j~����իغu+���A�gzj
c##���K ����2���������CB)/Ξ=���aeu����uAQ!j��s�Qj�:}[k�~D����c򹟚������d�uC](p��T�SC6�|38La{ʲ���̑A�~�q�.,�T.I�k׮�����|�M��������H�mO�V�k��+X,��!�S.J �W�w�������Ep�R&���_��?��T���ȧh����+c}	�5c�
�彗D�n�k:?��[�n�����_�eշ�vջ�:s%���}=Q���%������@!�B!NkÅfa�53�rpW�-EtS��^�e}|d�V�1�������?�D��_S�N�t�t���k�Կ	SSS �Rl߾����	JD͓��D�[o��6�3��8��c9J��;�LW9����ִi��Ԯ�B�{�<3p�:���N�LA����vd��m�~0-��/�rJZ勿|�2�mۆ�Q�����;hinɶ���n\O�f��P=�4����u��T�����K ��+����1��w����� �oΜ=����-,J���;b�R��5�AE�J��d}�_�_
a�5��y��@�A$����	��V��eX6KBʺG��Jم�9�v���t�Lb7���Ƶ^�TC!�Bq3W���3c�՟�"w�)�Ic,/�"Tҷ0Ƣ�=:z�07;BT�UC��[x�w�H$@!$��������x��@��ٙ���;�16�r�r�N��>����^3L�h�U��\�а���wo٦�ֵ�yo��!34�ĵ=�XY^�[w:���⬮r)�\�D�awc��r�|��5i�/^�Lݾ}��@��O>�[o���\�e}躶G��36����{��^�����M8w����!�ē={����]�~��-��N\�����Jsm�B�h9y�$����������n����}�� _UM'I%�?�$!�B!DΓ�j�:�����=���Rr��1���Q.B�B�oܸ���v��̀���o���Sl�ĕψq�|��x�W����B!��7������� �<��n)��ҥK�5���߷e|l{ _[W}N���-�6�8�ч�0�6#�8���n�۝��P�9���n��#I�8��ݹ�5i%�U�G���"����Y鸶[�T�sW�D�n1,����u����	�}��NNM���C�@?!�ċ��f�:{_��ƱGo2S.��R���`]a��X��y���KÊ/l�Ŏ���OOr	�(�կ~e{���x�ee�?N��a��%��ֺi様�'�B!���H���F$��������3�R�k\����]���j���؈�7o�?��?@���Y'N�=BT,,.���'8��ݽB!���ի���/XZ抾D���
z�w�D�����$�q���S6�i�wp�isU�>k�ܓI���a��w?P��ˍhO%��\nP5�C+A��潅�^D��7^,7�s�N��΂DC���5]]UE�vG�b�J ���b��n������B��m|��o�νo{��;��G�.?@P��f�����їD�n�_퓇2����oF�V��>v�O��;Q��-Έ)G{�M�0,ն��ۄB!�BPײ���y��mm��J�)˖�TW�W�U���v�a�%���_@�aue��$/C�xi�6�ۿ�== �/<���E��/�?~�D���F����h�홱��9�E�����؆u�mY�ُ1�7�����q8��MU�Y:Eq���r�Z"ws�92����{$��
~��,$!��ӟ�����|�G��\�%vmw��+˵]���}���������?������B)b9���!�v/�!��#���E��+�8ߗ�^Va�G���,��@���ٳسg�g��tfȿ̠�s�}����h�zgj�zc��B!��f,ьF��[���m������].�Uó^hi+c�B�V�߾}�6mJ�I�h[���He�������701>���9B����x��~|��� �1��|�$:�n݊˗/��Ԫ������0Z�����f
ߝ�*���c�?�Ը��*�>�G�����ݛ�8;c������w!>���vdȄٓqKZ+��7ޠ�=b>��c9z4�8�����rm�����@p�:f�?�z9>=�S~�� �-Ǐ���,��MW%����!��*V) n�%"�9qK+��{ih�����<|�	j#��V�;�s��i+t������p�#;�=<C� �7�f����{�^�VK��ƽ�ݍ݉�vbw^̾x���b&B3!͓v�Q�>�eZ�k�&	z$  A�{W�ŭBUefݬʬ����/�jԭy��Js���s�)�d�HK*U�x��!�B!�D�^�6e�H�z㏀k܈�5δ)�R�m-&�1�'7���,�1���C��>����悐H���%�ُ��}�w�$��(iiiرk'N^���D������8ǁ|���4�2o�.@U?����^1���|,�K�W�Ⱥ�Y(pw����/n{ج����e�C_|�"wu�*�Ɛ���'�P=��6`Μ9����0�xX^�ڗ/1g�ܘ��]�M����Ǉk��\�Ip�v-=�=�^X�7�x��� ���EE(�5%e�Z���H��vӱFk���<c�v3�{Y��v#���x���9���}{��i!a�FLL����Jj���dc�IS����I�B!��ȴ�� w^��8����l�K5�W����A���a�%&���g �QQ��wa�u��U�ܽ�_ !�gٷ?.^/�#b�G�C��v�ޭ���6'�#!����7����}?+j���h+�)��)��z��Y(pw�Gi�E�>�c���Y� T��Ǥ��$�$I*' j�|̉X0Q��g��@����;����o���=�M"n���Ʀx�˖B�k{<b����b�Z[�|�
446�it#��X&M���;w�ҵb��>bM�nFDnu�V"��v�ۍ�	�vQp"αc�_��l��xc��n���i�*�2���v�����m$o��aB!�BH4��S���6\�O�5'rW�cy�5ƊD<��֭[1c�<}�����Ԍ���@H$:��PS_�U�V���� ��k׭E��j���h4�֡���9/^�իW;*\7�����:��"R�P=����V}����fL1��y�fL�}yUKF�B�*u�* tO��v�!�U	�U�b����`6~׮]����o*)F�˝��p��1LKV%µ]���wm�k�ŵ=<ބ�τ Oߵ=vQ���*�ݘ�]���<t������!��� �<|�.߼&�>'�>�8a�nl�&nE۩)��4,��v3�CCC���q�<+����is2>�9�f�T�d��2�Q��1����HB!�B�1��fb��|u(�)�b�(�+���C%F���˒��=�>���}����q���rl߷�D���gشn=�͛�/^�BHbBٔ�t<�k01�x�#�r�С�չ��x;]���5�Mj =J��q�F7X?�"j�{T�{�:�T��Xf���!��d����^����Ny���U�N�}j���B'�ڑ�mn�>�+V���r�D�����W���9��=�M"n���#��wm?�!��C�jU�gY�� 1�����<~��N�'���O<G!�~<���]w���X����ܛ���8����}V?��}�arrr|�&�p�j���w�M�,�h�v�k��e���-�`*��S�N!�B1FI� �e�M����\�C�?��?+�*7��K;̚�Xb����T�ėښ�l���) $7�����{|��mmm �����0w�\�^B���܂���d���2�j�ڹܡv���Z&V�q�WeN�4˒k|÷��l<l�s�&_
��v #����-�*JVE�K�G��{Ff�8���}�h>�}�(pw������������E�Y�|_����JodZ'�P�=��F�tc-�l�[v�5�i׼�ux띷}"w&�	!�^v�ٍG5Ot�>"�[�{��3u�Y�����0���KkS�ڱA{Ճ
gٿ���k��?>���KR��c��̩ ��J!�B1�Ǜ�I����d�f8������?Gͱ��3Ɗ���֬Y�%K�����9*�`��� ��._ġ=������!�{�:�G�ӟq����γz�j,_��Q!��}��Ǫ����FK�~�K'��D�pR�,x)n�
��N��姨�۵bwY�<��A��H�j<�1���ѣG��}��\��)����K8z��qm7gBЦ��.�í���b����q�C�h�hÑ#G��矃B�=�]���him�%r�]ۭNr���| �Y�c����(���z������ ��\߆�v��]�n[Ǿ�`eG�� !�B!��ù����3��&�1�7���R�n�^D9���1�[�F������a�?~��׬BNn.��8�]������>�]	!��CZZ��ۋ�Ιz�"���N�*=�Y�1�'��v�e�ƾ�q���h�X���$����I`�06(pw����lޔi��lS�u���4#�d�li���Zwc����&��Ν�6�ڵk ����w�>Lʞ�j��k�,����7k�=6bl�����"� ;v��M� �_���
&M�Cy��`������=ǲ0�L���=��d,�X��	�c�?W�=q�iӦaǎI�l�z�����1���&�F�I�op�m��={R6*�� !�B!�%�#؜y�(�&���ci�o�d�e4> p���7�d$�:����A����p�z1:��'O�BH��I�:{��e�ST�>���IOO��s�U�n&^YT��֬�l�^�m3j����,��vǘ�B���t��#u�%���jS��91Dsc���?��b9�ÇS��0����z�
�8�{�k�,.~��&D�m��H����v�z7�'tlooÌiӱr�J����BH|�>}:�/^�;�K|�������o�F��ٯ7�,K�v˓��$J����sb �r��1ddd_�A�K��c�*6�I*�x���fܭ��Ҹ0�e3
f�[Oq;!�B!�m}#ȟY���Ni�P6&��C�X�E��z�@���y�E���F�\�t)V�^��w�8Ǔ�GX�j%2��@�zzzp���m߆�+� �_�a坲���
���x��	��l޼�gώ����p�5Cm�r�^�6�6b�fl��o��"��Q�+�;LIS
֤Jfo踸�;a��B;1xn n�|N2�1Ĳ!p���'tR��(�??��۷#''�� ���!�iwm�d"�x�}����D�eA�M�{�n�6�*���	K_]�;kjj@!��yyشu.߸�{����?҂0�L���=����cEK��g �"��9�����h�7��D%�Bz��Q-�P�^�:$
Q����0���lp�AB!�BH,��OW���:bw�R顱����^�Okw��.#-��X%%%��$�exh���ƺ5 �(ͭ���?k׭��;w@!$>lظO^֠�����q�#����=�z�pݙZ�dRw�=�,�dq=c,��#�!v"�G��B����wy�}�d���9�EZrP{�Dr����KB$֍��DVnn.8�O>��9���q�����.����n�/c���gM�k�� ^��a���>y
mmm ����8p� .]/��`��}���/�"�޳L	����k�o@Ow7���Y�+V��K����H���m�)$j(��*!�HH�r[����sa��aޭg��B!�[S�T��+?G�zC.��0gw��X^�9�w�cEBoǏ�w��]�#4q�G+���אEwb��Ϟb��7�l�2TUU�B�5�����A<}N�#b���A�|��Y


|�H��zN�e����za�M9��d���7깷��}yW}��.��=#��E�a'���=�8/uc�$���~'����᷿���c$����Sضc������V\��qtm7ؽ�X3�?KBAo��*V�����>CGG!��#--��A���Ȅ����X���k�õ��q�χ�.B�+V����	��h�����>��M��
�V|w�%�����~Λ:��B!�Bb��u���ahpP:�Э#*k���X��|�L$�R4�l�<y2��ۇO?��9����X�v51ý�R�ش��ݨ��!��ؘ�`>�f���;7A�Y�^��{���&M
�v���>���s���wc�B�����xQ��
�]��L�1�� u��;1h��nwc�s�7oƒ%KP]]��=��z�
����{�W��k�_-�nr�k�?Ԙ�ݺ�0��?�q: ;��ϟ���c��>�%�!�CL�<r�(n������$"Q�k�p3�^��Y�I/��L3�q̿|V��.��_���q��!G\ⱏX��$�cb�CȉA�Z�4I%�{��e	!�B!V�)�H�tըH.��0w�)�̓��^n���)xx�P�j�u��A
�]@��]�<I�.߸�};v�r6� �b�3f`��E�2z=%�,�}}h��q1�uC��bm�5>�0����y�D���K5��[�m8�������a,����aT�\B]�@����
f�!~��Ē��YN~��➥qq�cݵݪ�ݲ�\1#,�o���=�|�u��4'�/!r띷�O~���^B��o��'p�����5�&�>b|��X���@��p�/qQ|/,%I��Jt��?�?�T����f��B�v����&N� �B!�X��/EQ�H���jbn`,6�	�uV~��'�1֎;�`�<��9��|.YB�r��>���!����B�1�M��U�����AH,<,-�{�x�W�n�:�E���G<�5�Wcmх�����h�KV7�����އ@b�w���gLG_k��ҥG����$V����7'���}�{q��{1��ߧyG_�K]�#�=�?y�a�����u���c�x�M��w���� !�����>|w����G�n��#ք�fb훸eQp/uV�nf�/�>GG[;222@�C��B�n&�H�����S��L�J����x�"����=/� u/�� !�B!�%u�845͜)�v<3��F'�P��l�e6�ic���4_�����>��T=x�e+�#�.�$�_��;��z�Utvv�BHd�L�����Q�NbF��?��FF:%�Ns��	��-L�b_�YG��S�z�\?Ԏ���\]w����t��S�j^M\B��$LI*�L���.�7e���n��G<Y��s�b���x�"�����slݱ�Yِ���F]�ÿá��c��ܲ��&��8pm��3����A'��!΄#���GœG���R�Z����d'3A3"r�����'����`Μ9�����S�$��D���&vW����\F4c���"D��B!�B�!�F��)����lX�*Əh�����,3�R�b7�J�(�f�������~���.�Utq'1"��/._���{q��	3z!� ??��n��ۉ*J�3<L���dff�СCq���p�j��6��=l�x�`�P�f�j7P7̙:�&��«�K��rG
�ͻ1��F�n��T2�����#��D��}9r�w ��.\����7[��ь�{��%����>�X˂6;��E���_(��^���o��6~��o��&�����h��P�&�>�lTn&־�[�?~��f�����>�v�<!]�,��6�x6��2�����ɕ�k�����t�U����L'B!�B�u���=Ҡr��C"�%K�kW�JM5n�����i�������vK�,��͛Q\\�,B���k�"3+��E\��~yGĹ3g���B!j&M���w�ԅ/b�"��+�@�g׮]�={v�'��ݧR���Z[�Yo���=��ڃ��9`��:����0�`:zۛ�UV�Ė�j܍A��/N$����;�����A���>����|�D��܍ݨk{�
~l�[��$�wܵ]�5~�fD�C�x�X������o@!���;��--c-�����eYDn��e�����In���@�;�н��eӏ;f)�V�v�x�b3���%�ԛ7�jZ'���$wt�R��I*B!�BH|�Y7�]�)���?�OQ,�_c,_@�^	���=��N������V�_BbA\7??w�����@!�Ovv6:��ϟ�=?+�%�i>�Ę��ѣam��cmsbZ���u
ջs���5C��g1��vχx@�����E��^Z,��Eqc�o���ɛ��S^3�ѝ�H�X�����/~�؉��	!������$F���O~�W������>&O���P[G��e���g0'�3AA[ͳ�x�|������Y�������756���I���Ϫ=�����:;;���S8�p�ɲ��>G��]U�H0���I��Ku�p�;ݿpA����mN��g�ZWW���w���n��_<kh�;w.N�>���n���L%ikknAEY�$��5Ȉ�|hh�����}Í������*M���������6<�|d|��M�ZZ}c���\�k�}�aY9i�k�S�ց��B��-\�0b�[� ��>B9)�#c&Q5���DLR�%��\<���B!�B�E����NGog�����M��#c�~
c2��ݯ���?�3���@�%��>)'�Ă�}q�<�3�N�B�_����~����cuM2>�����G�A�gƌ>�d���ǘ�v�x�`�Pk���F7�R��s���@�3���.�F�0�MN�]�<Qnj9��DKq��B<����7�|?�яl�U�����8%v����I�����~�k(�2E�.���/���g~���@�x��x���A����Bܾ{�^��5]#�Bܾs�n��j�k�����.^����	v���:�����N�BS!v�9s&�����X�`�B��-Z�H�����m�ԩ����gw����&���ů����.�5�7o�#����aڴia�۝�����������U�����"��r��@OW�o2��ysUǤs��&Y�qq�㇕X�|Y�8�n�=ߚy~\Q�E˖�}�ZĽ�l����z��7�|=88'�'�o��_�ͅ{��-R|<���86��KT��+]�ck]a�d���]�WX  �B!�ďo>2=M�b������*V���b%&�[1�
_E�}�V��ǤI���[o�׿�5�D�E�NM�w�K����6�G.�~��Ήk�=]����Bz�3����v<��v�o�����C_�#�;�مA���|u;�͙�ǌ��D7g�`��N~vq��ߩ�8�D�fE���ɿ}�ϩ��g�E-�����}δOC��N��ă�0�r'?{�������@<�4�N�1���8u�{��T���T�eJ�kH
kn�g���rc,��WR7l����.��;�;u:��[�&�B'�|v��p/��Tcn)c'����b�,I(��b�m۶�ҥK �"�O~v�'r�㕈\�nx�b-��M�����-�M<D��_7&�[p��ߏ��|��������'>%���Ğ�{Q�܈��F$�>bM�n4־�H���f9v��#�T��J�N�c֬Yؽ{wB�Opy�"1h����OTI\%����1�x�����Z&�!�B!��v�5�q��fp�S;�[5�R�����D0�:q�>��c[�s�D��Dw��n�8@��\���'ǭ����ȟR0:�wȨ��ڰaE���G[Kf)�B���=-3�֯GZjjPl�H��)��D1�͙����3hr�͙�9՜9�(d��/_��ٲՇ��{q���O��H���.����/�c��E�'���-�H��Lu�z��gOd�BH��uճ�0��/�Vp�K����}��~�1V���s�=�w.T3T�Q��1�2c�%3��w�>���
�]F�'�<���'�70{D2�Ŀpc��%n�#ل���w
��A�����0s��O�H�����kT�gYDnB�������Po��E�v������x��i��W>� ���7�$�!$шg�����Z�Z�1V'3���X[�#���m����H�W�> q��+]��7�|T@خ}#4&6����0�N4׌ս9�@!�B!�σ��������A4Escu�ݱ��v��}�c-[�7nĵk�@�E|��K�cˮ �
���y����|q�#4Bq
1�c��=8y���Pz�$.5Hba�5��q�ڳ>��-��c������H�ʺ��u���i�9/(pw�j�ؙݍ!|�A���	-Q�h���<�"�1�p����}�۷s����"%�"�ϟ�G|���"������n��ܲ���=]�#�
��Gϟ��w��~�{��;!��W���#ǎ���J�����o��C�v�N��Tzx��Q71B�0?~ܶD�'\*7A��U�1��2�è�K����B!�:S� ���0�
M�U��KV��#�B�X��"�����
c,
��A͓gX��uL)�
B� ���;��{����/���B����cۮ8}񼭫Ӑ�CKc�^P[��F��mf�k[<�kfjC�P�ި�=d�%[���0��z��n�Q��=y`�0~P��2�G�7w:�:[�KHg�x�Dd'�4Y�I��<��#���}lB,"�U����@��֍�س-^�x���k<֨�]���U���vƙ��*�4k�%�?�����?2aE��g��G��~E9:���޷�>a�n�ν���ͪ�^'�i�z<��}�}x����I���͋�f���LK�GNRi7�n�J6F��3	����Ƽ=!�B!�D�f��2�jW8��]5~�*�6c�hE~c� ���1����x��СC��w����z�)�[������k���p`�\�r ����ԩS�e�6��������xp�v	�;5�]�v9^L�˻�
}�f�*ǵͱ�c��� n��O(pw!m��O��.�r����'�dN�D�:��U]D����h����\��%|�_�?��'��݌��M��M��]۽�8����nQ�nU�3� ��{����'x�����Ą!d\!���@ɃR�h�V�zIv�v�����Ǔk{�����3���n@�W�;�fv��ٽ_�{����х�z�*��^�|<e�A�Cj��}Q�N!�B�����/,B_wG�^u�g��MV�OM�P3��� l�ceff��Eݐ8O݋Z4��c��Y �*�y��8�{/n_����fB�x���k7����gm������5hnlqo��6��CR�d�Z96�dm��@�z��,���Z]7ND�����	��wr�ދ�Y��=�|�"x��$��41#t�_(�N��O�$�Ѿ�Ν�={��̙3 ����c�޻�UkV�^�um���ܲ��h_&�tm������̇�U8|�(Μ<���6BH�#�m+W�����>�{�#��!a�{��i������6���,\�;w�t<�����;�skfPjQڄ�j�\fp,6�2��Nè��핓�	!�B!�ѝ^ xZC�Bc,�8�;6�78�	:�k7��ϒz!����X?��}���)�y�<fZ�C�q}<}��n߉���h�X�2�����kW�&�/Ľ���� �@h�1V�k~n]��?F7Y�ea� K��sPgn�%�`��|>��m���������>�f���=����y��jڵ'�p�Ԟ�A�g0����,nLB�9^��:{�3��o~�+�����sF�&D�m6	�-����(t�*�7k������I5>��KW���KBH������������g�DVV��ݾ�����5'��X����:+X����[|&v!---���.�ݯ�$KBA?I��믄a�A�ds�2�YY�(m���B!�b/��S�.-4>���YR]1�״)�F�>���-Z�l~��y��hk���O�p�����>�{z�C��ւB���3�\x��2�'�+����<�9s�D��K�ﾌ�{��G0�VL�����by|����zz���ݥ��NA��Ew�G��tI�~1��+^+/����$�ō�-I(3���%K�����yZ�[p���ڳG�M"r��6���{\���&�k��}���'��q�fL��B��RBH�1}�tlܲ�����s�(X�	��X;~�X;D�n�|K6е�-��������`u�������n<Q%GZf0l�-sb�oƔY�42QE!�B�������K5>��_���Һ�̥��XƏ���ޢ��Eܿ]�� =��?�_��m7#7/U�U ��de��#� G�k��-!�bhp���jS�6���g[<���pիmP��c���jc,o�q��n�?�mOG@�G{.�����A�l��B����8�\VA��6Y%�I��%�G_a��I(#m����{����m��᷿������h5#"7kB�'�n�#X��+ݣU�[��b�~O�?��EQ0� �/s3!$yX�t)�,[��7�����9f]���l�-�,
�a����"n�������(,,�N��]����*�P��u�J_�.KRyu��a��&����Q�)Vʠ�;!�B!�~z2��v����Fc,+�ݽ{�����ӧ ���ׇʲx}�*O�o^����M[6�Ƶ� ��dc�ƍ���͒; $ޔ��bp` ����زe���D�C�S�G^�Y� +�S�Q����q;�q�w��50�ܹ3��������_^=5���C���\\���$2	e�~�ڄ;�~�����8O_?N�:�w�v���0'h3#�7�=��{]�-�e�g�����ô�"���[�㧟rb!���Y�ٹ9�~�V�ͨ���}Ą`�L�����{���!����_��a{ .1�.��DL�5ow�]��:	j�T��������^�8Z7IHP)��9��(��r8!�B!��ō:`c�W�����>''�]���4�fcb\���|�T��c�+K1)7�ē҇�X89�M�fHI�s˶;PS�5�/AH����FuE%�{��W�6�X��5?{D�!�,���ߩ=\'nY�&l���7j= �w�8��O����_|?��N�HM�8����)^���T��3����D�{����<ߒ�?��A���3g�}�v̘1C�nYDnP�����x_�tm�EDn���ٵ]Fsk�s����C���;�B�Ȗ�[�34���I��#���'�eJp/�G��6q��� ���;v`Ŋ�LDّ�
806u�1�иX�̠�Z+
�h&������ENCB!�B���;�ɋ����]��.��V~��yB�T�X�7FSN2�1����w���Cttt�8���������[AH�yV��=�8v�8N�<Ś!!��ddd`߁��q����A�ܿu�7V �@��,V~o�W�⵲V��������(3���L�u'�KVV�+���j�ws�փ����ur����OXɜ��5#��&��PF�I�v���~�A�K�����_����#�fYDnY�����{]ۥ�1�#��u����C���W?���)��\Kq�Q���C�z�-�-�6{�#��D�v�G����:\���.��� �;����1����!a{�g���e���#��x����=c�8>$�B!�$�o2=-Q��'�j�򕮴�v��Ke�%q��7Oc���|������A����'X��2N+!񦥵�/���c8w�,zzz@!n#77����]����A�4����������#''��Q"�����ۯL�ѸeE�!���F��ZS��Yu��~h2X7�
�]����Sg���>b�J���'���a�����8�zÖ�H�$�D����o�>�:u
�<,����X���w����ƃk{X�)�[���iFh�?�wE>��	���@!N������.-AOo������{�(����#Bw�����OU����K�b���I��2ۗ@��
��D��I߽=4��q�,c+&���
����I*B!�BHb�V;��y)a�LE3����+]	S�ڡ�M�E��<����������A�G�ݹv��1=�#����/N�о}�}�Y3$����ӧc͆u8u��y�;ㄒ��A�Cvv�ou)N��}Lr$ZW��C��[��Ħ�𦥥�z-�vA���y�7	Eڂ�$Aeĝ����I��Q&q��dIBY�_�N�>�Pa�̯~�,��ː���h5!"�,h3ڗ5�^,]ۍ��*���
l߹�e��� !�8�̙3�q�f߼���g?����k�E��)���XcǤ;�\�ܽ~�Ͻ.C�*%���̉(#}�Ƨ�ve�JyA���uAol�ua��2�G!�B!��3�E�ԙ�io
��[�9��;��"#�/^�={���ٳ �����% ����乳صe;�rs���cB�ӈg������� �N�+*����:�9s�8^�K���\���\+��:4.�7�RQ+4�J��I��0�b���;���%-�k����w��ܣ%�����;Q��x�NBE�j_[�l��5kp��]w��ڊ���Б#0-"�$n�&X��ںQD�V����x�={���,��чC����hV�\��sg��kWl��X��3u\��Y^M��'��cǋ��i�c476�����;v̱���ɱ`ZJ-l�:Q��k��v���ݣ3�\=��nc�h�t�!�B!�$���y���'=]];4,r���2�:�{���z!��Bm���.����p>222@��k�ū����X7u
�ܢ�-!�96oٌ�����b'��(�{�=����h�dqf�kw�����M!n�]��v�&�����b{֗3�+��w��=�2
f���eXaݣsb	W?�C]��#:1(^+/�����b䶄S�m������?���QTT�j7%��E����`݌ͭ"r{�����g��x����yy��W?���)���@!v#��v�ٍ��N�,�c�c�>���wjJDn��-3�e��!Bw��]044��;% ������ɓ���$t�ǅAo�_^0R�J������T��&Q�?u�R�N!�Bq�/�p�0#�=NwL��*ꆱc�j���Ac�H$��=Rێ;|�eee �  �Z�i=��;��0w�<|��~��BH����ۇ��>!v#&��!q6l��u�\&>�_���S�5\�e�ʺ�n�Pn�5�̬,ܩD`lL��I@EG&�y�GO��,c�Ɛ�
$�:��׏�,3�&{�6����uuu �@<D}�?�����l�~�,ڌ�]��n&�k���ѵ��n�а��=��8�֛�|�2�jkA!v�������Ni	�::u���V��-��V���#�c�*�wZ�]P^r}����&D�Z�e�I��D�ڳ9 nW)��^mJ#b�}DW"KT��v�N��	!�B!N14dO����z���Rǹ�t��HĦ�b6Ƃ�f�+�E�ь��x�wwQ]Q�E˖�`�b'/�j��юc'��ʥ�hmm!���ԩS�e�6\�z��|$!����Y�w���������g��иT�0 n����uEO��u`��B��]8�F����$��q���axpP:$�r��U�%!qf�z�'��Z�$��"�Hm����dտ�˿����wKP��._.0(h���n&֭"r�5a�u�'�mW\oVWa�����b&�ܾB�7���Ǫ��q��˄�V�#�'~Y�'�e0N/v����l�@��Jwq��!��&�M&�H�{ ���:7�cTqr14N��kU�uΞ��B!��7�=ãc�C�X�՟哂�b��i�u��q|�{�CSS�;��;Wob�у �nz{{�ǳ��e�F�44���
�b+V��܅�q��Y��Idb �gw�����e,X� ���O��_|�
d����B��x��[h��0*��G��+�	�I�H�tx����$Kss����. ���6�̠�cPaJ�'���}��_��������|�����_��A,ڌ��ڮ�}�D�H������>m9�3�O�����o؀Iy9�t�N�U�E���8�f�\ۍ��t6��nHݾz��3�!�_�����dqF�b�?�m�ra���"'�d	�@�*�p��!�B!�8˝�A�3k����-����X�6co�����'���+�{hnlD͓g��x!�q=�z�V��;v�ĕ˗]��%��ĳ��m���݁3σ�D���- ���?DzzH��&�{��d�uC�M-n�b�*�Fwo�7�
bi&�O��Ei��vC�{�PҒ��F<a'ˈ���������� �r�^��()1h&RR�/b��VPP�w�y?��A�CkK+Ξ9�c'N�tm�V�C���#p��ܪP�L_��S/��Ѹ��fL���WG ���?����+b �w�>�l�CՃ��s"�k���_�E䉼g�ӋuZ��b���Ghn�ۘ�عs'V�\�x�I�����jq{a����D�J9�V%���8\0z� �B!�'�򔼙�4ר풉�ac��B~d�h�X�#S�<���~򓟰>�2Jn�¬�����	B���
L/���o����g���B���L'j�7��AKk+I�}���.��(**��o��*��5G�bӠ�*k�Z��Y�v�)�:�Rڔ� �C�{��m����S��nԉA~�z��jf�A�����῀(�S\�p����׾�5�����e���$V�]��s愽g\�f\<h�>�"rsBI#���M�k�n1�3��ׇ�G8t�0J��Gee%!�,�f���-�p��m�Ȟ/��Gd����b�pm�߅��J�v?(�S�.ĸ㣏>
k��9�	;]��*�vu�*z�J�ܮ�T�������B!�B����t,Q
�u�a���f��]%nW���| ֕�RR�/b��6e����������e�)��-�@H��Xg����޹y��� ��X�3w.V�zg/]��0s�$��ɂC�� �BL�����vS������B�H�uB���R�Ľ}dă��i�={@��$�=m*�=m:'Md���M���*��ܕG漰�,V��={6�?����7 �A|������_����k3'h�C��V����wZh��߽�Ǐ0o�"��lN~���zL!FX�a��B�ɻV�#&��c���g���uZ��a{���o�D��]�Y�[�nE�8KDYuaP�ݵB�p7�do�I+ɘ;�p6�A!�B!��Q�kLEO��K�V(_�9��]��]�f�ө�j�,7�#�Y!0A�W����\Ɠ�GX�x�fL!�b`p 'ϟ��u�`�ܼy�b�l�i�f�>O��x�$���:�<y�.rss����#%e|�ڍcƠ���b�L��;�G2�ҚQ�O��gO�K�'�/F�'/E�̠�Q.������BȍAv���Ag�1*�3�L.9��.����1̙����ӧ�y�:�l��Z�v+�v��:�	����õ�(VcM�������|_^����zB��y�سw/TW���$ª�ܠ0�L��ޖ��E���+W�G����5O���1�Њ�$c�����̱�0�O��{,5(OT��#{�g��!�B!�;�)��$]�Z�W]3��*q�3o�%�xʜ�̗,��xc=z���oA܃���}��8꫃�H�߹���g���c��aOO!$y��]�UZ��f:���#�w�qr�y�w0mڴ����b� ˨�=��9�{u�J��l�g��VL���IDϠ�
g���^:3DZ�OKsn�w��KR��D�(��jwu�j<��#�-[����ǩS�@��'��5��X���U�Dqm׏�*�4�+y�D�N����(�|��֣��/^!�hY�|9�,{Wnݐ��`�>�3���NM��w����>�$�y��� ��W^�5ܓ8���=.���.pa�*I��P��_��/(n'�B!����^��AX�=�)�gtKS��,Ky��*1�(�!c,_%1�'�1֧�~Jc,���֎��X��� $�445����m�&�44��� �=����-�]7�Z<q��J����.233�կ~U����2��ޮ�!d��F�*Ǹ���X�U�[jj
�׺��?^��=�x�3	3��qcО�"i����|/��.]zP�:D
��qɐp�������Ӯ,Md��������ڨ��+m5g.6a��^㟕���c�}�׾@���x�+��_�]BFIOO��{��ՁKׯJ"��G
���&�>bQp�����(/����Nw!��(����j�ō϶`jʰ�]-r�sb��̠*Q�k�d	G�B!�B����"w�,��5�L�t��v�1���?&x_+� +P;L�G`�4Ǣ1���bϞ=8{�,��9�� /?�$q���W�,ŁCq��yB�Qغmj�p��y����,�d,7"V�Z�p!R\^���z!��+��������^2��G+L�m ���u�DA�{�q�n������`����L��=�DMU�R	&���v��]y���q��h0�%����_�[�nEqq1���u�&�oڈ�sd�.Xw��܍�{��;-44��>����щήnlݱ7�]�s!�Y�fa�捸y�.z��4�Z��X�����>bQp/u�}��*&�܉�V�8qnOR%ąA!n&�"�۵n��=����6Q%^�}\�!�B!������(R
�5�X�L�B����J�fGc,sm}����W�&"�\�s�v�B���q5j�j���A�=u-�� ��ٳgc�����������ϯ��������HKKsĽ�i�{�`�P�!�]=���y=��a+>k�uO���DA�{24i<��ԅw:��6z�S��cnju�*��+�,�"%%�NVڄ��իW��r!?��O�������3�bM�l&�����E�����~ݚ�эn��L���g/j�_P��[���3!d� ���m�oz*.^�M��*"�����5�v�2x z�f7�G܂�7ݸ|�I*�"�����׉H 9���B{�
���#v�NbJ7Y5�^^��V�\!�B!���[�CxgV���B�B��\4�{�A�ܹ��X��6l؀͛7�ڵk �O=ƢW������é�_`ڴ"̜1uuu��#B�C<7�۰i�8y����y��-M�|�F�*Q+W�tA-Ͼ6-�1�N�*Ff�5���>�[[7�5���srsq�nJ�,�
ܓ�[�X�ꑞDF��*���RS� xe	+�ɪNb��$g�hۮ]��v�Zܹs�]tuv����~�#����(��(׏�*�4g&VGi�H�v�ۧ��]�mj���D�Ç(/+!d�3{�lظ%�eh��м�ዛ��`�����@�^_�"�:)nO���������V�1m�4�����9 ��;����1�9��O ,Y�NP��T�x��)y�J5�k���<��!�B!č�:�7w<-�U�QE2����M��KE�ʣ�8�B�1���ד"G4�(�y3��¤�1!���I5�L���Ǐ�ڕb����2q(**¦�[p��6ZX�!.���ew1��Di�dq�-d�eDܮ�#�̟euC��6l��6�L�z���$��˃������=l�H�tr��	���0�wJHuLX�/.�3��III��S�m��o~�����W�`���X��rU�U��u�]�qfbM���n<6>!�o���
3f��{�_��S��=:X ��?����];����W�H"��G
���&�>bQp/�ݕ����щ���d�V����#///�:Q�[���GPЮ�h�*܅!���ޘY���2��p�Xy�.�B!��r�)+��|�l<$��׮�po7c���Lc�`�pX\�f�޽�.�q���ؿ�8M{{�ϵy�u�N���K���&!����͛����;����D&���cxh�}�U�7n��"���m�q%$��fo�ڡ|�T7���s�(K�jo6���$qP���4x� ��<z����KT�%���w�M<X��*g���X�7��T��$g�h�޽{�~�z�ɪ��U����ɾ����?���dggc����&��ScF�,i5(�.�}�}�b�pmׂ��^C}�[/������4CǪG�BC�g�}��8�&7����{���1=�y�������A������>4����N���=d:��D�ۋ��w�'?�ܹs�_0eU���^w,^[}oD|�~�G��zrL�"�'3��x|�|˂{���H��Y�C����^�v1���;y�{��\sF���嫾���YL�Ϸ����|�AR���+���x�0xF�v�dU`l�5e6<��B!�B�͋�al]8}�ac�Hc�HYF����BE�04�U&�1����K<��,!N#�7��F����� ���������B>v�n�D[G;q��h��qb\�o}+�M7�ڼ�-$nW*��Q��d�MS/��#�b��?�O���'�'
ܓ���L������4�D���:2DXrP�.�I#P��ĻM�ɪo|�����D��p��X�����I����_��~��_a՚5h[⩽�c�]�BCsar�_cC#���W4Y���s>�&�(�_}�&�F���C_���Ի5�_3����f<,`h���f*�;�|b_%��1);3f�D��G�������a���)�K�S�&�����	Ŀ�D�ۋ�wuu9ҿ�]|�E��e}?~�i3fh"L\Ǥ��~����������1ԻQ��{fwW7�^�F�ܙ��V��������z75�J�w���A��I�^q��_ i�o@��uю簀��)��8��dF��G�½=???�z<��cuaк�k���y�0q���0�f�]K!�B!�5e
2=��q͈'�_Q�
�+��cj��zZ@�~�n��ٶo�>������a�W��\��_[�I$⻘�����Cff&2�2�������K̩��յ65;ҷ0g���v�'?������ ��.��I�c,�� s��CYi��n�f�:V3w'����)����S�]|n'��-��N���N|ޙ�f���?�����z�"����;��u�H������<������N��N>ߊgz����/�v7mڄ����ihk���HY���u@U=�#��j��U�Eݰ~� �&
ܓ�!�Sfb��VZ��s�S%�Kj��nR�;��ɇ�9�M��G��x��/]���݋ڿ����i��x��C'It��e�{`?fΜ�{�p�"X6�b����q�f�XSn���vE��7o��˲k{�����X�h!�Ƅ[�:��;8���nX5N�l-�����X��5�~�5dێ���_8w>�I+��y���)D�ĩ�����z�ԩ����gw����&��� 77ב���W��/]��[70���",ze�"��}D��:q�l���T��
潦�C�8q���xa�����X�u\$j��;0s����K�DQh΂�p
���E��uut���b�@�ĳ����IN ��k�X"�/**»�;!D��mr�2{h���'����n�:��'NC�S&�!�B!���쟜�.�덁d��ʓ���ͱ�c!4nK�1�Q�0����QRRb���b'p�o'��K�V�j�:ߪ���af!�"55ͱ���=-}b~v���v���E}����i�V4���EM�-����+8�����E.۩��^g���2�q�ϙ;��ǵ���ى�ӊ��{���D6��n�\�T�n��G�ו�ܷ��W8��}������ʱUJJ2��bkS�P��Ɵ��a�X^hM�e��X�U���6=�^�n��'1�Z��J���*wo�IpcP^ �\��v�z�.�nqO�c����g�g>7�Xl�^~��?�G��3_b������L��Gp5֦�jE<hW�����YEL��'���ǻￇ[7n�ٳg �����BlݶO^<Å�˒�����ucm���\�����	���ĳ����:}�


��'B�J�_m�%#�0����ܽ=����PlM��x�B!�B���a`R�l���E�J�4�X�X��5�Dc�KoGmr���X�r%�޽k�����@��8�w@ ����
��.Ƥ�I���C�CF-�Uu�8�@_?������t��<�^�U�cŲ�غu+.^�w�q�b=y�d8������0fMN��g�Y����_��,V0u��9�{����[P�Ԉ��!=+٣my��������t�ã�����	�����ֽ�<��F}����V�x�v�=_�����m`B����s��͛�����o�&l��K5cY=c��cfM1�h.�[�aBC�{S�:�����6sDof�Ȉ��.�!U�Ơ��f����2��҃���-vɪ5k�JV����щ+/a���v���Ċ�-
%%����֦3�N����	֍��r�]�](�|�ů��UkV�����܄�!�;v�@Jz.߼��9o�>bP�mUDnq2�~l������du�n���R�6���1Q���ߟ���^Ŧ@������ubso�_�L������B!�B��Ҏl,��)�cV~3��q��1��6����׾�sqO֜�x�v�u�߲	���Ux��)��ځ��V����B܍xذqr��q��u�ĵ�D����n�q/v���k?���ǔjc�`;�S#��)�>c,Ot��h5Ļ͙�GAw'��=�iB!�=m�Y##U�qii~��r��W�Ƞ��KP�(]��	�ɽ�*;X"(���r/�X�t1.^�{m\�,�]ۍ�o攰Ghh��5���j�}�����a���ϝ� �� ���׮��ٳp����$Q�Ms���u3���gY����d}�kkiEEi9�{㇩S�_O�v%�a�D��P�,I%OV�h�T�IޢM6N��܇�U8�.�B!�����i����KU7�3�
��\��c�Tc��v��A���?���L܇��<yT����A����_bƴ�8r�*<���O@q.����v�=4��p����z��U�O\�ƍ�}��q)j�ަ6����m�0�s�Dm�f���N
��O.,'�;�I��a��)]R]�D��=#�H�%�RG�Ґ�ٍ!,qHP��B�<�@'9�U�L`�d���d��9��[�S�H�u��<��{3��pm7J"ŋ���b���E\k+?BvV�|�-�|�ׯ]!�9DrJ�ۅsJ��:QV�#�����w1.X7k��j|B�D�{��q��˾{
q'B���$q�)����R��Lܮ��
�޵������� ^2VV���vK��@!�BIFZS
��i������\�}uDci��������!i�K����<y��o�!n���	��;�W_Y��Ǐ�Zq1���@q���l޺/�kq��9�v�)VSC#�;c�?��?��V,��D[�f��B��@c����f�W}����"9�k��aTƺ�SP���� ��ga��f�J�
ڥ��90|'pj��؄�])lW%�?�x�2'�V}�))�#v��wĤ�o~�����{w280�_����O���(n�n��Qpo�7������X{>��(���e�1etp��{����[���!$q��Ԧ-���َW/���"ߟ]���$�>b���b�xI&Jn�Awg�{E�)�I�ͽ=� ��ݱ=��gD#^� ��}t+(��gta �B!�$)�^xpdj�aS��C�HZ��+m�}/���$v?t�~򓟠��ĝ<,}����a��f*U���jlX���Y�Z\L^B"337m}�J���i4D����6��Ь��lذ۶m����6�b��$j �K^?Ԏc�v�J�Q��cY��8��uC'��}p�1�R�'�T�|!l�.3>���M[nP����]x���0^I�8MV	w�d�͛7A�I僇�z��vlGB]�-�!�7�k�^�9���X[��h��@���ڪ�X�f.^���.�	�������� -7���v�;���nE�nQ�oJp/s�}$�h����*�2c�|��I�|�2�`{�}E�JW��˪6�z��h�v�6��b���B!���dpH�2-/#�ڕ㣴�13��1V�+�1�J�.�zi�%����o������K�����ߋ7#��7��ANNv�ۋ��6ܺu+��ل$��j�*M���wn����$����bN�p1�����Ͱ�TW4ڦ���	M�0�qU�֯*��ca#���0�
�c�	�A(p�vc����l3��.��������P@W�.���$�HII�dU,�/~K�p0�n~��O�ʲW0}��`�;D�	�K�Z��vut�H�k{��Ok����{�CO._�ā3!q&==��؞_0%奾s���ĺ�[8&��7q��}��n��$��y�*�������k7$��a��L܎��֍Aw���pQ{$�B�{�Yٸ�bJ�!�B!�$��2�W1މ0�W�b�f�Km�%��+���X����5�@H2��ۋ/.]��Y�q��Q��/�
Є���ŋ���[v����d����hkq/;w����S�f �NUU/���V}6�ޮ��5	y��9(p'�����M>A�'w�̔��7-$r�:1h��&�$ɪP�&$�NII�dU��۷o�m�/_q'bɶ������w�Y��.�[J���`��X78���%�:�o,��1i��E����:^�
��{p?<�����E
�	���<�n�:L�9����QE���H��b(6A�,��6��G�!n���=��,\����+�O����\����bw��zS/3�	�q=х���[�y�4��� !�B!d��݃M�����ݔ1�����Jc,=���X���c�X���h��r��}֜�(�>�$��u�mū�qh��(�w��� �ď���c�����EN]��$�u�x��Ľ��poW2Q��k������aX�F�nt���E3��1��NC��8���a�5+�C��ɪ���tq���a"��;C��]�'�+�N~qJI��*�HV]�z���&���'��޻a�%��\*��Kpo����=�v�;c-�<�`��ء�!<z���w� ��|B���~B�#�߫׬���p�A*�?�[� �X���G�������H�RU�u/^��q��������lU���D�%>a�Ulc��["�ܮ��
X��#rU��p��]8:�hːs�F!�BI~�S��i���@Q�c�4��=c,��n�cź�-[�����r��K8��qdff��d�Ae�o{u�+8�~J��E�K�	���ٳ�z�4�4���s $�>߸\<�j��C�a�ڵIch����Q����]o�g#��hbv�6<:��(=�ag��}��=a=���iyfj���+_�A/9�"��.�ިX%�!Y%n>��S�@�˗�/`٫˰b�J�k���5��5Ｘ�a�-V�W#�|��B�~� �zzp��e_;!D߽z�:,X���Kq񪿸�k���ݢ^�����c��@?����K��ĉ��۹�p�v٦��$���1���fUy�3QGB!�B�8��fǦeE_�Yf����3��h�5����ŭ�kضgIF*���q5^u9�X��ܺ���&B�3s�L�Z�Mm�>a�x�#��W}v?>c,%�ahe�-D�KV3��N�Y�ꘞ1�Q�vaTv�Vh��k]�=P�>��Z��^��*�I�����'�ҍA�Ȑ���C���_��z�>Q��dIV��_�%Ο?���A�����	���?(�2%�M�D�Ƅ��q�5k⳺�m׺(U/���E�,nPݟT��N��&:;;�克 ����o��������.����^�b��ڮmM�k���v�`7���d@�"��y�s�&�����}ɪ ��۹��m^�B&`�sc����핊�#�6¶����@>��@!�B/� ��gc��ቿҚ!��h�5y��O���x�R����OY�C�WV`Պױn�zܾy��� �������Qn�g��Sd��M�Ҿ��eY�,;�c���q��/���؎�؝8��L���d��93���{���Ξt:�N:��vbY��K�}-IU*�JU��J��\.?�  � ����"���G�x����� 9���b�����D��+ݽ��<���X�z�Gk�ۥEvn�3�Ҋ�C)��)�v�g3�/D��� �D�H5+�`��ۢ��OZ0��!_l�A�f����]7i%��e�{<q����*7�G���UW]%94��7��_�����/��u�"�D��BGG�e2�Bl>8�����N	�������8�4����*|�s����7TTT`l�O�⦴�7�xf46���Vl߳+���2���Vbszq��JG>�z���br�T�;r!�M�7�X��vBj��Z��tdJS0����b��jZ�х�B!�R`���z�~!?�����X� v�1Vas`Of5�c�D�s��1����u�a��p�i���@I��؈�7nD�`?>ڽ� kH���뽂�˗A�a^���O��y��g_l�6�R�墢�^o�g��a0h<�sZS�@@�W�{w���������Z,vE��R�����E^�	��)��JrcHra�
�%y��d�Sɣ\o�_�*�{�=�K�3g���͸��{���Jڋ�����|ݹ&�bm
��Mn]?��W���0F�Fq��	����?�2_)v�څ˼�!E��1���P?�ǚO���3��v�1���,��NM��4b2�(6_�#^���ε�Emm-H�"��P�B,���gv��y�Z��yq�F�v�k�z^�ae�E0M�*���'1��T�"WB!�B)$����]2��I���=G�X���2�J���X�.�!��o�=}F��!ċ�~����|���108�y���BG)f�,]�U��r�@?>ܹU:V)S�ٺ#�@��	�=��.]Z&WV>�o�fR�����M������jf�C���
������z����ۓU���=��'� &79i��&�Dǥ|��.�v׳h�"|�_��~�3����?���˖a�����������.�wYh�/�ҍ�y��m�%���k�E_��rF*6�Y-n����Çp��,)d����K�Q�O���q�rk��E��[����O�]���sy)��������[o�m�����Ė5�v�䔁�=�aKK���Q��!�B!����bv��Xq7w8c���gܮ
c������ ��`� 7��7�B
���{��sX�z�}�~\�Љcǎl��-��f��¢%Kp��6m���Rp�Q��i������eŽ]�|�'�C�,���0]?4Y;*�u��818-�� H~@�{�S2U���ɪ�"w1\�_$��;C7�&�c�)�zB)[�qbݲ[�pq����_�o�'��!�|�[�����9��`�����m׬�Ӛ�զ�^?0�.ȩ�/>��y���a�����ށ��tRP��J�>\��Z�;zXz*W��d�?�d��"r��#�ꯌ6��9�k���]m���H~#�^z�%Kb��K4e6/q���:�%�ԓ����h�*���LRi��E���aFz
�� �B!�7�xtQ=�GG�`��wFc�L�#c���?�oZ�O�q�L,^���mg�i��y���{11:�=�w3�L
�sڸq�ԧ=ul�B
��3-8�J�C/��SOa��ٞ2���z:vŔ��a�����ڡ���F5���8v���|��d{{ ͪ0��.�~�	_0&f�%	��4�*u�F�ae+Y�̈́�S�L�>]z�����	���?�^x�%�a�
�ӵݮ>�{��$`��}����̮K��a�|�{�MMM��� !^D���֭����y��؇#'�&�Y{��(�\�o�x��yā�#?�#�ā]{�����<���X�~��	�|po�'��H)� Q��o�>�-���a�RI��I��h���e�!�B!�����Fy�%�X�s;���G�~���������߽�PW_B
�ή.i����ͷ�
�M{�bdd���ո���ر}Z:۱��QR������} �Ϝ9s��/9ku�L>�^�1���C�	ݓ5�r�0&ne6곘.���a~A�{�ڹ�������ك����$�Bw��2tc�qdH�dU6���O�w��Ο?�ߴ�9�?��>>�3-�����vD�^wm���[�y���Mo�l�,�Rm���¾ҙ���'M�Խ�FEY9N�l�ɓ'A��5k�4AiyN�mAk�^�X��Xy���J-��{�)�}�ۂ�B�ZO�A[K+H�#�h�$�	�l�Ǯ{{bJ$��F�����0�1���$UM�\t�0IE!�B)l���4�ʫu�1�3�<������oS��x����(-���&�CCضg�T/��ƍ�,+G��f\�� !^d���Xy�U�Ǟ��z�K+� �P#p�ڲM�	��G��\[[oWD�]�v��G@U+L]?��M�1S,�1��}��{{Ee%>��1�o��@�~��[�J�)��~_�''��&��a�
�'A����K�4Y���TF:B!n����?��?�?؄EKc�k-���
%��R��v�kW�����Ѷ̶ɰBQ+�f�oZ��-�^<*^��S�-R�왳���##ؽk]H�!��֯��s18<�ǏH7)Q�>�bi�Ϸ{�g�<b��e�v%�N��m7�����^:0x��|�+X�p!�ە��H����FCjTI�vy���:1�LP"�������<*��v�B!�R�L�����)^?������Oc, �q�v��͟��2�^�c�n��Z�x	n�󓈜p�������|F�q�o����8�u�wn-
C$BM�wahp$�Y�v�4�"�|��煡'h�Ӛ��S�b����b)F��/D ��F�A�{��7´�0v�KW�ʉ��rP� B�ɧۡ�MV�א���BHV-��g>#%�:�������o|�hll�ϳ�ڮZT��6E�&������oI�j3V����Qj,�rO�4U���O݅����̩Ӓ�;� �M�P]�\�Vzr���f��k�Dd�'��Vb�;�d�oˇ�H1�Qa疏�kz���~멧�r�y!��dc{�c:S8Iܮ��R�ۓ�[�a�:���%Q�<E�k��p���vB!�BHq��Ӈ�+@c�,�;��1��h?{�����V��BG�S��ڤiZU���:4�O���V�ٝ�|bѢEX�j�aߑC4o#EG���p�����˪Q�����^���d�ڞT;Tc�9�����n��7G�A�
������*�9(�$��~�b�A�4�A�/6䠺c��t�tD�2�:�|KV9���M$����
$����c|���QVVf۵]��]�M��p쿤�6E�N�����ܛl@:y�X�vZ����ON����zά���#���� <���>��M��u��cz�t���a��#:Ǉ3�Xqm7� K"rf�C}[>�G
�=[w`xh$�� /����c��̼L>�{{��<!.h����)�d���B(�<Ġ)E���?LRB!�B��+�!L�/��.�˥������_2�jjj��i�i"�XÞ�E�_���G:����D!1q���*i����h�8�ͻ���b�Jw�<�>��O���ow�������{�D�PF�h��aXs/��j�����z�B�.�����?ͺa>B�{s�/�����`�5�����!��SJ'M���&:�������7�x�t����~��t�w�׿��x��O&/4-�Ά�n��4�u[hh("�)J5���.�V�m��-�+���%iz�p�M���;48$��@H6�E�֭���p��N�=cm�7����c�"�/�k�<bS�o���z)T�:��� ���k�Ib�̈́����:��x�ڹ]/I��*���!ɪ��rl:�$!�B!��8�W��{�<0�.�F���`h�+c������?����m��s�Ayy9)6�;;�I��7�p=�**q�B'���9�(q�x�f�̚3#�c8t�(�'�AH�2>6�[�J�'$�Zqݟ�v����2�A�0�+��>y4h�+�,d79譈�" �P�^�Oգ>�-]�V~�4i�x�Jvb�L>�r�A��EONViV�dU����J
 Ye�3�=�6mڄ��Q��g��&,Z���~{t�a�N�VbÆ�����Z�����.C��~�ɭ�/�&����NMM����uY��r�ףzZ5�FF��>��L7t��^��ƙ��%Q�����2kǻ�Xk"rz�{1X1]�!l?q�(�wx饗��M�M�{&����b����KR���A'��.'�􅘺\\}!�B!��������+c,@NI%jl�f��q�F�w�}4��#�Ò���{>%��	)F��ư�i�����7�r�UT���'��؝d��.]�s�χ��ͭ�q���;�Cwo�D��<�裒9����ro�ͱ���o�����C�(�iͰ4��u��p����|��gWG ��Sc�3 Rz���!C1р/�qc�%%��	+�EiE��e�7Y��g�E�c�=���� ��w��-�̙��+�'-�&�4g%������m�R��wuL�jr���N����T��܅�p*����PYV.9��kj���I�~^��j�_��RN�jF�Ʉ�׹�^�"�:����t�<����h�;�2C��سmgQ~w��O}
w�q�#I�|pYH�n9A��t��5I�ԉ�p�~U�k�UVU�g�~A�[!�B!���zMcISd>����
7�>�@����r�E;x�6n !�N�+�$�7g.��.�����y'���؝XF�/[����I�X�ζb��= �$8��	=�.�x���z<��3�y^�f=�@�cEEs�C͈ϲ)VP6�ү4�vy�ى�VL��'�C�P:�
i�$j�k���C����pc�I�>��/)Y�JX��(�udP�.�UNF�ɪ?��O�x�"H�#~�?����7�BccC|�%���tm7۬\�������ܺ�X�����
�m�A����Ϝ��WVV��O��Or2���!2��m�5kP[W�`�s�l�؛gW�n�rʵ=�eC�  ��IDATl"�hvV\�m��<��I�����9c疭�����<��+��M()�U"�M�v��
a��>2]�Jf0jPzm��ALU��w��uB!�B��=<<����$S,=c,�h��1���W�sh����vyޒ%K��O��?�!�7h>z\�s/]���(]�.J�@��o��NT�����?v\:��8.[���,FYE9ZεQ�N�mgZ�z��wx��g1o�<�_e۽]y�'n�d��%c�`B�nb��f�������3������C����>�H6�Tn�"wݡ#�/�$��am�V��*A]]^|�E|�{���9�?����k�c�tm׏�Q�F��3��)�76k{�Y�Zm��a�R��Ǎ����S�k��0k&���g$q�`� �;&Ő�@\#,\��W�@�*������V��m����\�Qlѻ�[�͇�H1"����;���x�'�|�V�ʻ�T&�ɖ{{b�:Yeֹ]5Ġ҅!�A1%����"��FB!�B�a81V9%�jc�tu�lc�j���C����\��ψ��=���������ދ��1Ca�E���/^�w~�S@(���}ӦM���(HqSSS������u�>�9׊-���b̕���Ň?�Ċ+��SOeT�K��u�Qc,����P[;L��:�X��1c,��Z����%�-@�
܋��ȕ`�z>BWΩ�L#t���nꄕ։AvqW���ɪ\~�G�������&o��ى_��Wx�+_V��s)X�"t�G�]�����iQ��uc͋E-�+K\��b8���A��	ާ���{�/�������L��ۋV�Z���֢��.r���.@{�<yL�wξ`��1�k��Xܛ�u�o���H�p��atu\ �s�Ε\����5�v(��:�v�ACq{.*�{䚤n�|�k���B!�R�l>�e�c�k�4�Jz-���o��oA��8>���<� **+A����i\�-���k�P�󣵵g#S1��q�[�h.^���
L�p�T3���3���a�G[9���>W*������;��.�굆X�{D�ڡa-Pa�7�
�`V�.^WT�c�y���
܋�-�{��k}��bP3̠R �n��$$Mʄ�ϧqbP$������gD���^�VBtA���� r���;��[�����m����ܦ(|W��&�oI��qk�@�4	J��X�b��n�����/_�bD�+WbF����bht��OCkg�&:���E���?�u�iIpo2�h[0�dl��G�����8q���I��ӧ;�(��N;�ɚ{�2)�K��6NVYua�'�8:X�0B!�B����mQ�n��c�4bw��'̱lc����5G��z��v��	�FGF$�����#���LNN�����kq�,�7��q*��11>��ǎa`���BA���\�e���O��`?�> ][B�#��w}�U��p�w���]�˧z��y	�XZ#,����X�L��)��Xf���~���H�C�{�02F�����@ii��`��L�������3�E�Ps`)��%IN�a�d�ӟ1Z~�u��/��/�_�
�;��CcC#�\{M�B��D���y���T¾��q{NE�ľ9�m�n�z^ @[������r���jl�č��sg���҂��)���q�L,_�\ri���111��p�+*f���)TTVi>�}���:��z}���Z�����C/و-D�z��i�.o�O|>���u7�ү'����{����A�.r�J���k����B!�B����YS�?��K��X�:���$��{���2�L>c�������̋{����8�w?���FB�#��:�IP[S���\��i�G�J�X��� �`ƌX�b���H紡��<s
m�1� �����	�w�Aow�w#U����5�\��ݪ+&���Xr��ԵC���|ߙ��M���c��p@��-�cK;���C������t��M9�pc�]܃A��#����� '�r���g�NV�Y�׾�5lٲ��� ��?�9���k�7^t��E�n���: l7h@6D��m���m
X�ؤ^7���b_��p�#!x畹����U�#G�_S��u�--�����K�`��E��������L�'X�=��Ll�]�5�F�k��u*�ccر�#���1�}�po��XIy!���v�$U($�0Ӻ0�I��f^���H( �B!���D�b��]�˰f��a)̱����V(�˥vqW�3"z�Hc�������_�"�����;�4�Bm}V^}!�14<��C��kkj�d�Rlhh�F�LM�|�9�;w��y���Ι3K�.EeU�8�a`x'[[1<2BHv8y��ZZA��3�<#�`�f���:�նd�X��XH�������+��~����aY�bwӽ�P�^Dt�Q5o>ƮtYrP\�����J=�bP9��t/��;�3�5k�{�9������4eee�6m�B�%��ɢ��,>���w�ug䦭Jg��{^�x	�� �F��H�~�/]���oɒx1��]]FEe%�	Xu�f�M���˗q��XŬ�5��vll�CCL�-�w-��ݗ��|�8�n��� �`��=�h>~2�J�D�'q\�~Z�8���A��zD�]�s������0��!��Abߋv��@����n19��n_�����1}�tL��������t3���v��.��1��T���+ǻ�d�F�.r�oE�n�M��K��S��>�om3�����,�@���Orw*-+��Nd�os���������GǤb�@|���?�-n�O�8)��������[�xN\cY���K�#�<�6�Ny[�VL0�ޮ~V	ۣ��p!��
���$UM�t���vB!�BQ��˟�1V�>-�1VT�l��́1�a{�c}��4�����CuM5�-\ B�}���p�d�V(t�.��w}Rʣ�ĥ��R-lpp�Y���1�|̚3%����.vb߱C��i!� j���s���W���<7D�N_��gǽ]Y7L)L�%ʦXAS�v���B;���i	�^��"cwO�Er��/'�R��eG��|����&��uqϕ�SɬG}���=
'���q�����+���9���.M{����Gy�Z`$������5W���wm7�֡�!�Z��T�i�]�N��c�����I+�9�6��
���V�]���4�DOw7��\��Z�V:���(��X�����]m�R�F�G"�_[�����1P?��lX���Zi��l ��K�q��qId..n ���&�����ݾ���*��+�G������}�s�Wr��Z��~����xי'��kkPSW����$��X�Yc����H��`�KǠz��T@����`����+�3}�F@�̊���M����F8�Ϟ?ב�&c��nth�sg�&��1k���>�{��Bߕ���/�;���DaA\c��8����ˆH�h&I�n�ׄ�2V������\�ɨPP9Ԡ~�*>_����` 13�X!�B!DI�H��K�Rc	w�ce�|�����/������4�8�-�wy%��v�m1i�s�p�� �PQY�6Vĵ�n���Y������S&9n}w��?�c����������TK�!��E�cU��,zr�ꄢ�%ȔN�b�h!�w˨e` r̷���m�ω�o&�/j�������_�W���n�ik�h�`�
C�Ҷ��Ν��߽y@4	3@7(��V<�������~w���3��[�}�%�n����[�Ш8Q�sω=7��z�B��]i���KU/L̯l��+g(n�
��AܺbF�.K���T�ܣb�`d�:2(;���KVes�����ꫯJ��'y�o����������+�����'��O@���N�f���"rk�o�?:<X�8+�L��+�{EE%*++��f�j^�S4��k�v���(�&3��+ȸMz����{yE�鄁�}�m��ݕ��'r�����G��6��:=rðj��(���W�Z����@�#�@� zzz�iddN!@e�_r�����pK��{����>�E���A��1�\���]����>k�D����uY;��ņ��w�l_�=:�a��5۷� ���K�.-�l�,e\t�v��dD��lr8��vA ��t�	�cI��>�w?:�;l���k,�z߭�y})�ͳg�v5�de�v>cڽ=6���$��*Ɂ!:iE��$��������vWL!�B!z����1V V7LU?�c	a{�����(F�{��wq��������<y*���+��/r��K)��-�N��>��&'DoKW������^�u�m�������{�H�Nolpe�Ű�+*���5�7{�T/��9v��%��E��!n_�t)�@�ubT��.SUU%�g͞���ӥ���y2�y�"�"�R_YU���d���f~B0�c��ݏK�p���qe�mE�ߊ�]���l��w�b���d�)�Z��k,�n�n}�[n���w����|5�J���ͱd���$Kq���$+j���1Ɗ�����`�>X�8X;�
�!G�����!���?���p�Q��r�HJ��r`�M7݄�~���oA���#G���������z�E���X'�Vb�������� *5n�Ia�c�{�";�s�վ�7u�Ŀ}���|�t�;�Pŉ���͑\�++*�s��	G��ztt��C����G� ��B�E�_r���	Q��|�+���ҿ�����$�q�t3��i6x�������]e�x7����oؤ��n���y�jl��z�N�8	�=6l؀/|��8+�[�[�:Ie��Ҿ�s`�wb��C��z�Ae�J*T�-A0L�vB!�B���@7/�����1V��$9���1�$nE33�ʤ�X5�z�W�)�l�,�##���|�{]sR̈z^��sҤdxh K�.�5�VH�A	)�	����w�=�������n!j�bD1�W���ɓ��7�O�c����Ckg��������f[�v���}�פ��e�ŝ��:���/IȮ���'O�eqa{L�n��5{�BL������{+/���"�dw �.�����dG�ȁ,:Y1iQG�����&�|YMV	��^�Un��|7q�۹s'._��->ڴӧ��M��lQ�h2�����+J�C�����[��Tp�Dl�ž�D��/�b��e�J)�5��
3������ʊJ���J�!�B�'}V��"���yrrb�X��A�?��>��3:6*=�,����P^8��ϕ��I���p]�c%�)v���X&M������@/�.v(D���a|b"i߄��kD���Έ������;�~��|<�3]�8��	�{������R��g3I���Ʉ��%����u�$����=��r���$F��t�I*B!�BIő�,	^�7�ҩJSd�/�c�����X�e�&�oN����!�7Z~�7JN����A�E_��ݱ��y!��0�j��@o_�2���^?���쪕(�N)�F�����X�(FF�1<4�9*�ΝB� ����	VuM�+�dX�_q�E�+D��}�҃��˸�y�4!$�׃��n�@_?��xꩧ�v�ڜ��-�n=0�g�?�V$�+m�Pg�gف]6Ē��)D��I1�`u�%<z	
܋�։�莊�S82h��"	��dU\�HV�fC)�2���7�l�s�̙x饗�_������_Gn&k��ڵ����I���R�l>֒`��\G���`s�Y���W9�g�:6Wb_��2g���H=*T�S�Z;�E��P�1S���`�[k��m�d����k�q�̮Լ��j�N
���H1#�\��n�����x��'�~�zǓT�*t�&���q�*[����uA3Ġ��_��K�w!�B!$�k��F�$cɓ�'��V����"�U=(�������،�v�؁�/�x����8R} �n����F��z��JS*D-D��b��Ƃ�3���e�ҹQ�ʅ)���d�%�#1���wq�'����K|UU��'&Y�xr*�y����Fϗ�u�q��(zGq��Kzo�w%��?��CW��x�b<��s�y�VC���V�ە�X!�)�~�Pֹ*G|���5���V�۽�E���)<��cÃI����{�{�Mwe��D�yA��Rw����7�)^7�͛7c��� ��?�9^��KX�d��ޒX7G�vg������x\+���%v�&"�����V�j���k��U������w�&X7[د9�ۋ�W�v[��l�uC��<R�g1L�f�x��z���U�vNp­��gI'a�����J��Jvo73̠<�`ii��� E�N!�B!$F�T=�Q��9V:S�`��/sw�c\�1Ɗ.J��9e���.�3f���/��������h>v�Ӫ�j�� �x�Oˮ�@���^�ԅ���B�8q�(Z�O�xq���o|uuu�����=.`���R�ci����J����X��@�ܣ��)��i�������i4�1p���INFn�v]�u�U@R�J�ٕx>��r��_�u�߿ccc �B�����_ŬY��L�Js)V6�S��6g=ָ�&��C��
X͋}aK�k�]�q��H�wq@�������e�x�V~W�`Wnk�7�k{rX~�G����	l۴�c� �C\����zWD����J$���̹��vaH��-���3�k\����@!�B!f�{Ac5`lx(!P�b)���^�1��ϸe����cӦMضm��8�t UUӰp�bB!�hi?ۆc�x�x w�}���Vn�e���bv�~/3�v�1��k��KY3���f����{
܋��<�d����+�U�F< �۳�������U������իW��_�2����{����G���x��WQ[[�i��͑�=lO�l_�k뀸=�"r���V�����>����M��h����T�:�ry���3��W�v��k;���?�ÃC ����ý�ޛ�$��I,{�ǧ�=�F��MN�IV��T:�Z��f�A���� �B!�b�󁙘���͚bY1�*)�E�U�Cc�_.��p��X��� �B��lہ��
̞;�B!2��.b��] �D�����+����!�S��S,e��h��t��F5De�P�ό� �۽	�E���*�5���]$O����:�g��R���v��L���~�����q��i���ׇ�|��x��PQQ����\ۓ�s)V6��-"7������������žV�e.ΚX8sa��X�������a��ߕ��6����V~�6����aa���k���#���Jw�7����kI�܈�3qoONRe$l��Q�$U
a�ֽ=���oX��n��B!�B��H.�Qc,�!V@�⮬�5�*)��W
�i�em�ʕ+���O�����A�����ܲ��̽��>�B!}����6�:�x��^z	�-r�F�d1�g�k�Ɏ����F~N�O�ޞ�n(���x���v�B�{��LVŇ����]ϑ�L�J�R%�����&��I����
N��h���Ւ#�[o�%�{�=:;.�g?�1�~���;#l��،u@��h��ľ��Y���m��0ڼ��l�V���	������^lA��[i�����ۍٷs:�;@��8����X�x1���J�<���0�k�U�Ĕ�}P��
��������~l�aF!�B!�lD}�+�)�9�d�{t~v��
]خ\�����1�ɓ'A����$�o��~�~TVU�B!����0�m�,]o�a�<��cyU#tG螬�1W+�^KN��XA���ں���L6���ޅw�JV�\܅�ƍ���=�^���&�R$�"�O��dUt�ۉ''�if�m�݆�~������MZϴ��?�',[���\۝���X-lߴ�7��{{�v��ۮ�F����&���kr�s"r'��v�wk��Q6��Vb�濫�!r�_�gl1rd��E��wY�v-���/�U*�I�D
�Iߍ��{�*e0Ġi�����fD!�B!���#�G���Ȑ�+��{�ߘ)V�+��9Z7L���XJ�,�C�	����䋉U&�4����*����9�>����>������B!�����}�c�c ޤ��o��&�������۔8m\�Y���a8�di�g�1V(�� ��
�I,Y5�#��.��d*Y�%����LV9��ufs�x-�U�w�Fww7�79y�8�&&q�'oW] �V�l>֎(�86�bes��D��������m��:m����(6����m�B��F�����Z��-�.,	��g��[���z!	N>��c'@��HN���ۨ����s:I�ny���$�R�0�JR�b�ȅA<����/�Z�	!�B!$S.c�ܗ�5�`�y���9Vd��+1�s�1��}�b~��4�~趉�NlS+��y���7��&��ضi�._B!�±}�bhpĻ<�����,�����ν=q��5���5ŊNA�Xto/\(p'�3Q��MV�M%�"��KViUJQ�V�+pqRˌ��9ud�d��ٳ��o���.�w�|�������?�c���X���D�v�f�i��L�+��ޮ�c�~W����uLD��_s��n�3�tm��`�����4�Ʊ��A�ͳ�>�����4I�F+�:�T�\�U&.V�TF.��K0�Mq;!�B!��a�cc,��{�f�_���{��`d�'��5C;�X����5�c��{����ě\��EYi��Z9^� �BH�#��?��W�@��ҥK��/���F�fQ��W�g�eT;jꅉ���a-��
܉D��*����bSP�̴�*�2Q�x��,�>�Kɪt��A�ne�C=��۷�����.���@MM-��.S�/:#`ͥX�^�~[-�+�����V�����LG~+�`�X������n��vm����$X7g�].?�b%��vs��m��=M �檫��W��U�$��I�l���[���J�����	�S	ܭ$��\��~|�B!�B!Y�+<��X��XA��(F{���BP��McA�WU椊�kƌ��7��w�yĻ���`���q�]wH�!�B
q���m�|Ļ�7��M��չ^t���&��R��bI�B�u0>�s|h���3"�
�x
�Ie����]�*7!|ɪHg�����i:��{�D�^�J���U���Ӊ#���t������Ž��	��� ����ǴiU���cr)^tB�k�]��{��&l6�}�ޜ
���/J5�]mÍb�z¬�݁�꜈܊�^g�#�{`WD�����4-�7�<]ۉ�K�]ػ}����;o��v�m���&��-7^g"A�c"A���R��HRI��{Ҁ�{�H7�7B!�B�;ڧLc��
c���Q����'p�d����K���{�̱���?�x����۱7�~K�\!�B����۳m.^��6�>�(�㎼��Z螸oӘc)�!��hv�g��=�R
��5�3��y��
�Im�J���6Q%'��	�H����d����OV%92@-p����J2���ϟ�W_}����@�Ϳ��_QVV��6nHZ朰9sq�mn�v�[�q��[��Tp�Dl.žf�d�N��ڦ8��wuFDn�����|Ws�����r�8ЏP�m��]�c���u.�6O?�4n��Fx)	��$�n�*�dօANRE]�e���I��PZ�Öv��!�B!�;t�g�.�1��n�o�ҭz��n�1�ۗ����ۇ�/�x�s�gQQY��7n!�B
������<��Y�p!^z�%ռ��«�_�O�ꆖj�s���=1i�i��ۂ��{{a@�;Q������:�{�2Y�OVE�4��Һ1@�Z�O�OV�M,�˂��Gy[�nŖ-[@�Ϳ��/Q�+���I�s)lvB�k�]Fq�Xu��ir_Ym���vY��|�iC�����pm�ݼM���X��p��|�� �"r�ǻ�8� G�Wa��}���:��;��=ر�c�:�x�U�V�^P�s:�dkv�sI��bBJ9A�LV��T3��UtJ���qo��%�B!��Mv�O�E��a��{�W3�����;i��+�l�o���x�����~�9<�s��I�����ցB!���}�z�������ַ��А�5�t˳UCL���̛b����X�b��a����D��� ����Ã�d�*Qe 4�&�CJ����U�ӑ�L��� �K$'�F�*%�$\7��L����W�C���������%%��\���gl����R�l/V�����\>�`�fŵ]3ۑ�J4X�Uf��ι�g.87�Wf�oi[0 ��y'\ۭ�Zܛ�3ږ�8������I���1jڏ�o���x�W\o����4I�+g{I��ܓE�	�3�*���b*+�cS;!�B!�8���#��qwq_��c�
����h�Pi�U��7�
��c�Q��*� \�E}�h��>(c��O�6����k�_B!�x����Ա �G���y�y[#�E�j�PO�.&=S��#{�����t�b:;E��B�w�ĩ��\��ڵBw=�A���/����dUII����ua���P	ܕI��]۩�p=��F��-�׿�u�����@������?Ǔ�|�פ����t��D���;�M�5�"rb_�X��]q=���?�"�,�9���J��n�9q���ݠ�s�A��{�M9"Bw*� �W��~�SSS �����-����$��$���'N*�ۍ�T"9��T	*Iܮ^0_@�aF��N!�B!��4�R9�+G�N���A?|¡=�F~����X%P>�4�����(���Wu1a{���HUK|��7%c�K�.�x�cK�?_}�ZB!Ļt_��s�gA�ς��+��լ��ܮګ!����(5���Za{jS,1�s(a�%Mi�Iu� �f������$up�����R%�dwI�KT��jGw���&��bw��aMG*w��y�L,��f��_���Ȱm�6o#��_���x�٧q�իuc�
s&��Ю�X�f��ka_e��ᤰ\�R�׬���j��:m��m
֭��M���C#������k{�D���\�S�n���~|��QV�۫B`ٲex饗T�
=I��<!\�bJ/nO���VJ9I%����k�������gB!�B��D��zMc�uÄ9��K9�s�K[/�k��$���6ƚ7o�d�����f~� n���Zk~�gB!����N���e�#��_�u̚5��̰�����L�Rdc��4#>��
c�c#3"��!]!A���`�/G��D�2Y%��+�Vqa{ܑAt8%�$UB�LV�"�'�d�{�d�]a����pQ��\�Z�-�y��8q��� �F��ӟ�+�=��+V����;&`�)��6�u������V��K��������oC��9�v�+p"���*�ǻ����o���$C����������� ������QWWWTI*�r�	*��[rp���bw�[{��������1YN!�B!�9�1֪es06xEe���i��^����!���	��XJS,�1��^�c�|�+���L�6m��}�; _��Zy�U �B�w8}�$�D����� �������_�fX֖�SlN�{:S�ĨωZa(6iGz6����6���V��*0�.�zX�b.F��S:2(��j7B�`<i%:�D�x-��:2��hE1R���9%����ƺ�b.\��^{����(J+ ĉ�g?�q\�n[D�+��v9&`5�}K^'�������)��+�ς�ּX�¶��n@��k8���`�ǻ�:���-���m����h�ُ�5Df����� ��3�<�[n��I*��4WG�n�y!�����`�A�}մj|p��vB!�B����,p9�K3��n菊��џ�I%nO�9I�Y�V�n��i�,�j������-;v/^�>�4I�,[��B�Μhơ�� �����曖�J���Ś]nv��{0�Y��!idg���Jc,i��K%rW�cB���5��@

܉!�z����r�SP:2�ĕ,f�
��Mv0�uc�%%���:�*ّA+p�]4�*iN�U��`%q��#����	��A��,r�`�U�����-�mp-ę+��t�Y�w�x�岀�8.�b_+�2km_; ���k��v9�]ͭ���n�̩k��88�������ׇ�� ���5k�}M5/���F��Zn���6Ġ�켠�'�0��I�v����{������@!�B!�@�K;��v�g�1���}��?� ˧�WL���W/E&�|��!
���Fbw�c�
����*�r�عs�⭷�¿�w��0طs�t\�XM'wB!$�ii>��{���G<<:s�̼���V���Q�c���P
���c��1�^�P;�s�h9Cq{!B�;1��?��W��ؕ.]G�N$���qd��yr�*1�`A+t7���Q�N5_���l���7��<x��� �G�|����K_yk��F7�PD�+�ѧD����E���C�{���W�u��p�v��3�[�+V6�x.E��(�7g�K�s�u���n��X'z1ؼ�u5}�W���͘���`����_��_cڴi�'����̓X�$�4�t�Jx�T.�@za�2IUS[���'at?H!�B!$�$cE�ϔ�C��=n��u����c��d�1��պ��>�ܹ���oA
����cb՚�A!������q��px�'p�]w���Jl��'��4�X�eP����c�ҍ��c�%�p8���@��w��m+pCyX��
7m'"'���x�*�Ŝ�J�z�DבA%r�Z�''��dU>&���,X��={6���oKO���G���;��g���O>���U-���R�k!Ζ��b�Y�w�x�eUpos��ͥ��l�>n{_g_�O�v��լ�����>�um��_e�d,Q��݃m�6cj��х��/��k���I*�$���~�Am�*�HN�sa�'��΅fE��c�B!�Br��+3Ē'�{:�n(��*S,�B�����tE�P������r~!���Ki�u��9�������I��ukA!�������c���R�PI.�~n���k녲9��ڡ�^�1�
&j�1c��|�)&z�&y~��E�<Mq{�B�;Iɥ� *V-�xO{\Ԯus׊ەw��Ȑpc�&��Wrr*���:����qd��i�l:6�����;��c�ᗿ�%Ha ���L}�Ql�x�����be�dEDn���^�������|��}mM�6g�ޜ>4����޶ۇе�|�ۂu
���s�2�o�SS�7�t�|�ɬ$����R#'����ҭ]��JNV�D�DSHG؞�ĠMRń�u�x�,�AB!�Bq�1V��K�n��
��_g�gq��5�J�F�!�S}��^W]C�Wa���Ϙ1���|�M��A
�c!9��n!��>��&R8���I����Ei��~��f�6�
��^����>�cik�w��β��� �	�$-�;JqG�/1�b�Ay�A����/��Tn�!�*��]ב�DUX���I��7�M��qdx�Wp���>}�p��_���w"w%9�Z�sB�nMDn �5)nwFp���v�ľf�d�q�b�����n����k>`�_0����k;1I�������X,$�O���|�;(//�]^Lnj�:Ae͉!�vl�b0*r���%��)�o���wB!�Bq#c,��]�n�0�
J#?�����F�P��k��O˳{뭷⩧��O~���A���q�n�B!�=ăg'�),��ylܸ�hͰ�u�dQ{�z�~�P�gu��ص]�*k���a e���}���B�w���� J,B���:I��jWԍAv0(�3�UQg����]�l��G֯MT�'�	�BsY�[__�o}�[x�7�.Z`��������ƛo��;#`ͥX�\�Q�Y���j=/`5�]��S$���Zi�~��6~���bs�Ј�{{�tm7�`��v�tu\����I׺���u/[�,��'+�NmK;�t�
�e��^�*�����$�ERJ���k�K�vB!�Bq�$c,�)�_�K��Q�ea���]k�%���
c,m�P�0(c�+��n��Ċ�/���d�u��Q�¡��q��s���@!���spOΜ<RXlذ�>�����/��-+��"we�PY/L�9$��
��k���:bd~ii)6��"�
�.�S|p��5T�9�+n�:2$����z��%�����h+w����\����zo��&��_�%�������o�ѱ1|�t�: ��爀�R,xs&�7�|���Ή}Ͷ������y��.m͆�=��u��+�����ݬ����Vb��o�>�϶�i�.隔��?>�����a!�I�t�R��k�JP�qbH��S1��ƠLRE&��4PiGQ �B!�7Ic�%��1�{@��T7�w�)�v�gu�Pk����'r`�#@;e���u9e�%�����o�����)N=���Il��ƴ�"B!�dq��o���i),jkk�Q����t�Z�0�1�y��u�䑟�\�U��ͱ�
a�4?0�����f�С���bl*��i�Q��j8�V�.�W��ew�h�Jv0��'%��ve�
��]�ɪ\
���v2�������СCػw/Ha��O`|l�>p�o-�D�+�ͥXY'>+"r��\��Nۣ�z�vžV�e>�����~�Nã��'���9�v�v�}��v��S�n�ph�>��dѢEҨG�>E�n�\�q�Jߵ=�HR�9190(RF�ve�JρA̯��g�P�N!�B!�����x�1a��4Ŋ����XZS,�޸n�4�sd����+��v������/����RX�4����>q�-�<!�B���.ݳu:Ν)<^�u�^�:oͰ��fo[	х�V����k��uG}����+놱��beU~�RP�NL�Q[��c�#�"w�$����/;�xMR9h(r��EJ^A+�R�28�Ȑ/ɨtɳ��r������y����;�n���y��O���-��gE�j�bs�4l�M��6��V�����8�؜>aAp����ᰅ��S���u��������o��\�aA\O�������.a֬Y'��rc�e��ȁ�8A��� '�B�2��/�HT���-��!	!�B!$? CUQ��b�+�+����퉺a��ݠf�CΡ�1��"y�mx��gq��alݺ��h?ۆ��n����#�BH�ײ;�lť�.��C���裏:V4�L���rum��K�~�5��3ƒ��Q��ͱ�������%�
������&�Z�0+0 i�4Ԡ$lW$��L�����rP��Ҿ�R1���{ul�����B��n��Δ����WU�������S�o���\پ�nuuuV�u�L~���5׮M�ʐ��t^�DӮݖ4�ר]`��+���뽒r�[��Z�|t��ȍƁ�}iV`e�fE�����FG1<4�.f�"l�t�PX����a�m����i�im���4:2*��=�=o����	���<r��:��M4�Jd��GO�ޘ����H��^�S�2+}~�n�/E�r�Tl��N�Z��u���`�+�b����z��0>:�����vڝa��M���D������]����9��k�l^gX��k,+�^to�����э�n�J߭�ع]��ҋܵ����%�롸�B!�B������z�������Jc��џCIuô�Xr]L!vO��X�XW����"g����hmmEW�Z�%�=�@n�[ۗn��gc�Bl��͸���#ksy��t��S汝��m��}ї��}�������&���}����u���nQ��;����oK���?55��[������y��k,e���k,+�~�x���9k�z����5C$��qm7�9�9V0f���W�����Sp�Br���������MRi�Ը2�_!|(jP)r7rP�����EC4f�+C��*+�n�,XIb=��طo��_�E����/���}Y�499�����>��]�����?��+*5K�_B�~��7�^�i'n�߲r�'�`�B]�ё����x��v���7���k��� z{z�l���Z`��TN�G������P��l���S�V��}���`�X�OXqm�zq��3on��n�l�Ѿ:q�(��vmR��m�h[��B�~��5�Ӟ��ŎNT�֠���DK��6���i��/�z����+þajr
]X�|���M[��]��9g������/]�m���J̞?� ��};v�|۹����5V��3� ���<��5���w���%���S��1�KR�3�q_HNVA����MV�0TTV��y(�B!�BH��%8=5������]���9��9�P��n(f)k~��X���&��9���K���s�J��~��q�����UUUp�Wrk�⻋I�?r��l}����ܼ˯Ziz
�{�q뻋<nW���P��k��藄I����]��pd��cc��OF�\��B�.�P�P���y���Hn��&&091��b>���vdx�"FI9{����-��ݾ�rs�b����)�73�7���=˿���3g�̉x=_j�Fˣ�Sl�A�P[7T��
�{0.n���H�4�slY����v��^,P�N,��W����h�#r�&��	�`l����];�`ԕAߍA�����G;^�s��s�@�溲!���|�M477��ѣ ��pr��?� O=�4jjd!�� �쵣ia{4�\���2k��7)̵)`�&��<.ulvž��F��]������n,�"�p�^���� ��+�;�Ě�m�A���m�9�sK�7Ļ?ކ��N�¤����***t��C���Z�`$hW��]�b�����T���0IE!�B!�ȡ�SX�|Ƅ1���]�k���~1O������亡Rخ�
i�Os/%yh#c,%�P��.�m�뮻��#��?���3n�&���_YY���)���NcMNM��ލiiFz���h�.\ 7���K�-��~�i���]�~1��˝QSW�i5��w�L�/a�Ⅾl_ț�.��;257���Z<P4k�W�`�q;<4���lK _��X�K�󸅙���+�ছn�k�s5B��DM��+]�PL����>k����55CQG�m���-��˜���U1�ۙHRiD�r�J��roW���C&;2$�1�ܣ�&�2h�UN%��-�E���jjj��|/��2FG�y�8���.|���{<��3�5{V�r�BIkbes��D�������Vž%ڇt���V���m2��"xgD��*��kǵ�(�����dlV���~�@a�;ǖ�~���+ ���&��e˖e%�TxI*��	q{����=�Z��J����B!��Q�^��5%=�{=IخqqOvr�Gk�:"�Ľ��nhd�%>�}X[�g�%)o�sQ�溲e�%�<'O�DSSH�!�r?��p�=wazC!�b�+=�R�pb|�0���[�r�g+��Z�\/���OV��ʚ���];�sP��rr�N��zv�L��͝�S�;P�N2bsG��E�Qr�J�ZύA9�V�.'���jG=7��]�.|Њ�ԮF�^wY����k���^�����0������ɧ���K�H�r+V�k�V�bߜ
�3�K��7�6.u���������pm7/X7�!��|g�0�������i������N2B�/l�`��/)\�x�	�{�YO6���l���H��3IR�LP����TCtU�` '�9� !�B!��;����a��˧c��4��5Ŋ������Fu�0QKT����ʆY����+z�\��X���*|��ߖ�����A
a���p˝w`�� �B�y�:.`���%CR��Q��~���9�fX�c��v(���^�P�KYC��S�c鹷����q���b�w�}c�Nh�B���K$��!	+��]��Ҋܕ�Ɏ�"w��+������1q����&����СCؾ};Ha21>�������_�UW�6�9���,��͋E-�}=/`5/Vv��<�Bd��F�Έȭ	�Э�߆�ݡ�Ftc-	��f�os�o���=z�{�c�G���.�AO�LfՁ�knV�T�T"A�.I�/xOva���Ӹ.���uU���p�CB!�B�'�X�����u:"wm�P�'L�*��N�rmP9����]4FQ7L�?�Xn	۵�W�Z�7�x����@
��T ;6��o���ZB!����L+���#]k��D�S��=���Vb�yz�v�	�z���=Q3L����Z0�Ҋ���~ljRg���$c�|.��ά�7�qq�KX%�%��q��,nOvd�{-�,����NTIsJ�;2�C���甯���s����R����?�'����q����/V�k��6)��"�Չ7ܺbSU����}�����.&�Ypm7�k"�|�� ��+�����Z����ݢ������B�SWW�����AmmmVSVב�X+m��3����+�Uz��PH� O!}Q{�vщnﮎ���B!�B��d��`½g�5Ø)����]��=^/L���X%I�v�~5��a>ce;�����/H�X�6m)L��o�n�����ցB!�?tD�Ha#�a�ﾜ��|.����Ê)6GY+Lc���#&�#?�������u�)�f,��e�ۋ
�I�L����?�HRe��.%���VF"w�9�SB�r��$�WFu�%���Ƞ]�f�w��믿���1��������Q�uϧ�cS�}���Xk"rb�|�ڊ͡��t���Z��I�$V6k,�\pn��r&��k�w��������e�:�7P��.gN6����ܷ���׽�W��zb*�r��JvbP:�+]B��v#���{{E�"t����B!�B�ğφ�9�059���c)E����h�P�9�1�@�.������9�����&���p��a��E��FGF��OH�!�B�k���p�������ǫ��j��M-�Ͱ���A�9V���ܕ5�T��t�XA��]���V�k���X����b˹ ����Ã��+V%�����=��23�`8��F_G;�h�N^e#�n���(3�'l1����������6t_����(*�˥yFb>G��a��w3�̱��^���J�v��	��	�ai[�b-}W�������[�׹��3��G��C{����S �ϓO>��~��y��2�l�!�I*�����Cl*++æv?8� !�B!�x��`���P5r���ݴ1VL�.�eq�c�D�Mm����Lb�~�h{b���|�;x�W088R���i���(n��(+/!�B"װSS���v\��	R�̜9S����:�uA��p+V;O]3��6�֥]׹=ͨ�qQ�A�P�=K��X��������^�t*�����\��{ّ!��J$�tE�vHI*��=�z�A�d��$�2��x-�\9}�4~�߀6�O6�'��<���t�[+���&"� ������w�/�5�&�u���Ní������[����r�x���,<a�m����{����w���� R�lܸ���ZV���в�^��&���ۃ
q�����
�������1t9B!�B!����|i�L�����6���}�Q��N�F"�T�X��f9�m�+۱�4�J��5k���������2/Y�\�Ѕ-����.�}~B!����0v|��|ȯ��b��e˖e���K3,+����R-��#��L�5ĠB�n\?L��{]�8�R�^�P�Nls�7��V.�ؕ.��=#w)a��ۃ
'�dq�*a%�MZ�eRՉ�آ8��`�Y��累�z�-���p��"�bg��������U��X-��M��mǰ]y+`5�]�tmOw��5�Z�}mW�l.�9y>
�a���U��w�߅��p�\ۣ��
�YD�>#�����G� )|�����i�\ML�C�l%��\���r�jjJ5��n:�?'�T�Y!�B!����f`U�7zߧuq5B!x7��^�pq��C��aJ�;27��D�^�X=��?�_�� ��@_?6��'�x�- �B���������s�<����h�{���Ųe�5n��n'��۱c�]����q'�7{��&q��-�Mb'��E��"�V�3��f4]���$H |A���_?��_�8$p�������E[k+H���_�:.��Ҵ��n�ͱɞ������fuC�`,���v�>��m���u�4�g34�Wx�X�/͕�U�Rܵ���Ƞ�T�X��Q��-��`p�V8�PY��;c��Rm�o߾X�r��v����w��Ԅ훷b��Q�>sf‴��m�}�2�[��X��,>V6ҩ�W~LV_B����#s�C���+2�po�`�}��������{ة9��^쌥���@����U6 �=V�Z�4���	SV�K���"���=E�����,�=�\;��t��B!�Bz.�;0w���W�}ƚa��^h������#���ڡi0�keU�ĤC���lƺ��;QQQ�6��nZ�[��;�0m�t�3�BH6q��!l\�!:C�&��w�y�ַ��[���`�a����OP���bi���������G��8PFs{�C�;q�ږN������D�J#H%�&�q��,�A��h�*%�A|�
�{�w8!�!6���Q2��7}�t�X��>�(�uY��{y���ŗ_��˗şH��ܢ6��{9�M������u�Z���������mwbnw�p�}ú;�y�������/,�Mv�Fs�&t����8�M��|�������&.���#Luw=�"U���^2�R�TS{<�!Uz{�wc���!c����vB!�B��~$�S��Tc{P��97e���f��S����y�u%��4����R��ѓj����x衇p뭷����w#L}��+wx�5o!��l`���ʃd�F�>���BW����o��V��J�JR7�q���Nmb{����F�{A���k�s���B�܉k�q�7�돖3g�b��ԟ������}�V����U�
�J��"�����.#�����g�g�������Z�:N?����


���Dn� �7}�t�}���6����]1�K�:1��l6�x_0����1��ذ�����o�I�X۽A�^wlފ�;v�d˗/WZ:����nû��P����<���Š��=77o+�:NތB!�B!��ƶN4�����xr���.��Zab�0�3���@ch3�{��`,�8k�XZ��	vw=��9a�<���(�TӬ@���46b��s��SB!�7�b���ء# �A~~>V�^��cǦ% ��6����x]PolO�e�On������n�ţ�t<�ڙ�Nhp'.�� ��:�C��D����hnO�ȠMqק1$3�KD��ஊVF�JY�"��e��]c�v��;�@YY6n���ޱ�+�p�>��*˜���ߣ6̾v����nS����gSj{d�3c�7&�L4���&r�72Xg�8�R��p��:�����B剓 ��ȑ#�r�J%�A�Fw'��c�w"����Bz{G���`B'����vB!�B�M�q�7��֦F]�P<�њa���њa(��J���܍uC�`,q���3��Z��'B~��_�d�fC]=λ����B!�7!n�����P_[�=�~��X�ti���UO�_&���2b��j����ϝ��B;�v�(�? ?$�>'�!���U������#�\{���nLb��U�D��`��McP�`%�	k�*�e63m�Ay"C&�QN��2����~����ѣGA����J<��_��[nI�86��0�z`����n>6�f_��d�M�fa������Æq�o.�lX�3��k55�{pӈt�N��n��K�/���g�$�hll��-�PWG�*�())Q������0ee=#����w�z��L�
�E�N�@��Tک�QR�9 �(RB!=����Ĥ��<�~Mc3�����e!��<�� ����Pm�����Is7�ۭ���]��)�f&�ȱ$�Rki�e~�e�QK��o��ػw/�{�=�젮�o��*ιp9��B!�7P_[���>A[kH�p��_���Z��uA���f�6�*�e��l%K��cu&7�'3�wv�����1��D�����;'���(�w1�Z��)w��n�b����Λ%2�1���99�Q�Fa͚5��������4�����w��EX~��'���XG�v��v_�|�S����6���ڃ����v;c�,�_��~�aYr���s\q;�q��&t��{=x�?ژR4 ���}�=�`��i�������*.T�E�pT��=$-�*�Z�23��$���0�� �BH�c՗.�]7/�|?�'���_�B�;!��@v�`�)��RsR�wY���n���)����F(3����w�6�ҭ�QMЭP+7B������#�(ɗ�4���ڰ���0k�\L�}!���̉��Q�g���F���3g��{�E^���������_���z!j�F��ՎϑyC0���Vh���â�c����v�w�:UM!�G�C���������X7����V�J0���ј���^�R���Cvƺ����c�/V��x�	���7�F]m-���ӊpiĺQԹ)U���{/��1�¡���1�lӱYءa=#L�����3�1��X�n�ph���װNc�w�����۰g�N�|S�Fz/_�җp�7����%�)N�����T:3�{"����G��r��	!���H���o\u�r���/��N!=�7�by�x����n��9�f��uj���,��=!K\�F�A��}�Xɶ7d�<��c����ǎ�Y������4��c��%��+!�ғ��:���Í8~�(Hv1x�`<��8p���@7�v���}�5���p,�P,m0V(V?L�eZ7��H0�����c]G!*4�OX{�׎*E[KK��`�`pO��I�*c���@%��2t-�Q?��I>�����2]�rc��믿^i;��?�$�ؾy+N?�>w����g�a��!�ސ�.=V�0�ߵ3ú�q^��~_a��6���������a����F��{��=1�3�=3��{_��"�����q�m��fn�4a��zFTS{�'$�T&�,���He�����ݿ(RB!=��?a���*_��b�����yI�y	!���Z;=�>�7�Gk��g��Ě���,�][3��@��H�0��n��il�n�k3�ټH�|���z��X]�d�*�Lc#ν�|��B�	4�i�o����Z�d"�}ժU�:uj�jz^m�ͱ��`�?#�2�	�?˂�B��ϝ���p�Q?4u�Lo'zhp'����cx���C(� Ms��U�D�@@op��4���(X���+�����l���]w݅cǎa��� �E�J<��_��ǔi��w�d��4�:4�:4����q���N��f���Dnq�w���o�ll:Sϥ۴�[g�/�����mX���[j�k��;�)B�>&L���+W����u�(S�����#R��ۥ"U�4��؞�ܮ�0x"��in'�Bz��~��/�e�_�|!�]�&�+��	!���ZE׍ꋶ�f��ݐ䮭ƌ��Rj��`(ftWk���������;@�c����ow=/��b��+�@YY�}�Y�좺�4^�e�s�29�BH&s��1l\����A�q�*B�.��b��~l�;ce����aX�B����`�`��,�=e��~����Dhp'���D7M����q��!�A+V��Uc{ "TE�E�$m�{��nfrW�*%�A+Z)�*eI��D��y!@Y5ډ����x��q����� �E[k����������/�T�{X5|���z������qfc��ߵ������{a��s\޼V���x���3�xKž2lٰ��QYJII	y��92m�t��)��H��,}!��S�J�0Oo�U��E*C���~���
!R%��B!$�)꫾t����+#/�I������1c��Xfwy�� rB9�za V3��U�j0VHW'hk����X�]��ڟ��X���wp��!���� م����[�9w��H�qB!�F���޶Cy����\~�����Z�ϫ ,��pg���]b�2��)�j=��eLm��
M����a(�Ζ�]׍Lo'���N<卣�8�_^L�2�2�&24���P��Z�*��b��`k9���4.^��Ȑ�t��lo���X�f��4515���G8q�8����������J�6lX�([���jl����t�n~\��)B}�`k�dr\��n�ܞ^ý�qfc{\j��qf��	Ǧ���8
'�!R�?��n:z�0Hv"�'z�!,X��w1�+q�;�ӟj�E*�$Y�Q�2m-hG��=/D�!�!��Ƨϙ�}�*d"�=�ƃ��x�E!=���A̘2-5'�>�5DmV��.�՚a@�HLqצ��b������h�{�D���X�XK������h2ǏǮ]�@���صu��U���KQPP B!$7bmX�>N?��̝;W9O��Km��DӻW��k��p,+u�x��������X�Q<tv�gݐȡ��xJ]k'�F�EA]������VB�2U9�e�XZC bp�ъU�R�J&X�ZF�*dP"COHg�7o��^<��� ����G��/��u7߈q�G��0�z`�M��5�f_��d����:�8�d����&����{;��a>m��fc���Ә���F�t�%�i�o�＇��z��E�/\}�����NaJ?��7�T	���ʘ�.�%�H���`�͠V��Η��e�!�����1C��)N�*kϠ����>EJ���M��ꕋ�)M�ҳX{� �W��]�U�{b�{��ܣY���|(v�,ȂX?������ ���[���ӠA����"���$�8q�^���8���<t!�?9]Y��Y�֖��d�СJ������Rt�.hwɞ��!�j6��k����ΤuC+�X����	3;�94��y�`�L��z]��\���\�J4�kS܍b��`�&2h[&&2º�{J���H6�u��ȑ#x��h��R�����������/����V/��}�=��jݬ�ɩ��֎�dޤ��7b�D���o����W&���_��ƍ�2��mX�w���8��nT�I�r����[oU�T�0��-tuwV�K��� TI�)Yz��0�D�Z{8�!���C�����Ϣ�8uJ�_����?!w���|�R|��L�&wqJ���O�;!���:�P4E��	]��5D}�{0�f���F�?�dŮ����o"W	(�1f��=���t{3f�P2W�ZE�.Kiij�;��^��ӧ�B�};wc���9�N
�f�L�<��Z�W����/~��<���&wY�P̧LoOQ7�.��b�Gu��q!,��^hp'iaC�@��Ztt}@i�۵FwU��&3��4����V�2&1Ėu���I���ԽD���2�2����w�m����/��H���{�D���p���g^<41��-�S�&M���}��i�������홅�7��D���{'۴�z��n:֖���X�oz�3֫�b�����O>ڀ#�d7���H`���8�M�N��۵g[��s��`\����IA��v���"!����ɭW+	�xm�~W�����2Mfr���$w��	!����� n�4��5�:��nh4��ꆁP�~��#m�0bt7��wH�z�{dU{�XZzc-��K/�ѣG�_�$;W�?ڈ�'��slkv�BHwikkæ�*]EHvs�]waٲe[t�.hoښ`<+fj��eu�����v�h��n��>��W�Y7$ɡ����C�A̛2Շ$i�C�hpWD*!V)�Z�J��`4��S�-U�
G?�ӑ�`w=?��V���Ã>�S�NaӦM �ˑC�������3�2}��I��^�#ce#�}-���k5ݗ�C-�����5��ȭ�����o}loHm�o�}s~zozq�M�=jNWc�{�q��Hv3z�h��?��|�2C�21�kE*�8��Vf-�Ȕ*�!�
V�����!��^�.���/��r����q�Ϟw�ܮ"L��<��뗚�&w1��y�&wB�!|P�s��E�����=Z�D��ω)����ƚ��XWR7�c4�{���6�3�կ~'O���������#����9矇!Æ�B�ʓ��������݈s��}�s�������6d�ˌ�aX&uCuj��?'��Z2s{��]�%y]e�����d��N��+�kF����-1�A�v01�!bj���S�U�p�ܵ-�P�2E��z?���J{�;���^Z[Z���	�/�%�]���|O��5����k��LVwlvnX�4f�C��pg�|�u��5la���s;�צ�-���arw��c���w�:���S�g/�m�̶�%%%x��G1a������D*c{A���(X�ZS�۵"�jt���!���ŤQ��䷮L9���_�8���ٱ<��k�V{�u�&�/_�P���N!=���!̟2A5KS7��Le&w��5���H0���Y��vHk���ab0V ��"�r�&�F�/fv�*�����Ǐcݺu �KKS3�]�&f̙��sg���!����=�wb����\|�Ÿ��L�9�0����2�^A�SQñ��C����˳4+h^743�ñ&�D9�$54����
�@�H��Z�Rڵ��JIm�ܓ�UZ�J[�5���T��Ƞ[;�(7��8?f�<�����;�����l��	�9�kn���=�.����X�H�f_���V�k�fe�c�3�g����؞��ng�s������;��=���l\����@�8�衇�hѢ�	PZ�����خ~j&3���0��
f	F�J�fP*Ti��(RB!=����ˊѧ� �����%%��k��k"��^w����	!�g�jE׍.U8���ܤ�X��a �Zu��U�;�u�x�0~���nOW�΍mtw?��Y\\�tݻ�s�N��E�}�ںU�*�d�y(.)!���MM���Q]YB�̙��~��kZ2����mĉ��5�N��C�����3VC4{XMn���S��uC�IRC�;I+�Ot�)��RsR���L[�)Q�{ fpW��D�J+X�S�]"CT����	&w��Tx!n���s��G��ի�/��T���s��k��EX|�����wFSk�v�f�LNmO=z�ޘ�3�p�d�f�k�72�`����Fg�o6֋��3�c����7(�~���~;���j����2���==Zc{�ܞ*}A+X�j�Amk�Dc�Q��ۃ�!���g/���SG����o���lG���o�*��^���~��?��w@!$�	v{ۇaL�AC��\������E��0��H����ƚ���VX��9Z7�c=+k�^�E���'�?�:�Њl���)�����xٹ9f4!�'=xX�v�{�5��F���{��^��`��񚠾fh��n���vh��nflW�C� v�C(L�!��$�y���(\���L��	V�x���&�!�X%H�Ȁ�K�D�G�S�exe`�2饗��ѣ��/~B���ۯ����e����A����O�0�ה�.���X��պ��� d�2�D�ý��N_�ߩ�ˡ9ߖ�^:�:��CG{����@����_��~��ʹ��_F�t���T�Jan�	Vj�A}�A}kA5�=e���k��H��u(B� !��sҿO�1"�}կ^A�Y��4��}Ҩ� ��3�q*��SFG��D��^����jpW놱���y�g�����b�BE��1������<K��D�ꊓ'OV��x�477�d7mmmX��;?y",9y���B�k��HII	֬Y�	&��������Y���u�XH^C4��uB㼾n�t6�
�������C�a�~�ۉux5A�NmK'ꇍGq}��Š*T��d&�@�����rbI�r�J+R�%2h���8Kd�� 姙�l��_�2�;���<����Y|��q��Y�1�X���{Cj���+����p������ՙaݹ	^��f7=��nnp�p/��g�홅h'�q�8�x��,[���{�r]�=��nu2c���l�����a�մ�&0����S{L�����D��!㱻��vB!�����w�y-m����}��;y$!��|�8V���Eꁚ��1�]\�����X7T��dݟ��B�k*OrWǨZ�{�XN�ᗙ�l����Ê+��SOQW%
�����J,^�C�!�b��Q/\�z5�>�l�k~^���-��BM1Z������e���a0�v(��l�vD���x퐰+w����N|�CA�2y8��N�����hnOl;Mtb�X%0�ݵ��
VP��Q�y"��Ft���"N"��>466��7ߴ�^^�??�Qʯ����_���w���/���;w��硸�HY��Ԅ��:�����[7��8���6���X�n�wf��t�II-����d�������[�^{C]�=s~�m�ؽ���vԛ�߳���T��ĉ{C}}�}Y;.{���D�������jٰn�D]*�nolhH�	;7BX;.����52�N9��X۽�x�g�����YGE�P�yK{{;�|^ڻ�曻>w���i�'.VS�vq�V�w?�U(?���$���>���χ_�y�������O��$~�$�L��-L���꒰������ۓ�jRۃ�-�UQq	^>�[��B�<�ob��S�Cs��!��P�B�б(�/ӥ��?�S�՚���5�Kꅪ�]`���ؖ4�=Ffc��=7�o��F?~�=�M�DA���]�&Ϙ����5B!Z:���vnݎ};w�<�����q�W�fnO����z�>�hjצ�'�ڵݝk��a01 ˬ���VN��vjz�4��x�D	���E(Y�A�ԮNc�U@Me�Ls�D!V���Q�h��D�`%�����*��vaa!V�Z���zlݺ��~�4����k�~��t���#8������a�СhinAcC�b�غ$�qc�~fӆz���|�E[��ܬ�M��O�e����mm�kO<9vh"���"�Q���v��ܺ����[��wb�M����l������ar>sƅ�s;{��{�޳u#��}%?~apW���3��kMv���Hji��õ%������;���?݈�w񹓗��Z�\�쵋���=�����w�Z���{ޭ�����M|Nn��9�?�8�����}v�X�"T�J�� KaH&TS۵U*QJL�F�c���dz;!��ۨoj�/��!�7Y8��'�@sm�i�gY�gm(����
h�?G��dwy�P�v�!�]yN+qfO0��y��q�m����/��2� ���������EO�?��뵧SG=v�0j*�0a�d��(�DHʉ#���n������D�o���߽��o��Wj"A��|�	�Ų����c�9>�PD�د߽�Ջ0��OzyO�����OIQQ�k��s�}�W�N��D�������������կ~Uw�\&�۽4�[݆�^h��YR7��e�Xj�gY���ܮ���aHq�3d^-���؇w��͝83l,
�*t"U�wm���堚��$��*B$�=�S�Z"�T*�����5k��������S�8�i�&��!T	����ɛ_�]��߽��[���Y��`�ĉ=v,����e~�:�|\dy]m-�M+e�Xm�ߵ3����_����������ʏK�5cƍ���:|���%��uu5vL��zj����/�W>뇍�r,\x�F�k>Z�2����7ld��m��-��Ò%}�����Ү��\"�Ю�w/>oR�!.��;0d�?mW;:�1x�Ю��/�����.���ڃ�[�)�^�
%~}��y������]|�t�������Į��"@���d���0���5"��X�����^�Ҷ���^2d6���N!��FN�4*��B�ۼq����S�3�ݟS���X��������o��ѥd5C�*\��n�R��\��]�Q�K�9�-����{�Euu5�}�]K��K���������kW�~�ڿ�϶O�`��0i�d��=h�����oȫS���e����j���(��p�|�o�]h��ί����]�ep�h~����&�����3�o>�D���طk�'�Cu��v��{�ﺡ_��<S�u�K.�w�u�'`��9����)|X�0��6�ai뇪��X;������A��Y�Pch�.���Û���e�xH�w�+o�IC�\_�`l�ލBUlL@�r0'�N"�*X�q�v0]BS:�.�H�|�'��ɓ'A��J���#K3fʹ��sS�u��s���c2٦U�sdp��ɍ�V��vƆ��c�پ,�ȅ��S��/���a��zeBw~�qq�Ѧ������{�1̛7/#��~������Gj\��='�&�P%K_�����4wM�BP�jдŠ$�]��=,9(RB!���:UB��Զt�a�X՗'��w�Fh�j�ܕZa4�],�u��j�9�5��녑e=�ޗ
7�)�Wy��X�۶mK�_�W���j&~���ӹ��������cJ(Va�?)ڂ����/~����������p ��������������}��w�����w�~���`,��멯���|���՞�[=?��6�1�~�����z�j�������L�3Ʊ���3l�ޞ�vhLmO��9����kK&w]�1�t܉�W�g�FL쪩]�~P"T��wE�Jh9h����^5�kJ����w~E���D\�R�%F����jf7��6m�br��{���B���[���E�(�ŗ^��b��Rn�����F94���=0���-�Ӝ�niG�&�ݹ�&8}_9����8[�e�F���oc�ݱ�>�奸�i����])�8}�}��.��ߦws"�v�H�
O	I�a��v�@%�Zs�����TA3�*:=�?g�)RB!���&���!��~�>�-�����>��$K;��5�Xj-Q��Y��Ko�LE�P���Y0�nK=��ne~���x��'���!Z��N+uC�C͘3˓dVB!�I::>��͔)S����[�n�'�����YV7ԇb�������X8�y��I-Q���2���3q ��wN6��2t�j*�,��'��Jd�?کN����U\�
�?��63����E����+�����f׶8PV��.�g͙�{ι)5�f_��d�M�fa;�ou�W&rٸ��M�ĥc���LHm�tL&vlη�Z�0��؞Y�"Ŧ�?Dc}�!�o��V�x�aV�D��R��A�J�ޮ����������JLK���'�!��^Ms�>B!���,�5�'��j���&�='����푀�x0V�T�'j�T硽v�h�ᰶ~hnrWɶZ�1c��SO��;�Du�w鬤g"��vE;@���\4�Bz7"�}�����6l�r�8r�Ȍ�����iq{?�uCՖ�։��u�X&�C�#�v(���t�vc����y��x�?��,����N2��+B�e�`47�%��R�c����]�Ȑ��.P�c�0�T�ct/���Pv�/��2�t�����?!2Z����__ā�r\t٧Ч��k�̾��_��fa��{��[v�;}����.h�ؚ9���;1�{eX���[:�.|7�	���wM�r�-��k_��o	M~�^���aӇ�{���P�Mk�	U]���B���h�̿{B!�7��ƛ�!�xKus'����ri �Hs7���X�I�w�#!�=Z/D�(�cuM#:�ZgT��Sk �ZK�1c���):�577�#�����k1���5.��	!�":>�ٱ{��dj;1E$�?���J�{&��Q����6����X74N���ꆲ0,i�0��0�7����*j��4���ლ���WI[P[��IdHl;�(V	T�K��������YKd�$�������,N�>����74�S��ڍ�r,���_�0�ɚ��d��]���3�[k��J����X��+���m���9�����	�������c�ؿu�u $W\qV�X�ܮ�|-~M�<�d�L��`4��MR�թ\��TRڃ&	Ʉ��`%�����DWB!������{B!���� n�<�u5�za�a�N���`,s���8�%�#�n��XV��=�\�Y�F��,��1"���;v����X�t	B!���&���W�����Ĝ��B<��#�?~F��3����J���Jr{b�3��9Yr{Bz��9�t�!��*�>���dG�C�=y<B���S��G�D��0%7�dSm�{\�
 2Dk.	@fr�᷁=���'��z�����������ގ�־���wⲫ���a�Ƹ��nѰ�Yj��͚���:6`\�Ny&�a�S�����u\�n�����a��voiin����p������$cٲeX�z�"Ve���Ix=���Pe�ª�=�<�]�b�3�b0
�[����1�3d^-�ٍB�Z�Y�"���U������V�0!�=����cm'�$)����	D��\�gc�{���/GUU~��S�%�����W�b�䉘�x��1�BH�D�@�����@SS1C�������K2�>���c�����>S��k�C����P����ܜ\�}BxB �)4�����!�4~Z�MM��$U�R1�*�R�܍b��^�\�Ҧ�k��[�N�W$r�}�ݨ����/�B�q��	����a�ًp��磠�@Y.�H��W�{�Z�x{f�$�u+cM���2��-����nB��ku~#�Cýt���uK�E�7U�ۏ���)���b�x��PZZ�"��x7��4�Am1�1�*�T��)z�*3�u	R�J�4�b�_P�7��"!��t��O!$=�h�}�x��V���k�j�0jn7���v��l냱������ֺ?���f�.����466◿�%Iơ�8u�$�,���&�BH��P�l��	�Z��ERr�w��n�vm�+2�Ψ�@2S{�$K��k���ڡ�n��c�C�L:?�@k�ɨ�bHq�IF!ğ������r"�~��ܞ�"w�M��T|��փ�yDl#*X�q��`*�)L�ݙ���W:�����o��d���'6�l�~\z��?Q&ZY3�:6���uh��gvjV�6�;����1܇-��oמ�ܡa��8��Non����>aܤ�&x�=��N�7����Xa֬Y���A�e�A=M��H�{��d����Θ@����a"T�.�����B!�dy�9 �B�����e����IjpO��D�9�wM`���] ��D녝b��Z/T-2�NЛC��!~����wp����3�[��֖l\��U`��g�o�~ ���45���n@剓 $������(�V�I׼�b�Z/t��Z�Ϋu���Iz�����ax���v�4���C$24���Z�*�U�����.��VF�*jt�<9ֈ�b-�!��f����X�fZZZ���T4�����#&N���.���ڀ��l?�M�VM�^��XwL��q�o.��/���kej���*�\`�W��,�xG{{;vmݎ�=��{&�?~<�|�I><#��~`��vui�.%S�*�@��"�v�P�
T��Z�W�hn'�B����|B!�Bc�U���iP�G��`n���a�v���?�L����Ѯ�j�PS7��]0Vo�+
�������܌���/ $�'O��_�Ysgc�Y3,�!��q�w�.�پS9w"�
��r����&|�gBm�����y}0Vb�g��]�ʦ��>��X)j�2s{^׵�ۧD�~����d$o�)��T{�R"�V�R���=�⮊U�&w񝠊LF�J����6��4u����Z2APJ�|߾}����������A��W���CX�d1�,]���x�c��X�\{fa�fe��v}>�c�1�;�?��p篵G����O�9�Oc�ݱ����`Yvlފ��6b��#G�駟VL� 8e¼9�B��؞L����#˂��`t�^�2
Vf�����|0�B�.�YR ��^��B�<��m�c�C����eqC��6F��.P��S%�=�^����j�^��熁]K����������T��֮]BR������T�/���a�� ���8z[6|��3g@�U���Z�s�=�ya&����ߞ��.��l|���[�Mo%�
��Fs����}�����X�]�F����%X�7/��`��`0&E����F�{�!0N���ӸȤMo��,'S�#�����z
=��m�B� N�6~���܅>u	�͘��W��S�u��Cs���ꉉܡ��޾`�U�S��������8����?7��l�߆u۽��T%�l؄��:bq����ӧOO�8�&��R%0Ȧ֓�5˂���Xr{�ւ&BU(ԁ���d�AB!$�`�;!�?Xw�7O��S�k�Zs�����e	��j��!�`�Ȑ�F�e1�|���?�0Z[[����+45���7�Q���^�Ҿ� ��g�e��8y�8�ç>�)<��(((�S��x�j��ݮ�qs{0I�дv(3�w��a�g�4������'����2t$Id�&1hS�uFw��=�� �M��b��*Nz������c1b{�1���C�@�U�.�^���`��	���K0h�`e9S����D�v�f�����X{&r�&zc�֏�����{�4�`��-8T~ �إ��T��3w�\WM�~Mn���Pe.N��������v!P�+��B����<;�hn'�B���B�	!����#��dP�r}����ż4�]ol��H��x=���YL�`,��]��;@3+�|�>}�f��\�6l !Vi�������S1{�<����B!�B�o�۹{��T΍�Ò%K��KJJ2�p�	����$��$ݞ��w}�P��������;L��E�x�H>��g�6<�'͆c�i�h�ԜH�)Z�"UL�
h�+��]�� ����U���"ȉJU.�쮁�O}w�;~�x%�S��9y�$������>�y�`�ҥ(*)���Ooj�4]ܡa=#L�����3�1��X{�{����eq��X��4�{�*N��z���L�Aqq1�x�	�w�y�o2APJ��;	�*��=>Ml/��خM`0�����?����'U�B!�ҿ��B�4��q�1<X&OpOR3T��j��Z7Tky�:!b�X�r�l���j�PS7��o0VO�8p��%j��w�!VZX��8~�(�.^�1�ǁB���@,�%��˜9s��O���Q���ym �6+�1�ǌ횺�ݮ�AC�0h��Y�vDk�ښ�:�`�ژ�N��w��|� W+FG[��؞��`�^�JLq_�JkrH�*�4���$���w��Ϙ1?���p�}��ĉ ��k�Ə�s�v,X���,A^A^��[4�{dl�l��e"�s��e��a	{&r���vƆ���!��{�Ą��Xb�{=v��}��MM �;��GŅ^h�$�X�ռ��@�.��+�F�T���"���Ik�L�jz�Y�����#�L�Ǎ�
��B!$[ط�B�_l>с��Ek���@,Y�P_3L��9��92�k��`,h�2�қ`,;5F�p�>O?��br///!v:�����C0w�BeJ!�]��N+����*�f͚���2$m��t���=^34>:�?���ܩ��������5�Ȳ�O�hn'�A�;�xZ::�?8cC�ʇ�,��htכ޵-�)��P���U@��`$`1u�A�e��	M�`TwSH���̙3�ar���0�O{{;>Z�>vmێ��/ǌY3��s[&r�f]�fa�fe�խ��0�;4�[ܗ=ý�qfcәz.ݦG7789&��~��.��f*O�ĶM�QW[B�K~~��V���.�,2e��ӻ�m��d	��vm�*X��0$�T�V�b�s�D����B�f��蝼4#��/��gF�A{kK�F$�j��j�P��	&w��'��f�Xq �eٝ`,;v?�n�رc�`�{ｗ&w�-���W�b̄q��p>����B�3�MD;�lS��	�.S�Nŏ~�#�9�3C��5?�ǥ5�k�>���±��:��%ʺ>��]��V����Gqi_��@. 
��;hp'=��:0y�8��>��nP���UZ�*'n�7��L��/�݅��S�7i�AU�Q�<�&�L�D���Ǹ���Q]]B�CcC#־�
�oނ�/�#F����p홅���7�{a��s\޼V��[��L������?��8u��aℼ�<<����k�
=�`2�{�nC�%s�>�!���O_P~N��`��BU߁���;B!�d'"��K�-Ŀ���B���]m�01T�܌�P7�>;>[��2�
�S%K������̞	u�t�Ǎ����TQQB��й�>�Iӧbּ9�/( !�{t��cώ]ؿkO�7EHw������3fL�0��a����%c��~���C(V�wy0����ʼ!K�-���<!co����^.���MMq�J���A�$wm�{N ��x��>��*m*�����tu{�pf�N�����?�r��0���׃��r��	����)ӧa���0p����c�3�ݑa�5��Dڞ�<��ƙ�������;iin��m�q����q�0�?���4�[�7۝&0��e��v%���ԞL�����ە���!����ۮ[�la�ޣ�`�!����߸B��-;�_XEqa>!�d/{���:e<�Շ�����f�7�'����fh��R܍Y1�ciɄ��߆�I�&)ݟE���#G@Hw�X��8\qg͛�IӦ*��B�#>?E�p疭hkm!N7/��:1�C{wM喙>'��	�R�V�>w�:���s9�'`_9���{hp'=��N`S�P��iR>4#�
9	�2�{d^/P���`�&���U����h1�ir�c�x�b%�A�hr'N)ۻ���c���X�|���{ީמ�ٙa���{G����Z6�{`7k˰nq��1Lv�	ݫ�����ػc�"��sB�"η��s�!�鎹=~�]\�R���L�jZ�i�n�T��&���"!�8A��ʧ�-tt}�|�'��7��}���_�	�~�Y�w����_��&�!������N\?�?Z�u�B5+Y���n�} ��]�����h���ac�Ygʔ)J��=�܃�Ǐ�����ֆ->F����1w�M��z"!�d�{�ء#ؾy�π������z
'N�V�/��������N��$5�d�Xj�0���I��]���X���
�8Hz����(�1u��Ք'��V�X%����8���9�J�v0�� �"w���I��t��V^�IB֒%K���+W����8A����Y��b΂y(--�-���t�|�d�S����N�
Lm�w#��X�����W����m��Q��}س}�bZ%�rss�b�
�r�-i���%@�"q�=�*uCb{A��`0�b0��U�*jr�J�����in'�b���\<�����O��W?�ɽ�Q�ؒr��#���_��t"n�����N�4�BH�'��ځ8��L$A0Z+�e���؀��YMs7� -P�S�!jk��`,��.��Q�JT�զ�g��]K�u�M����E�g�܉S�q�طs7fΙ�1ƁBH��'���ͨ��!n0b�<����M�=��翹=;C_?�����5Ci�g]8�y0VB�g5���i}����1�Iz����8^���#�T{*!�!���vP�̠m9�#��9�85���b�A���"�6�]��={�Ťt����ҥK��U�V����8E�mo��	��맜|�_��Iױ��,kbVv`nwj"��Z�]Im��/k�쌵g"w�n:֖a��X�7b���:S��Cm'�k�v���6�ban��������7ڻ{�^'0����*��bP+RE�������B������oƷ�<^�hH���܊o]�3�K:�W-��������]��Kp�˒�y��x��� !����Dc'��GIC��(7�Kñr��Xڟ�5C���`,�SM0V$K��J�{�:�v~�̙x��q�����
�8������w���D�n��Nc�'[Pu����0���'?��3,��2��矹]�q�E��$]�Շ��vyb0��n���b��>w��t
�W1L���I��#E�lh1:�ڢTb�A�@��7Ot7�1���@6U�ʌ�q�B�v�س�@FK^��.� ?��z�j&��'g�� [�.�.Y�9�梠Pot7{�[7;5+����Dn��k[4��7܇-����ü#s����-ý�qf��	��mX���]c��r��EsSqq���_��=3��[hr2/O`�$.$����`��)D��D�Ǳ�iڃL` ��}���W܌���Oi3A�tt�K|�g�c�3�FQ�y	A�����bǁ�8|���cz�㮛�'#��>�<:B� ��=�{8����FK��x��f���.ꆱ4�@@7�ĊeɃ�T�;ľ�Bc0V�t@�	�f����E&��gϞ��E�{uu5qa�lmnAmMf/����B�����ؼ��� !n2r�H��>k֬�4����n�.Q녩ñ��v�`,IH���Ϛp�����J��$���Nz$g�;�?8�:+�mL��y�@��"�H�;���@�ʀ�(�R�úm�m`�û�e˖)�=�M��UDz��＇�?܀y�b�����ݳ�v��iJm�gwf�wÄ.]�����n��L6�Jj�a��QzeX��=��;�8z�0��؍3�� �mĹ�+��/|�Ss�ߦt�捩��H*��v{	r�J���T�����.��&����vB!�����/��}�y���n�����U��o��Ƿ^�t܀�"<��-���ߢ�ݛs���"����I���N!�͋�}���"��lV/���1�����������Y���x�~���?�ɔz��ǔj������<� *+�2K����c�c�ј5B魈.����у�A�ۨ��~�ۓ�W�P�&�hl7Io7Ȓ�u�X��a�@,Ӯ�Qs{QI�t0I3�x�ǲ�T&L���Cq� Z%3�'$o;(0
V�w�f02,����{��ݎ��t[�{��ʰr�J��y�E����6l��>Q���-@aA<���,l\�Ԭlc�w&�L4�;�8�ܮ����.��9߳�v�64����P=r��v�Qn���M^^|�A�x㍮�ۍ�mJwk^���x
�F��el��.�$0���*������c9��B�C��u�͸������3x��MX>w�9ﬤ��N���~��_�ۗx�}�B��������BH[0���C1-|P��5��ljv�	Ħ9ڟj�F�{��]�cA�����fBݯ;��t��Ν���E0ֱc�@����N�ʹ����w���N<c��ъ�묳�J��݈�uA+�zc���.��Sw~6�
F:=�u�P4 +dRC4��,�ak��.�I�����h^��������Z#B�[�	V9:�*� V%��b�1�]��F�X*�X7.��{o2�kq[�:�s�ӟ�T��z�xA����f,<{fϟ�$�'`��n��끉<�؀a\��lӥ�s+���zps���7녹�+�<1���<�@Y9�l߅��f����/���W��n��W�(��{=���ęU�������Tg��P0h*Pi�j*�(,*�ߏ�	��^Zۃ�#(��EIQ���N�4�� _I�����?�u}��T'��~H�����7��>~����n�h[ڰꗯ(�8n R�����I���N!D��:�)�ǣ�����sN�4�d�H��1�]npW�\�`��~���y&w;�t7k�"��g�Q�܏9B�Fkt?k�L�;!��&��VU���	�x����s��i�|1�gB���v5��v}�c�C��Za(	��Χ�ʻ>Ob�g�4���0��}�KK�TY��*P��D�J+\A3/o;���݅9��.�H�q@k�Ӧ�G~O���3S�J��%{nѢE�`%�B�z�xE[k+>xo=>ް���ż�PRZ�Jj�U#�w&r���S�}u����wj���rhηe���ƄNs{z�>��+�w�0���/),,�#�<�����U����N��V���I�Z��?Sۍ	:s��H��;$U�����6�T��n���w��/�G& Һ���)ǉ�{�o�w�M�q�d-��)����z\~�4�:y�9��{nT�_�g�N�̧���������@QA�r��?�W.��vҜ��;v؀�chn'�b���N�2y�j+����Qc��!��}h���=G[/��]SY0V$K���&w-^��O��c	����L�%ޠ�G���sgc��� ���Bu�i�پS�����x�ĉ���'ONKMЈ�fu���0,Ӯ�����e'�]]�a5)�J-1U�gY��!���2v�'�A�;��T5�pr�Xj+3Mq7
TV�*y��ؼؗI*Cm�����t���y�#ar?u����v|�a���>c�Y��x!�W�������s{�|k�1ۗ����������n�Dnzs�l}�XK���7������!�|�~�߽�� �k����f�\y�=�ܞ��TI��p�Zv��Z�d)�;h"����N!$5w��_�Ζ
�n�-�oj�W��/<�K�Γ���܅n���v�d>�+N���7�+nH9v��H4�B1��%�h@�r���fh�^7�[�j��z�1Kot�&w7넩�%B���Q1������8v���2l(��>KIv'��L���
{v��	�S�*��&LH���o���y�f�7��S�e�X�k������
:���ϯ�㩿�����
6��SƢ���i"C���wS�;�r�$�AO<�A]7b��2\��=7w�ܘ`u��Q�%��o���c�X�d1��8Іa�y&�a�u��pj7kٰ.]����2gϠl�^�W�|F����s�W\��B������ԈT���!s�J+LY0�ǒ�%)����
B!���;ۻ�K������߽���<��OI����V܀����m ���]��c��Ǫ/]�����N!$)u-!0
Ãe)k�v��j���]��Y�*)��h0VB���jlW�[�N�/���4�O�8QIr�X���!^r��
��|G	Ě:k�Mԛ�!�/�w��cǱ{�Ԝ�!�@t��cǎMKM����0A��Y���!Z��v���h�0�P;4�ծύ��L|�w�kx�"׍폖3�1I�n0���`�vИ�)�iE*�pe��5�DЦ��7��H&�C�܌3���z��I�(߷_y�?�/���l����~�O��f��3֩�ܙaݖ�܃�\1�K��oB��=}�V��w�Q�b��$�_�~x���q�d���ܘ�S�O��0H�Z�E���ݮ�]��`La����ۧ"��3�B��_X�֎ ���������N�����4���ן֡��߿i�o���wᶟ�@s;!���l>�uS&�����f�c����������5Cm�PE1�#^/�w��MF�����3�Nh����0a�y��\��v�!^SW[���>���1e�tL�:��� ��t#jGR��gAH��9s���>f���xF�c>�}0���.Mo�P7L��Tj�A��v]r�!�=g�$l-��������	���������Pe�� �?��Z01�!�t�9�w5�!2&"�DZ*si7��axw��.�܅`�o�>�.�:�<DB��ys0c�,�(����v{���p���Im�n��e�:���n�po:�_�:��CM\�EKAB�������SO���v,JqSd��Ю�W�)��].Ti��*�H��TJr�=s�Q�R��b��P��B!�m~���PR�o��-L�:e�_on�|~�oo(S?L�"���vB!Vy�<�'BsC��f��J��n��ꂑ4wm�P<dI��pT�b1,.��7�H:���:"9T��V�^�m�x�$I���c��]�2s&M����BB�״���B���ݏ��V�N,X����1b����tڽ��S��I��G���#?%��!������ϥ���r�<Hf@�;�U�h�x���T�,�4[�}���P��� ��RD,$���S""��j����=��[�L�8?����裏b��ݰ���^�_�Ȑ����}��/����/Ӈ�݋��n�vqb����رe��<


�4Jm�mhmnQa�/����@юL�������K�HuHb�¤kwg�_��Ȗ�߻��MҒ͎������^�{���ֶk�B����ZT��oe��mZ��L���=?h�������[�345�Q.
��ٵn}]]�{�F�����������~~ר�t~���گJ�wQ7>|�r�5{�l���q�"ju_�R���ZIo�	VR�J1�����O`��O�hn'��"��_�"�q�y�����{WaK�q��G�܋
��k�I�>��N!�.����+�ci����X34v�R+LU34�
��X���`d�z�|zM��zQ'�Ώ=ZIr�ᇱa��.Z[Z�㓭صe;�N�ig�D��@!nS_[���p���rBH�Y�l{�14ȳ�^wֱ�]��!��k�� \��j�0E(�xN���R~��ۃ!��X��aA~>^?Q�u=E�d4��^Ǧc�v�xt���B2$���%�OhD������dE�RS�)�P��Qѩjt(_d���v7'�ūQ�F�駟VX�֭�T�W{{;�@��kէO455�����b�����W�����br�N����c���	f�ƆT�>��&ꖛ{O%&r;�p��;wc���}���t_�Ǌ�QO����Im�.��:�|.>�z�y��k5Mm�"��M��X7X���?���M1ۢ-�ݱU'O����O�R��0�O�:ٗ}��SG�c����i�o��={#�T�Y����������[+����ɼէ�
?_��������a�ԩ%J9]�+,�6e����zc���	T����`4��O����k$�B�����9~>�P~}"t�A�J@zk~�w��𭫗x�/��	!�t������)�?�1��5ø�]�hpW��S������jz��{_�g/�2d~���'���~�-Q��
�;��p*?�R��M�i|X��K�1p�`���k�+�P,A]M-���ǀ ��/�kk��RX�]�kp� ̎�MMhok�e��&���v��3���]����[�練�������x�
D�.�����~�
��-�X˗/W�唖�zV���:�fh�����O�w~քbj��S�������ۃ�������	�ma0�hp'�����i�`45�F��I�)� �A�BJLd0�S���F#�Ơ���v�����='�-p�c�ڵ ��{rߞ��cА��9kf̞�u��P����[2پ����Ec�sý��`q����f5��e"�e��3֡�^:�}úW&x�}�<v�w�E剓 �ofΜ���Ǎ�(e�?�z������v�Im�br׊R�H�.����w�e��`x�"�k�K���F1һ7| &����f�8��߯��8g�8e~�#hmwv�!�������m��y��U�{��տz��TaΤ����t]���w��{x�B!�{l?с�J0��x�Ϥf�c������;�k��iL'HHqWuUu���Yݟ��V�q���S�E�z�)���˰BQQ�����g0�x��_KK�/��;,ī�����S����~H�&MH08
��`��A�?�������%�}|�����o�L�J8ըqc|�����1b�(��tS���;aN�����<3���J�P5�;��~�Z�� �>� �k��ʕ+�s&/k�n����)��Wk�zc�$K��9U8V�`,%KIp77�kk�f����8;*hn'��W"��=�l�����Z������[�փ��t)�5��p¶R�n�ʭ}�5N�??����U�򗿀?�9]��＋M~�ig���ٳt) �M�f�p���������>ֱ1��ذ�����5,��?�7���nѶT$���݇��f�	,\�P�ap��ᾋR�Yǩ�ݙH�OmW1ڭ	TZc�^���/%���)��U������V�T�wq�����7�oI�F�?؍5�Y�cU��D.Y8O}�JL)h�>T�����n��靈����X0u4H��w�~B!$�y�<��'CSmUb��]c;��CM�;��c�t�h��R7�uYqTc{d^����v��v���5k�(]�_x����7Dw��mĎO�`���4}*B1���������v0����?�y�X�B�Q+Sk�F�7��KL�>'Io7�!&�
�܃��ꆚ�a���c&H�A�;�Եvb�(��<�|(���bL�����Fw��] �'��6�|�i�ܭ%2$#BV&�܅P%�-q��?���񝶶6l߼Uy1�ƌ��c%w�;5����%��7����Dn��ō�2��2����p/�	��v��'��Q���U.:	��-[���]���:~	\qaJ�,ǖwjR�%$/�甶�Am�AU�
�No�̫bUp�$�b�e��Ogn|f�L\0o�]�[�<�I|��%x�[WB�Q5s�0��W�;?��l�s�wB!�������b\1��m��ρ�4�d�CH����XO4ܣ(ݟ%i�q��B���0��Q'���Hk}������~�;�'B���W�<��S�`������!�tv�8?rL���3�$�����{��r���2�&�t}o��.ϒ���>�=Y�0e0��Ƃ����=duC�(*.��G���UC�o��Nz5;N1v�xt�ԋPI�)�p�D���-�F�2��(V))��id�jt�orO&�h�$�Jy�.�G�5x�]w)���}�Y�)���B}]v�؉�fb��4d����V�E�'�'�NM�Lm7�=Sۉ�3�gp�� �U���t�ȸꪫ�j�*%��M���8��(#n�TZaJ�b� P�����FD*5�!"P�-CJ�{|Y�ʤ�`�����r�n�%���י�U�u-�6fH���L	����уAHo��x5!�B���-��#0��@��s `�t����;�6��?��v�x�+쐰)Ф(�B��=K

m�(P6!�UF_(e�Zx�{�@�jl'�^v�x˒��邏�Nw��>Yϧ=t����$ǖN����~��.���.�r����z�\�Rc���,�ǨkkVHu�{FF�=�\��}����7"$��t���#??���M��((*!$��ڵE��K{k�t]B�]���wu�	'H�J�T���H�z���js���5������ĶөNm7��,�d���a|3X5�y��EĞ��NF=�Z�qt��q�zC��l�W�BZ���G�R��*훟^��xc�\����G�h��=�w�#���>UUU��[�p8@�]�7_}--��J�ݎ;`�v� '7W�o�Dn�ֹ��#Rzhc�o46V��ǆdX�8��qY} z�&ڰNc�9"ma��.���2m�ؚc�=�w�����fn���%�Sjc�B��S�������*c�,X�*Y�r���z������6�#������� �.�BC�NB!�$��nr����m�n���Ak��-��;?�F)�J�{���9��+6f�D�詧�*%��~��� ��U�W�R�k&Jan���ːckV�B{�2��-��͕��~��1�Z�:��j���v�H�۵�X�����r9�����⚤��	��4��B�;I	���Ay������-�He0���*�H%�*���5�GSp��������xΜ97n���Zlٲ�؍�M����ه������v�v��ﯲ%�Es{�l�&�P�F�0��s������P��sń�:��ƈ����eXٶ\*�����;"���:�,��`�[Zm!+ZsY�<��T�R{Au�'�����ss�6yA^ă����CNB!��	�BI4o��0�y�;ש뀊��1���������u�:�ۛ����,cy�%O��x�8�s<�cPYY�����5Cb;�T�o��
�k��8��@������X�b%ּ��bG���p�Wbƌ1�Zs��Hj�ʚ�|�.�U�X�Zb8�}�X:�C���ҭN�P����k��R�.{C�;I	z�����b���`e*PV�m`*���J���Ms����F�cl���]�]M����փ�_~96l�W;zBd�貖Vi)(,@�6۠a�f�W�������O�z�&���uǆdX�8.���s��	=&�T�gk7V,[.-b] ރr����w��K/�!��ւV��UȲz>�ߢ��L��k/(�	�In)�3��R�v���BO�H`�HE!$��ݴ'r�(KB!$q��<��/�@_o�B�АC���v~�� /ݣY�k�R������E��?ۥ��qӧO�m��&�׭cj.�B��b)(,���F�75 7/��䣷��m�280����ۉm����u�]�)S�Ĵ>hu\<j�њ�_/������ImW������|Fv���nnn�j�y#�/�e��aC�-`%��-.T�5����/@� X
�J)X��ƕ�MeP
Wfo��4w(�*��M�b]�	��EOd����cB�������e�]��K��;��݃%_-��¢"4o���n;���-]F���i��9>&x��qKm7k�1Li��v�0�=|�����#4oڰ�$eee�ꪫ���Zq�����]ml4��R��U��v��@��\N�}����J��A�sB!�G�G�X��Ԗ�B!$Q:��bk�f�y��B4����c��=�=�����I�}j�A���)�rh�/�@�Sit���]�Us�ո]w�,�j�--- Į�tw㻯���K�Eiyj��P[_��lB�ːÁ5�V��u6���J��	�+;�#���?a�ĉa����E����KknW��C�P,�ڡ?+0�%�`��X.��v��azF:>��!�0�;|%)Ň+�0{�D86��ܮ�` ZiR�I���u�X�V�T��<���4���(�����p�B��Β%K@H2нu+���KiWV��m&�y�IRjS�Ck�𘥶�-�38U��4���E)aj_�f��!��d�n�V���x���^j�����`)}A��`�^Л�>r�?��X�r*��}%�x��B�mX��wB!�$�[\���GY_��g�1#��%hQY3�z�6�][s�Q��)�B��f�X������<O?zsk�4i��\q�����A����"dG,�|��U���Ԁ��Zdd��C���ڕ��޶��C�t�@,�*//�g�/�u�X���vm�0�P,�`,�v������N�E̵&s"�v3�$��%)ǫ-i8��}[:B���o[���\y���c��B�ʠ��'�*�փj��ԂM���UTTছn���_����$��:���O>Cye&66�q�fz���10��*�=n��n��ذnql��|��z�ƎV���NFF��T7�k1�����-m��"}a�zr�����S���z�vi�SJ�{VN�\W��B!�.���!�B��b�f5�c��=�.h1(K��[3���:���ʘi�w����1�����B�[�|��u��7��k���B��;,�Ų$�KL��Am�DT���|���!4~Q7\Ѷ\
�FSB���3g���/GAA���V�%��.�c`n�	�r[�k���c��vhhn7Jpr�=��[��E��I��y����<X����J��nx�O����4�X�Oe�o�I"��X��V�9z���+紛x�1�X
V��ŒX%�>��3 $ِīu�勏?���'5���	E%Ŋq�G��Je6N�=��qFc�����c��n��ݛh�z����X�zM�d�0m�4)����4,q�l�h0����򺜾�m+,�A?�]���i/('0i1h R	��BW?E*B!�b�Z�	!�b^ku��*�u���C���5��!������2�u)����%5�x�+**�7܀;��=�I&���޶LZ233QY=�k�Q]W��Z���#o��׮ê�X�r�����d���y睇��,[��=&�㭝�_Ԛ��B���cik��`,o(��klw��U�v��aA�x<�B�I.xuKR���n|�W��ۥp]A*�p��U��,V	dQ)M��}:��JNv����j�{�D�h��q�O�`_NN�ϟ�	&`��;!Ɋ2ٽ���M�k���q�����c��nuRc�}�&���Fj��?{LL�LmNOw։�����ظ1ed�1g�\p����K2�O�*��#��/LI[P�����e
��8e�ܮm-�Kp7I`P�/hD*�s[�к�׺�B��'߷�p�ٙ���#�k6mIr�2p繇c�m�a'����7����@�G]e�GG'}�l��!���<��b��ǴF(п߬f�4��������r0t�?�!�z�@]���=�Z^(��D�����/DYY��>����Dh�"�G,��?��k�뤄wa~'���0���9�Ծb�/X��dE\��{�8��c�^��j{f�en���]��6��ە�XnˡXz���ڡ���:uk��.����C�+,�K#�{I6hp')˲�NT�L���V]1*����m�4����܁�7�1
C�R����^�M��2����l���O<uuu��k���B������E��s��P�0�#���jT�}�V��0�GhX�:�;����o�T	7����[<߮��X�j��l�`�$]�k�y���SNAzzzL�'�s�K���\������j��G��On�����U"��e��n�d�����	!�ؓ�Vlĉ���^r��1�p���^ŏ+6���ń'.�5�Mi�y��0��'��+A�AfF:���8�gۃ�Y�ُ8�ƿ�bF>B�����K_"V#���v~V��KrW�jס������v{��k�ꚡ�h��U'�w�Phg��~:���q��ף��_>"ɋ�庇�ݮ���	���mvN!�����DJ;;=�ф�^s饗b�̙Q���K�Q=�c��+���._��bOm7KnW�إ��r����v����>Q;��sNI6hp')ͧ��8��C�jJ�zPF_��jS^�
aK��.��
V����Oq��*2���.�����*U�NBT4+y{���X�`���J������B_~��i����rm�D���kF[7����n5���o�	>$úű����n�\����p8ذf6�[�5+Wa� ��Fd�ꗿ���K�~� PE{\,����v�X5�M\P%2�ۇu�)��]���t��+���:K��2<�*>Q�p�B�	�^� �4����C�~�4���l.�۹v%+3g��6��3Es;!$)X�Չ��ZT-�s����4c����.���P3Ԇcy����n�S�w�ۃciI�:a(��QO<�����Ϣf�b�
���q����"(*)���jL��W&B��֮-�/�lڰ��6jkkq��bʔ)q�Z��N�v-�ڡ:�s?�uCM(V���q0�6K�jk��±��� �k�م�$'4�����a�T��΍~Qʤ��@u_��� h[z��i��e��PR�;�b�[ό�ڡ��nr�Q��<y2.\����
_�5m�٭[����>����QZV�ꉵ���AyU�d�Wb��n4������>Xk��,�M�a}�����ذ�׮�:7u���LHUU.��2L�:5*�پx���=&������v� ���D*���/Py�+e��^��P�kn�?'/o�.y<L�!�b��o���n��ogs�?�ً�4�B��o�:1�i"�|u7+FwM0X�л#���B@��?'��]�Ь�w��W3\�d	M�X~���())AgG�dx/���2�z����v��[�FJm'd���{H�6�|v�ZKs�q�P���P,m�мn�2�҆b�B����N�"B ��5��6��I��+U��$�E+�0�"��}���`B����h=x*}���Ms��X%����C3�kG�ūP��<����jjj�$��n�	���:�dTӱi��|����kJiy��Q3�cǍ�1Fj"w�1�p��a=s{��{���0��jl2���#	R"�}kg�n�
BR��w�]�D;�x
Tј#��h�M��ւ�@�1�����{o���T�P5f�i|�[��A'!�B�I�ȅ��<�ڌd�o.�+7nAuy1!$YX$��&U��cm�Z�aѰf���ѕ�U�۳;����L�J�Q'�em1�8����>�pz���n�[o�BF#BOl�o���Za��T��B��RVY���dG�΋���"k���~O�hgƌ�?>
�^4�g�:b��|.��]��9�P,m0�����t�nn����j�B��$^Bl���W=��9k%����*x��r"��\���5�q�}�u��X�ǟ���=R�)�BT(iV�H����J<�� $�G>���O?Gn^���0���UU(X|46��`հ��<4ý�qF��&ڰ>ڌ�=���q�zlX�}���}��� $U�5k.�袸Tf�!J�s����MaP-r�A��ւ��԰"}����R
Q��T��6�7�}#��B�>7�y���H�oq�[�bnx�m�t�)�\�B��yyYfO(B_owj�r�P�ߚ�D��Y�v�_p���9��Dc\��D��0�766⡇u�:!J�����SZ��7+;�+QQU��	�_�ZIN��X֬Cff&zuDBF3���8��q�YgI��v�Z����q�z��X?4�2�
��w~��c���f5�`����b�cYL\.�$4�⥽˅�	Q5���]Z���vT�����e��*��8�4�!XY9o��ą��~�;)��[nA__I%���}����,�WV����U(-/Hm��z�1�plH�u�c#5��=��� �1�c�Ftl؈�k֡����2�5��3ΐ�F֎��9kn����ܮMafn7N`��/�]N_p��a��E{A�6��V��	!�}��7N>x���>�a%�uv#�8�\����؋�~X�_�T�]"��d�1�����W�������.0���=�jñ���r�g!^�[����#���پX�q�Itk�Bk�7o���q뭷bpp������U�WH����PJu/KU�.DlJOw�T?ܸ�!
/!�@nn��u���^�*�C}��h���S�������"Ky_��XN���kvW�ӫ�۳�2�r1��$?4��`�!�Ѐ�ͭH3Ɠ�` V�&'2��Fw��.��`8�g�����'��ڂ�M�b]�q����c"�C�>��={�l�����C[�H��t`����"�Uƣ���W^(X5|Gj"7����#2�GjΏ�	=&x;!>�uut�c�&tlڄM�7b�����Ÿ��q�A|��.������v�X��Z�{k]�
L`P����)�0\�����k��R�S%��dg̘��S���C!	f�]�p�)�:�1��'$�9!z\��[җ "}��َq�!{�B���n��3��e�&w����f���3���LMHr=�J�gar��e�/�j���lΜ9����j�k׮!��0�eyK��-�A�V��ld�XcKǁ�D��Z+u}&$թ����W^��w�=�B�}ў#Q�v�h��҆b����͂�ԡX�ڡ�.h��4����{�EF4�����9qDs:V��z	*b�S��%b��KRʖ��o�R"�ț���b ���c���.���eeߔ)Sp��wK-?��CB<�+�-���b��.�,az[Z��#5���jV7�8���!�{��a=���@Wg'6m��Q���7�	ѥ��W]uv�qǄ
Tf��������J�*����@�m1����HYp9-e�*��v������ ������=��w��ڎ�&`��d�wG�Bj+Jp��DzC�k؍��~��vb�s���O~�x���ੋ�^��t>;p���Ď�� �$/?lt���%=��:`�:a`��5C�����<4A��?����h��徽����w���Z,^���2���Lx���Eiy���-+��!�Dh�;:�)B�F��M�08���(�k��p�e�I&��Z�:.Z�vm��(K�*�����`,U=�gl^;42��eKa3~Z9BF��$D��G5U��s��T��R�J�������+�7Y(E*]�J�S)�x�e�z4��X	V��UUU��o�=��򗿀Ȗ�-�������,��t��Ri;N������î�bal��{�a�1��s�HU�ҹ]�G����� !$83f̐��E{d��can����ZjĩP�����~mr{0S��1���Moţ7V�9l��{B!�_Z��;	�/}��:�����/:S�ƃ�6�Y#�G�� 7��^�����؅�]�!�=�p���Nt��>Y�ġM��l�\'ԯ%��k���>��B����]{�x���2N�z�vκ�:�y睸�;��/��At�Uv�/��E��]$���,��} �9�]��E���M��N��c��y睇��<�55�v�k{ј#u�P���n���2�V%�����b9��|�Js;]��N�B�yey6�.BOw�D�Ȣ�^��g�˻\���ъU�M��f3�{��	��OolNN�9����㦛nB__!�8X�r������zM�e��U<��8����=ѩ�FccaBOVc��=�-]]����eC�0kBB#=='�t�͛�����Tf�%^��ܮ0�+D+���<�!P�2Kn7j/(��>arW,���eO��øC!$:4M(�3W����|�[�?�T����1���&r�ɿ���	A�}�t5n��� �BF;���qԤ	��X�>���fx��ݟ[�9����><����5�"\�{2���!�FͰ��@JF�f�m$��� Ӄ	�"�f�vm����e�}���R]���XZ�R�1��L����������)���#:��J�%���.��9s���h��b�Ϯu�`�ve��j(�Y0�6�ݿ�
bb7^�˪��R~��>hp'Ā'�A�8�S8 ���P�KS�������,UG���
c�,P���9!�����E��hr��>�v�a����5�\���vB�#^�6�� -J���%A�d�X��YJJP4�Y��vӖ��~wk�vC[�ű�2�'��]�����{�G��:r۳e+�n���(PTT��.���կ�A�*P���]~U0�kZ���0lA�
������ �2c"ڻ� �2�ر�/�p
�\��o��9�r2�ĥs��@��6�C�:�w����x�6IلBH�y�5�3q,��v�
--�k�i�z�<�}A�?k���Z��/�������j&�h���_��ט8q"���:�]��s���i�Fi������,E%|vv6��D���oDOw7�:;%#��)2���𨨨��W^�}��Ǵ��ݶK0sD�����ܮJm�1��c�c���=�C�3��v��XP2/��LF'��&Ą�=.��[�F,W��C� �X�6���Ղ�b.e"����6-M6��s�E+y�d�����'oO�:w�}�dr���/A����^iY�J�ʼ��P�
E�C

QP\(����&x�8Sۭ�C�{�v�Hi
==�[af�����7�������&\u�U�i��l%P��øP��򺮹ݻmM��7��t�,P)�����r��	!d43��/�x*���)���鹪���Km)���~J
rq��g��2����t�BI���7�a���dٴ@���^��$w�~�����q�F.����R�����ќ��|��gt>y{��ƽ��+��,YBHh]U$v�EIfV��I���zaq1

@�|%��[��Xb]d�I���~�	�»t��W���.�^(cen�GQ������B���:�X.ej�y�0�۳�v�����|Nq3���Nhp'$?lt���%=�*Jm`N����|��/Zi�ӛ_Nd��vЛ� ��!~�E-Zɷ�`r6� ��������]w݅�z�=�X\L����[��X��_�
�'h!7/y#�"�!g��]n��������L��}}�"��==ҿ����[f̘��/��������a������]O�ro-^{As�rqh��J밨�!�$#"�z�M�y�
�Uc����w����Z��$��o��a_Z�q�>�Qz�#��Y?�e��A�=��7x���BI5�����
�3�=�X�j��f��_3LS��60r��8&�V"b	�����h���U3��)�w�y'���?�7� !$r�iO��.���-d�����/�-��f��ė���vw�{d������&��E-�9s�����/�M%��>;��ܮ�'Z��ܝ��v�N��J�зx��c�����Jt�3��^hp'���t�Цzu.W�K�~#|��P�o��`�fl���7�+��������Oo�H%>�s�����oFg'Ӫ���P6��[��S�}
û0���`�V��fdf�9�Dvn�s�G��s���TJmY088���~i]�O��}���^���vB�A���֩����N;YYY�5���/��v�5���]��`��n����&��c�{�b"V���s��[��-!�{�v���sמ���c-#���{űx{qn}�}|��*Da����_�}v�έ}�����G߃�NƤ��].}h!��Te�f'J��c�`+���*k��BE�PB�ˋ�-Yc�e������J������'R��=�mr�Ƹx�(����p�u�a�w��@�>��Atl˦�}�Y�RmP,��y��37/ϳ^�/ൺ11F�Ɖ�܉[����W
����ꮄ���7�v���裏�y�d��vh�q��9xoC0�{;Ak�=+��5À`,�SSC�	Ͳ�%�^�Q�U[�@�h�wB,�j�s���ױF��e*�Vz�)��g+!N�$2$���q�h�Yfs��+��3g����_=����]B����,X�OCMZ�H{��͑��"R<K�d*��ʔZ ���v�ȭxM��&�1H�H�AE��.}�Y�*#��Q���!鹉u�����W�ş}A�:!I��s�E��?�y��P�&�x���B�B�@e�^Pafwi��J�IW��i/�_T���sC�r!���b}��/x�⣱�v�����k���w�F��؊����}'����A�Fާ�F>�de�?��{��F>�T�b���J����.�6v���.���翣��B!$��z�J���`\�Z/�����a���W@�PO���&�a���4���]�#i!����-Z9o4��OolFF�Ν���f��r�JB⇨�uun�=�����˗j��6(��R�07٢F��#m���ъР�җ� ,����R��>)(�uEB�ŤI�p饗bʔ)��&���1��8��]Q?�N8���~0�q�g=�z�P,����,����~F��!1���8���]�+-Z�'V�o4�}kҢ7�v[W�&�`s�aV�D��~��q�}�a��x�@I�8#�p�8cFa���"BF�3��#�+�ۥU!�9�oҪ͉��[!�mq��c�f8��RA���a�}��%�\������Nњ'�sDz�`�vY�����[k�����ւ���ZAʡ�^PY�Z_�A'_�	!d4�~s���	\u�/qƬ=�JflS[.-�d�5���6����p�AR����;���Vl!�B���\�=i"�V�X�3��y����ϊ�fݟ�Z��5�[q��8F���4��]�����n�/�j������}�������3��}B��t{{z�%77�g�#=#C��yB������Δñ���R ���c�Z�t��M��Y^<N��%���+�-��"K�';Ep�'KQ����)��}}} �$��bƌR0Vyy��ꁱؗps�X��
��v��v��v��}�5[����%�7�:��T�X�bz�D��b�剐��˝�WV���b��l����Y���X%�T~�*����.��&�{4�	�[XX��.��'O�-������ �!�yj�x}���!��!��D��9�#	���3Ϊ�= ���*P��u�yr�YCff>���~�T�2�y���7����p�y��� vd�����m����@I uX�ُ �B���[ܘ�4}�k��Bx����a�qP����0�~��uQ#T���55C�^(��&w�]�F���ت�*�z�x���q���K�!$y�%�b�A�_����7_}mx�X�V��B�����78�䓥����26��A�sDfnG@�PU7T�CKn���S�=uC]�u:?�M��K�DBR�		�'�ֆ�?nHj�$�JJ�JO�ҊW��Ei���ʠw3��d�O���.Hf���|�̣7V,�g�Fcc#�������B!$���R���P�LV��l����:�j��X���خ'L9t�)���?�j�jK��<!�؛~���A���#���u�o~��.�6w����B!d�#L�/�e����г�S�O*�i��Z�j��z�z|�=�Lir�Ɗ����_h���
e��"����O�v�m�믿�֭!��s��,B�����_,u~���ݶS]1����ncs�\7��jð̌�RJ����21��u}XF�?�KJ�b+�$��o<!a��_�T`��U��R�R
VZ�J�R���&bbmr�:.Z�������X�G�)�"���;��{�-B����G���L⹋o����f$�Km��=m���{��}�'��ً��,('�T�������߼�;���Ĺ���0_o�N��]\7̟?_��\"�졌����9��#1�%/��*��]��*��v=�J���sn�mď��@!dt�j�q����1�p�Ȓ>&1א2Α����~w=�!��B!$�^YU�Y������ӌ�?k���ݟ�8wh,و0���
�Fݟ������q�d���x���?�	�/���Bh�@�;��n�Ν����5��G�!$�T�����g��$�D�މ������V�s�=q�e�a����b_2����XúF�p�>��u�y�Ex}U>��mIjA�;!a�b��ٵh�2�DO�� ^��E*�`�qh��.&�h���>A�c��eeeR���/���o����P�ݎ7�:nn.#b�lǘ��.>�����@B�/~/�sO��]����l6u$(A����|NN��X�H�ss�5�/-,�������A��&+�]�6{�8�쳥ߕh	R�k�}�6��/ȷ����ݥ����Q�-u*��2XҀ/���N!��k؍[������?������C������M�ZB!���㝍c1}���<��ݟ�5C�Ρ\I�ޤ)��v��Z;4���a�7��k� Zckjj�`�<��cx��'uCIm�M��5���D�_6��g���;M��"e��e�y"�ŹU�N��]��\��¯����x�s�?�x�v�i�Aj�0��2֎�A+���06�{������j��QZ��0,E�g�w;;;�m�^G����$
�	���68�[݈��6�E����)S�*M9��1}�J�� �b���"�w���<�#�����o�w�}B!����*���X�Ad�n�6����4������t�,�]�;t*������[)PBH*��+1��p���9�!'+>�m��>���x��/0�JL B!��d��o_eUbJ�*_��\/��Ú�����Q��J����^3�+�`�͛�����rV�^�;V��!���Y*Q�O�sO��Δ�?{�7)봉 �=�k~"��E8S��'��NxG������,��uuu��������P�&�>he����$�]�خ���h��\N]��Q�P^���1i�z`<6�&.X��DB�;!���!��P���eҶO�J�Or74���	������`&w�خ]��`lA4��k����;����~�BIM�u�hK|����v�
Tf�b9.�v3c�O�2I`0La�Kn&��%�t�oI\�B!�g���mϼ��}��LE��q1=ߏ����-A�@b
}�B!���.
*jQ���ݟ5چ�n(��69��O^�����m^�W�0��+����ӦMCss3n��V���{���BI=���̙3q����"f��P�M�:��9�)������:>�t}�����!���X�ވe����.4��Y����1�Ѯ��dCS���4���U�@%t
WJ�� �g�B�D�H,�vAA�ϟ�]v�w�y'z{{A!���A$!�|��8��ӣ�V0�c�/�v+���6��jH#L��e�J�ܮIa([�Z�A!�:���?!�BI.D�������k����oB�'�!�w���c���5C9�R�x����.HthV4�=�h;a�)���g��]w�B!��&���8��3q�	'HI�^;��h�ۣ��Y��vq(C��u��M��J��IjC�;!Q��7�4O@_�i[����1��ݕU`���خ$��_q�L�;
Vf��h_$c��%�<�l����z|�� �B��gҤI��K�/�E"@i�)^y���=����͠˰��X��vEC~Q1^Y���!�B!���瓕C��� w�2i;�[/T�e�A�P���ݻ���]`^3t{M�z�����ܵ��ء��X+�fdd`�ܹ�~��4����BI�5���^�w�1ej��#��ve�0h0VaX���55D�XJ��2��	����(��t�T��΍>�J�ʠ$�h�_3V���W�h=�ݎ�`ξPK(�h�Z=Vޮ�����#����.L!�2����g�ƹ瞋�c��M�
��d�onW�/�	T	^�J�ܞ���7׏ŀS�EVBH��ï��WaM�V؁�vn�!{oB!�B���_mØ=i"��}z�Y��s�A�PQ*���]M���ĺ���F�S�L��wߍ�n����*!�2���G}4�9��Z3{,����nX;t���ܕ���H/��E-�"����(�r��m98��=]��}�P%��=����j;`��q��Qb���+тU4�	�Ġ�����Yg��=��7�|3�.]
B!��*++q���c�̙���h��#�ˮ��	T���0-s���hjWTF��R�ҊTY#ׅl.CW?E*B"e��K"��U��O���>���6!�̙>�=����\� �B!��^Z
�\�~����^(�{���}�xMVZ���[�&w��X3�fPVqq1�����X�`:;;A!���GEE�T;<蠃bZ;Lֺb�s�5C��a4����v���ٚ�ݡ��.��-�����wB���0�r{�q��{�_����	+��W,Q�\�B�`�� �b���B�'�y�n��nx������駟��!���L�>]�&N�U�v;Y*�}�2�k����M�VZ��4"UzF�����NB"gI������㯧�(��>']�7|��
$����=m&�8P�zp�}��B!�2zx�5s�ƣ�s��ܮ0����X(T`T3L�������]��5C�c�r�a�a��ɸ�����G��B!$y�6m�ϟ������
C96�u�X�ۥE���v����uC��^���\PZ��Z��OH2C�;!1`�	�km1fV���G�/�+T)�X����*�ocf�G�S������c�:��c�mk�*,,���G��^��[�r�JB!$���˓:�s�1��Ȱ� ���3��}�JqJ�O+LE��ndl�jlצ/�jd���q�`Ֆ!B���O�+���K
r�ܵ'��;^�+�Ǖ>&:�`�v��c�������7�kA!�B=S�Km����R�vuxJ&5Cy[�n�ً4hǇ���j���c�ӊ���|�7����a��X�������^����B!�$/999�7o�Ν;*j�v�#�����I�0Ts������
Z7T���v��_R�۲��9��wBb��A7��4�Ǻ�P�LK�dT7�"�,�!-��[�*^�����V�w�����m���.���kLf �B���w�]t���#�Bݎձv��ܮL_���]ܺBk)��t��SjK�C�&��	��L�Y��x`��{0���U��8�������`8��vB!�BF7���++�pX�}[��w�ݍ�v�Pt��j���]6��ռf(�21����a,��233� ��~�M7��o�!�B���v�MJm�v�mm[;L��b��v���$��d�}��ڡCSK,(��F>/8��#D�Đ��a|�^���y�,�7Y��w;�E�V���pe�� ��#������X+ǆ;��]VV�k����n��6ttt�B!�E��;�8)}A�0�E���X;�S����|��~k�H���FwS�J�4�b�M����j��	�%�L�"Q����BmE	������q����/���w�3Cs;!�B!��������م����0�#-GM����]��#�� �k���j���~{<��x���裏J�!�B쏨��8��3�^;�C�0�������bn׆c�kn���i�s���ݡ4�k�?���5Et��Ę����6�;�Y!�aIh��>㻩@�<"z�L�i�Ie0�L�
g_�Ɔ3W�m�|���i��p��7��?!�B��;�/�S�L���=�m;Tf�B�<�06�{����V��C���v�oh�`f�֦��,N��4��,H�����/�K
��{^��]�X�矾�8L�)3Cs;!�B!�E������\����4�wS]%`��j���&w1Ә &w�z��#��ŲF���8�!�G�4���B!ľ�/����ԩS��Vʱv٧W/�ܮ�!Z7�;+���`,Q;����[�Ǣ�As;!F��NHh�4���ZԻ���a/V�H�0��&�����oe"�L�`�}���2�A�]SS�;�o����N��B!6!++KJm?�3���7*�P�&B��M_���e�{l��C�"�6�AޖƔ4��e4�O��]����c���SP_5KWm��g�*����ڇ9W>�!�B!$u��v�+��T�Hj�!!j�����Տh�1ɺ��13�ۥfm�z�k����v��<���<��s��E!�� R��Ν����7(((`�0����~��e���ˊ��}H�خ���&�k�۳���QW9�\ �C�;!q�N�V7����s��:-- W!�bUzz��T$�`ev>�}��g�H�3220k�,L�<Y2���� �BH��y������첋�Z��H沫xejn"R�-A*�K�خ4�MmW
U^�*��o�R�"$��Ի#�n̟;�p��;�IK���ڇ�hn'IBq~n��,�+ʕ���߉z�B!��TCt�:c�f���Y�ñ�V�UIT־$s�%����)w~�l��n�brW>�x��Ý�h����\r	���~��X�t)!��x����?�{ｷ�m�z$s٩vhnn��:?���±�en7Km׮�I�%�㱮�	B�94�G�\=��k1�w�Ȗ��n0�g��j�{@���T��+�9ceV���e��Xm�����nÿ��/)�}Æ �BH������ܨ
J�n���x�W���ւZ����n&R��۝f� �J���P�7�d���	I$���=����/��}�O��v~�#��(/��Lm� mO�҈Ң<\p�+ �����z��uk���z9���bD�f'�+jј�L�$�:���:nD���]�UuC�P����a���ѬZ�?Z��k���4�|���$}�B!�G���t�I8����l;Y��f���v��a@�P'+Z�v���]el�C�4�Cq�?f�i��Ųͼ�#�
4�g>]������1�K�V��so�T�(	V�ڧ|N�������x�t�A�2e
,X ����@!���"�E���?;찃nA�.T4粋@e����nfl7��(�7�;u�z�vS��'T9�UV��[x�F���ɝ�v�l��f���2�����~sHj1fL�&��uM�3]x��)eI˚�=�¼l��Ǣbl!Č�7!}|��$-A �$a�
���$מ|5Ñ���
�Rv~V��S�5�h�#�&:�;}�t)���~ !�B�ǎ;�(�EQ`W�z$�ڥ���on�3��r����C&�v�C����%.�[�&�in'�*4�� >]���'6���u�M�k���n�{��d���9�y"�7s+���WUU�n�A���N��B!1"??��vN8�)�!��T���(P	��:�-�۵b��0���
�ܮ�^p�6��/.���;!L�'.?逸���v����$���љ�B+��U�c�%�b��@l�0�?}�q82A��Yx��ˤjB���vc�P�l����C���m�������Ё5C��D'�T�Z1�Gc[��z�!<���200 B!������c��g�a�����XϺ�|�cjn�t{V�����B���v��}(Hr����jk���1��n�梟b
�$�ڝ���&�nmS�K�ұ��D��L5����cx�5�<VE�p�鍵��$��b9���%����ƫ���:�B!���~����Css���h�b5֚@%�7���h�ܮ5���*M��+4s�R�����6��/.B��X��G�m<M�4��ddBY�*K@R����j{�����_/?G\�8z Į�+��?�?�^��X���q;oq~���8�m!$�Y7�1�0ah���bR+�خ�y����T�B�Ь�>�=�v^^~���Jz�m�݆o���B�.�=W��ϟ?;�3k�qاgnW�hn7����B�"2��u|����]X�� }��4��@�mwbFCе,`_D�n(4����z��4��x�O�%3�zY�J3^b�Oz�a��zl4�e��|����kp�Aa��駟@!���)--řg��#�<R��_"ŨH�cul<�P[��Q����>��us�J����ʪ�<��ؚx��in'��4g�$KZ�������~1�p̔��x��_c�Oah争�RR��g�>'��>��򘟯j\���ɍU ��p�z���(�o�/���ڵHV���]><X��^��\3�[Z{��v�	��?�q)ͽ���B����"��HnO�����d1��5��p,X�ۍ��ۅ�]�v�1�7b1�턄�$����p`c#�ٛ�n"R���Y����S,	VдT$3�Ee"C�+�cO�(��`���>�:u*�y�<������!�B�#�ifϞ-��+++��(�Ĭ���MZ�[[�d��А3ts�7�!�l<�o����d@��ǌIì�m�s���y?����$�nC�{��'��!{o���L�1��܀��������HH���i|Q^6�~���.�Z�X1u���c0����1'!D�竇�gu���I�[g͌�t�Nc��f�u���F(F&��5�P�srr$}sƌR����B	��*�S��ߡ�����C;�
C��ݳ�nh���Z0�lj���1��܊y7�7`���6  ��IDATJ��		�	�o�9q`c�yY��Mn���/���(���p�*X)�aUL��(e��v��Ǔ���SO=ӦMÝwމ�>��B	ΤI�$q��?���E&�����*n%N�
?}A��hrWR.���%s{i^l�
�RB�}X�܇�B	dJ�x��dmG7���ǘ?w��9�'�}�f��Ի $^���p�uO�ֳ���BK�df�K�g�#.y�u�������������X���޴�?�6!Dar߻�c�D��a:֊�*��Rw�����5C��i��%�fI�/�5�h_�)677�;��;�#�W�ZB!�X���g�q;�0_�h�
��v��rl4���E�kP7ԫj��c��C2��[o�pHeno�'4�4�b�js�WM�pt�nr���{Py�B�
K��)yd�B� �*.ES�J���HD-����&,X� �����ΰa�	!�=���p�	'��OFnnn�bS���`|�T�
7}!���#VI��+�@e��n`n/(����p��N!d ޶wj�I]D��c����b�q8f6m��#�}B��[_-����õ���3�X>��;7ཻ���}��]���A�:18�OR��;����d!#ã�]�(?Y#ۓ�����8?'�ǿ�eN�����!���j'~>�[[U�[�*�����_��������҇W3��q=Z5?���Hk�b������>������E!�c���q�QGa޼y())a�0
cC�*���Fv��ݻn�������B����wy]��Z؈OV��NH���N��X�:�Y�pl
4��IKzFt�[!PI�[�8k:�P^$�Ņ*�]$�h�B'n_"�|�|����Mʊ	>��V���>��C��^{�{��k��&]�B!�����q�9�H_���9�%@E2W,�+S�
��J�����skfpw5��cn��J�КIs;!��QC]�X�e��.'n��wp���t�u�,����� $^l����z	o/n�mgj�5+#}�����$�����<��	!���݉iuM��V�ܭ���[���ļV��SZ���x��Q���=ܹ�n;�r�h�q��a��������o�?��[_&�BR��N;I��=���w�vL$�ўst����c9M�������_҈���?!рwBl�k-Ø%%�/�8c1B+Z��+!TɷR�;4��(�<I�O���k�m��/�W^^����Gq.\�����BH*SSS��O?=얂V��i;Vǆ;�����v=�ʸ�ఁ�]ahw�'0	UJA*0��/���vB!A�p�tdg�_��-/I���/w�4r}��h�r�sk�噎K9���~#�ɀc���$ux����ﶵx����c}%����e����k1!$�_�Č�F���w�5!M}0�y٭^q�ӽM���\�>Ǻf+#{4k�����5��SC�u�]�$���z
�<�z{{A!������v�Ν����QW+�n'�̮��3����R�͍����4aX.}s��~�W3T������D�WTIA^ku��m^�C+R�tS|���`�� '2x��y�!b[\�$��K*��VE-�c�L��{��-�c�=FъBHʑ�����>Z2��*bT4戗y=���!Pi�ĭQ[���a�J_�
����t�핒��9B!IDiQ�8�@��d�t�Ʈ^\��[���왇�"&��(s�o~���KBCnv&��㑰W<�O<��g �CۚNr�#���Cp܁Sa7��l���<ZVw�B����.L�oDږ6�1�X�z�[9�ʷ�-����� i��U3�EM�i�B#=�Sp��/�^}�UB!�Jzz::� �u�Y���N��a����)f�C�����v�`��n�N�+h(����Q҄win'$���N�M�g�0f6�����4�P+�?=���`��Ifٖ�ޡJb��>+���1�����f��/�9�h5{�l�ﾒ���g��.�!����~�퇳�>�m���mw�)���"PYI_0n-8���-]��А~{� s�V���/�Z��r��&�b'2������b�mk�:�r\θ�Y��؅)M�q܁�5�ۍ�N< �}�#Vo��:����~�g9n��,��d&�!I���9�}�͑�.BH$��܅i�M�71���z>m��������w�C2�ۨfI]/Qi�Ѫ)Z����W\q<�@<���X�d	!��TA�N�<Y��瞾��c̶�9�N۱:��<�ui`8��vhP7�3�w}4��&vC��Y(�^ ��V��-n�4�uhp'����m66 �����d-�|ӗo�+�j�J9��p�Lc𥹏,�ANfHK��1e"�Z�R>�h�R���!y��1eee�?>9�,X� _~�e�/HB!�Iss3�͛�3f��9db!FEc;
RᎵ$PE��hpv���AD*3s�Y{���	x�%��vBIB�L���]p�϶���4���- ����}�sI���de��?����z<��XҲ�=�E�z)�7����/���U�_���j�P�#L�:#�7n�,��B��ʺ�\3T��#15�h�c]#�G�����>�}����s��G��͛A!��fJKK�n&�s233cR���^;T��=�r�PYC��ܽ�C�]���X�Z�+�vh�e��Y��]؄�2JH,�����V���؈�nu*���^m��R�2�<�-����9���4�4i[�#0�A����(M�z�&�h��c!Z	v�a�w�}X�h��^�]��B�h 77W�N<�Di}4�Q�n��Xk���/��4��i/�W:/��������eG<GQ~�s-�ƂRϟKJ�t�&�����f��NGq~N��->�<��q�����~BH��d���n���e����!�A�
���V��W<�B�N�\�j��ܢf<��>5C���QS4#:@w�q�9s��������B!����̚5���oQYYV�ʘdގ�X�$�-_�PZ�=!����F&wW`�˿m�ܮ��,��Z؀�V��NH�����$��v�dr��n�nsI�ֻW7���V�U���P%3xE+��HwW]̈T �/���}E�dH^G�J�G����x�	<��3���!�������?��v����&N�s�]�H��*P	�#������ghw�TA*=�ʻ�SV����BI���q᱿��غ�o~��؅��M�A�|��J���5��C�|�����9t/�t�n(/ɏ��C.������ŏ��KB�%��vb���/��
xA2�u��B�;@�	�3������4w��X#���h�>�7F� }��K�/^̀B!��)S�ଳ��ԩS��x���1G��
���@� s�b1Jm�^7�1����������m�U�#����NHL����$A�ܧ�5!ߛ� V)D#��s�VhVn�v�/R��*�1I!RAn;�Hpcx�G���i��M,E�pE�P�H��>�p��S\\�s�=�gϖ�^y��"�BIv�m7)uA�
���l�]ŭh
TJ��5��/L	�H)X�)�P�Jb��`(R9�SZ�in'���g��.�Ӹ���AIAnHǮٴg��<z �.\��h�.��Ղxx�#�ɘ�HQ���w��BF��rb��zT,Ð�O�kfD�o|uBU����@s�R��#5�H�|��&´NQo�N;�x ���*z�!�^��BH2��Ѐ3�8t���h����u��.�B��*�jr�P�~hT7ԫw}���v|V��j�rJ��~(n�n�f5`�j��	�54��D��}j�P���i=(��b�Y��R�
8�/V�}ij}������E+9�Ay>Y�2�����F[�B(�U]]���Jv�ax�G�t�h����X�8NN�Z+�D۫D!R�E��D�ȟ��s��>�?�g���.H��^�[<�D��'���D���}����.ĩN8�P�����1v5��{l$U4��"���]���/([��ܲ:��Bs;!ɀxI:��=���
t��し?�Ʈ^ؙ}v��#��$��>�޿��w� �E$;��ۅ d4�����=��+A0r8����#A�!�W�\��.�1��L�/$��@k���U�T$����C�Z[3��ӭ�i�~�0���h��beZ�U�v[�9c�<��x��'���B!$(,,����O<���q3��sL*��A±t��w���p,�Sܧ���'Z���4���n�0�f5b�Z��	�4��d|�r��6����w�_o��֭	Vj�J��{.$�b�����a0mME�4��D�`�|���B���m��3��1����.���R:�ʕ+�bJ���M�D ��x��盨�gee%�܂D�����D�_�����^��s��߼x�~��|s<1��x<���RI��3g���X�SV�$Z�J�\���*�G�֤��/(�*�"���@edr�(��[@In�7'��o���w�}Y��̎%9���_a��ɐ_R�0�����r)H�Ѻ��7n�[��ɍU ����u�7�kA!�����C�j@�s����EY7���U��݊���f���*g�X3�GGҫ��i�Q3�R�-AXVj�� xꩧ����L�-���+jW�$�痃�䰚x��?{�3?�D���'����Z<w��E<���{A�~����u;���ӭ�wF�T��?�C9'�t���,����G�/s$c�P��Hh�����6�{n����Pp�{��ݻ.X�Ո��NHܠ���$D��w߄	C�U�ҍbݳjlt�]D�/VYi=��If�"8Q� ;D+�,\)��^��+J�A�Jt��1Vƈ��������^���7oF$����d"H��X�|ip�/�evM��^~�I�}"����a*~�@	����>��g/��"=H�,//��8eeL�ŧXoG��`���=4�J-N	ûn��N{AS��������ڒ��:;7�W���yٸ��_a��-�������p�/&���L����)�u��}�#����2|x�� �B!��uC��G��ro��[U+T�b���
��|G�w����Y�P�'��=�v1:>5C�eY}<��a���Ə��.��f����ߏ�?�8j�����v]K��e����)�$U�"�Yև��g�= �ά�w�&K#�F9L� !� Eƀ ��c��:,go���y��ߵ�������%$`�D"#,��Q�a$MN=�߼��vWUߪ�U]�]=s��ݷ�	i��3���|����y�ݞ�����y�3���gϐ���>������_,������Ax|:sƲw�tΘG�b1�#4y�#��nޡ�34�cY���;>�y�v�v~ΟG[im@�����; 
ou20u.5%v$+y�A�"�X�Tҝ�m��9)R�����u�,�m��73�w)Zeb�xNX���)̦� (AJg	�-[F�\r	��������^   cٺp�m�QSS�˕8�3'j�V.�e��!P�50��w��v�H�s�&4ӳ���C"  ���K\��'��|Lrc�u�vSTش��:{���     ��~� ��ϡ��v	�C`	�'�&Gf��ͻ?'���=y����A����y]x�a�`����Us.\(v�~���?��?hÆ   ��w�!��}��������w�;�xoi����^}C�b��w�����v>JJK��,z� �� ��9|  m����I�����ɭP� ������1yS!�'+�Pb�z0-TY�i�j�AtO#�*"�؊0w�����k����ٮq�4i}��n����>tO��   @��}�٢u�N��D~�E]�
��_�*mp�T�w}�*njl�cj�h_07/�ĩ�p�lo7T|���fzak�v�   0����I�vPT��o����_�B     �0hm��������V脡��%���td'���I��ŗg���I{�|}����u6��WO0�׺��5����Yg�E��v=�������v��E   @.ijj��~����}H�d��5��^�]��:����ڵ�����w|v�+v|��>�+��׻���vx� ��(p6�Q���tZ�>�7ni$+rnb0�d$�96��P%5�D�}�A	�ԸݭM�i�J^'W"T.�������|={�l��W�B�^{���x�	q�   	�9�S�8�x��y����Zwl,�߃Z�j]V�r��4�+�TT�D�T5��!P  �-��������"�    Phl;����t�����c��(n'�&��ٲ'��a%y� <C�.�#���ǌZaP�aО`<�0甕����_OW\q=���b�{�   &t��7Ӳe˨��"0_0�9Q�ú��;�� ��o���<CS1������v|������}
��w@�@��Q���!�M���ۨ��;%X%��av��!Zɛ�&��@��"��L
W��Ny���=����+�����R���wz����sM�st�͟?�����n��F��/~A�>��B�   �s���-��B�^z��g��8�gM�_;�˵@e�䶂CC���N������-%ʹ~v�  �{^۰���Koo#     Px���g�&�ES�Po��.A6���)�n��M����̕����9:�Q�UUU	�pɒ%��ϰ���   � ?~<�p����|�&L��w��n�{�����af!�|��o��cs{�;4z��r�ʚZzz�D:܋�O �	� �t���d����1V)�Jf7�&�*�,����0r��̐le0�K�DU�7!B�*2l=(E+qXW��������.�慠)]��N��~���v�Z��L���
   ~�3g��_s�5TZZ�wqJgN�Z�s��vkc;#�(�@��w�*0�jD�ri_�in磤��6΢�n  ������{;�o F�     �{��؞	t���j?dnq���v^��1lϐ�BR�M�!?����F�#�u�=�:�aÏ}�ct�W����/���   ������.]*v|�2e�oP5�+��Ϛ(z������z����_�{�v��q�o8��n	���]��k�O�G��Rw�  � ��#�CB��|V1u9l�SJ�J>U50XĪ���!-z��B���Zd3C�փ2�n�I�*�<�>�G)X?�lD"���l_�~|~��w��{ٍ�|�������{�9��OJ6l���   @&�u�������@5nܸ��t��:��c���N���!���d�}H��])R�)���Jz�s*���ւ   ���Z�yE���!��7ѥ�M     ���HЃ;�i���>|`���4�[��v�aJ)@��f^�������x�f��J����/H�/�{��v���ɓ鮻�%&����C��	   ��7����3g�1?���XT��^��*�
���C��v�b,�ops{��zzh[5�ǐy 
 ��(CV�j��R�j۟��V�
2���Sc�g��'�V����I�����dн(��`k�OZ�J�v���֚0��q����O/��"��g?�u��!�   ��1{�l�馛��k�����@�(�X!X������}����a7���ڕ������z�P=�F�  @nx�͍t�9Ǚƾ}�s�o��u��t��TY^�{o�j�@# ��8oQ3͙RGQb�C�f�V �0���RA�4O�����&w2��Dꂬ�3�w�Щ�]��m(V5�g�ce���Rϗ��u����0�����вe�D��w�����    '�/������[o���F1���w�Cw��z�hl���5�����lo��<�V���PT[ � �0
J��M�tM��n�m
��T%�Pe|�jeQ�L�r��$�M����:螺�H��i�A���U���pu�Ma�v�x���y���:��9�C�/���~�󟋠;   �_#�ΝK7�|�خ��l�Y��5�
Pn������@e#N�TZ��#�P,��j^�k_0	S���	u������?D   @���V�c��c���������HQ孍������+7PmU9m�w�n�?��vw0�9�q*M�PM;��-{Qԩ_E���{�W6l�� H>����'ŷcye�s�p �X|�sΦ2�z�,�;�CY�e���X�q7�0l'��ar�������E�]��q�b7�c9{�E�|�a>��r�!z��ͺ��&���{EPq���j�*4�  Ȁ��%K��-��B---b,߾`PsF�wh�����s�oh��5�C'��T��볭wh�۳�p{�,Z�ZL�� D���]�ZJ�7�۶'GD*�p�jb�he0�V	�h%稄��he�g44(�����71�д�w(���Vˏ]�ȁ�����f������;�<Z�f�򗿤�k�  ��	�o��F�=m.��\�S~�D��^P<3���sq�8�"LǍ�v{��lO70��TN��,P�Ll���WR�  �c�b�ﮠ{Z+��쥨���ʹ����մ�`;�	�n��t���.����{�8���7���u��S�`-��>@_��TWS!ƞ|�}��?�W�Г��b���3	  �:�Y������H�m��~��K�Р�94�{����ӵ�G�;4x�F���Xv���K�Я��տ+������P�j�������u�]G��կ��#   ��B.��b���F1��`�ε�~��wh�[�錾��;��u�۝��<ϩ��*Z��|��&Z�Z Qw F9��]��Ltds�&�(S�R�V��ɌS�h�67����i�J�I����U
s#CR�J�ܓcىPQ��%Z鼷�:�1>�>�l�����/ӏ�c��nC  �ZX��馛�ꫯ[�#خ�J�=�kxy�tNjw�┎@e�[��*_[*Ī��3iek)�  �7�KО�N*$�z�F?��L_���Th������T���������ڻ�(J�������7�]���诮]L���c�;���6   �Yݚ�����l�}CRܭ�!ix�:�?z�1�^�lpWy�EER�J�9cY_g�	F�S�:ǯ���8o�<�������鷿�-�X���  0����GߛP�=@��F�Wh}���˱����ή�z�X����/�-�R��|�&z�;VUp`����9���{���@f+CJp"��A�2��^Z����ײ����V�sqV�J�L���32��GΊ�وJ~B���^�/�k�9'�1>�:�,:��3E����^z�   �>�s��hٲeB�*---�`{Ps��:}&^�
��"N��)՘]��N�J��kn-�jl7�/�7��/ �    �b��zR��Ҭ�	4i|U���6NQ�7M�D`lû �  j��2Dg�n�����34�ۍ�!Q�6d|n
�+<Ñ+����*�X���<��3$ˎ�F���'�+O��5��	r��؜9s�_�"]������GA�  � ����[n_�(��~׍f��)Ԟ<���y����\|Cǀ�����%�����fzc�  �� �^���6SmA��Dj���<%@����S[�O+�w��aE\sD��&�p��z�~��ԫ"u3C�!� '?"QP�R�B�1t��O�=����裏&o   4�9���N�k����;�<�<*�v�X���A\#8��x�'���s7qJG�rk^H���*׭!w�n��fz�5F      ���go8�>q�  ��Wv��MtL�.�����к�gH��a"Q�k�g#�/,J��l��EZ��]���#�u�=h0bcc#}��_��n��~��ϰ���   �.jkki�ҥ�kƌbl4��:s��Z_;y��\��7�;?���*��Z�e���ȣ]���7䣤����E��BN	����; c���ґ�YtZ�~���5܍7qJ�:�$yc�z0}SSb�ҍd�~FJ�ۇojR�U����|�%�+y�ea��γ}m}��~�����ur=v�	'����Z�z5-_��zzz  @a������t�u��駟�2�������?A^+_��\�v
�[��T�J����ۍ"U`�B�b�U4��m�     0�Yz�B��_@   �y�@���f�i5���������#�x�5�=C�|�ݟ3�C�Gv}&C؝�B�%ړ�s��)f�����
cl֬Y�/|�>�я��;��$   �͔)S��o�����&MJ��`��u��;T�3�C�o�j�R���-�X�;>;�+*+�厩���! � � �1v����xZ;uwq��Ū��e��ܭaw�ΐ�TXE�l�g���� ��a��r�|�555�=��C7�|3=��Ct�����Ç	  @�)//�+������Z:��c�X6����B�G]�J�s�W����~�(NY����S����]C��mmW�Uee��nl6���      �v�m�J�v�U�qf��.���?���~�'���  @�Iz�S��iG���=p�34�cI_(��=��S�}���g����g��!:
�aT=�l�e;���@w�y��~�a��ر�   ���"�~�UWQUUUV�`�cA�mޡS�=y^�7t�݊���3��*�P{�gEȽ�v<=�"�E��Bw � G���Ȯ	t��R�:r�F�J���xe�S*�N)��T٭��f�V�I���i�A��nYEFK���������#X�R�]5�?�����b�
q�۷�   D�	&Q�n�:L.��|��s!Fe{k�]>f
T��q�0e��D)�9c�]%R%�)s��1�n'P�D*Ŗ�����*z�H��D�     ��NmU9���7PUE���/���y��   $a���i��q�uhr��7$����3���3�2����C�Zʱ�~�zh�&v�a.C����jkkEȝw}��'���w�y�   D��`�����˨��,R�v�X>��w(����*�����C��5}Cۀ�C1��� �Ll���WR_,N ��w �(��qz`K-m�I�m;m�t���|������	?;��,\��˸��5�.���f�$R�yUD��E�ǠE�\�XaΉ�X]]�q�t뭷�3�<C<� ���   �̜9S�Y��;��`�j,jV>-��faJ-R)�)�ւ:"�N�BR�ro_�����G��:zb�x��G#"      c���+�y�$�y�~�����   31�������Ӷ��3t
�KR���g�����Aw;�aw�_h��#��W?/�к��z�`��A�_��rQJ��������^˘   ���ŋ�ݞ�;�<*r�Z\H�v��F�wh*Ĳx�N��V����w}6��ߐ�Y�BU���;�p{U�lZ�ZBC�� ��@��1�P�H|�PK#ڪ����2%L�+kK�5�lq7^S��.�S����T�LR�"�6���D+�"��5�uL%2�r���%K�Х�^*�U�V��;ߠ  ���~:-]��.��@��-Dq�Ϛ0-'a*y^j��UN�v>�l�[
�k_��ZP!R�L�NnG�C�      ܶ��t��6�<H�ߏ   5�>�ZJW�k��6�gHd���8���-��7���z�V���g�hqWy���#�a���l�??����(�ڭa;�8����$�ׯ��+W�O<A}}}   ?TUU��_N�\s�hng����sN>����5���;T��nޡN1V,������n�n�a,6H����r��� � �M	:sv��n?��'��S�!�Zc��(X���N��aڂP�ߥY��7m����KA�Ma�ڝB�ټ��5��p%[�n��~�V�^M�ʘ   ���8����)��"����]��`�Μ\�Q��n�c�t�)�XR����3�4��{j_P�T|��~-oM�^      ����4��n��u^�@�>����7@   �y�5A��i���-40���<Ì��P<��X$�d!�9�.w�6����BU���3�B*�>Z<� �������ԧ>%B���oh���   7L�:U�q�u������X!�Uc��+��V{�f1n�u���q��^��?���]�q��;��ή�za
4(dp ^��c�4����;ykcp
��JK���%
��Ķ��vO�SE�-M��H�F^#H�)**�T��xcc#}�3���o�]��W�X!B�� @0444�UW]%�S��2w������U�Xe+LY���T"�5؞l_��T��*q�Q�2�T�D��k���VT   
�����Ʃ"l��{;	  �7�JK�??-U�s�����Oһ��   =����6S3�Hz��pWd|�η��l���ܭޡq��/d�*���'�n���D"rO�n{�WO.J�v?~�)S��[o�o���z�)���M���B  ���?\č��!VTT��Us�ձ���wh���<{�n��V1��o�۳�oh�K�JiSb6��}�  �� ��ҡ�t��6����Z�"�p���Y�R53$��m?(�*�-�t�!L�VA	LaP��r%<e�����n��f�馛��_��{LX,�  �n=��E�a
S^�FQ�ҙ�����I�J��)��v���8e����8e��l�)�p��H�Uk|.�y;��   
�������A�3&�����3��/   }n[r
-l��:��76�O�:  ���}�tx�L:}����I{~�9N�k�Y��靟e���oh�Sa��P�ݓX�B3~<à<E?��Y��:Q�2��lִ9t��믋b��~!  ��q���/�=�z�b�P}B�1x�f�P����!�Zۭ���?h����U�5��p=��D��� �  {;���މtUcu����lE+"�5f��i�A;�*%TY[��J���>��I�6ZR�
S�
S����uY�\�x�8>��O��O?M+W��;v   g&L�@K�,�q�'Ƽ�Mv�Q��$`}�0e0���m��*�����!�ւv�v-����^j�B�;n  P8����ޒ
�3��i˞C�z�  �GC]��=m�t��"��  @���Ct�w2]>������Nޡ�7�ls�b��w(���Gq<.�T9��7Lb���~<�|�ؽ�w���-�q>N;�4q�ٳ��x�	Z�j�B  ���3�Ȼ=�s�v�uQ����LQu�����C�b,�p{zh�2,7�06|���L�L��UM��C  � Ƞ?�����ʖ94pp��V���`e�KLAw���20f�*-V%��Fa+��z�D+�s�\�6�w���Κ5���/��n��z饗D�}͚5�&  @�c�9Fl!�����Z1�Ka���(�S:s������Eu�=S�r�V�)Ԯ�gn-��������^[WO���~��  j*�9S2Ư9�8�  @��	�����C=  �?]qz`s]�2�znOjM���k1i�0����[܍c�~!#�B5~<�0<E�9^��(����O�N��v�������W^y~!  8PZZJg�u���.���21�����Q��|y�V��8�W�e��y;�0�p{U�,Z�ZJC	��; @၀; @I"QD�[�>��B�G�؋O��͏b,� �s�`e�~�M�������)�ȩ�A"����:S!���&�bQ>�'��ݮ��l�{��ضm=�����Sww7 �X�ۮyA��~��b,�n<�"V��)?k�U�0e��[
f�U6��q��������F06"R��)�Hen�BԠ]�}D�z@Tq   
���U����$   ��������J   �g(QD�Z�.in�����mX]q������r#���\�%���B��;���.?^��:�zN��t�]cܸqt�E�c����/|�G���   �ĉE)MMMbl,���c�
�g{m��a�g�P�w��s�o��}�ۥ��RbR��'�^ &� yjs�N��Ds����xK���<4�,u��x�$�`E���lg�؉V2�.Ī�J-T�E���E�ms�2'�u~�������s�ҧ?�i���?N�>�,=��S��/���  0��υ��~饗
a���.5n7_w|4�X�d����B�,C���P�U����Z۝�\[��T�*R���,tQ=*   ���	������4i|��   w��XC   �����贙-4�k�3��z9�^a���K��n��_h���8l��{~.�5+|.�к1�9Qs���������|���Nz�'D1�믿.tO  k��R.���~�������?/׈�X���(x��1c1V����ש��v�B,�%���Ụ��	 0:A� �ʺ=1:2q}�z���P*��pã����JK3�d����`'Z��܇�;v/2������z�7�:�S�!���B��������E���;v���{z��h˖-�  �Δ)S�K.��8��!4y����KQ+�k8	S��N[
�(�P�s��lav�m���#���)o�77�   (d�j*m�-�;�֬�J   �cp�{�8�>  ��vRӤ���r/����>����>�C���'hW�%}C�?(��I0��d%���3$�5��������;������A�׽\�����.]*���Vv���~G{��!  ����3fВ%K��.?�#���g;�+�P5^a���F�ޡͮ�:�X:�X;>��~�r�gKН�9��o:m:�p; �� Zl;����lvuڟb��˛���2׹���d�����*PYǄXemf��������@U�U�!�0�|�ڽ�QAW:�gϦ;n��vZ�~������A  P���Wn[��+�.�ն�xԃ�(	XN�HR���{5'aJ�C�vBU��v��{EU��5�v�G�  @�3������Ʃ�    �ȳ�P�ګ���tPg����d������N~�[����Tv7�c�1�1r؝�,Y
Y���vS�m�ٮ�2Gw�Ϻl�7��:�����'>�	Z�f��
��y���#  -p���Σ�.���>�l�'2��f�>�~b.�����C9�����<�ۭ;@�c����S{k�p/�C F;� ���ӊ��te�l��,8��W� ��Y�<�I
T雰�p%�(5�N�b�0ejrigP7��U��]���u6k���y�\�97�q~<��q�]wѓO>)ī��zK�4 @���c,��/�X�-ps����t-��|�X����z�S�=}^ue��n��`��ĩt�=f��ۥX�p���J�l����!   FU�e��o�N      �z����j����znW������]����m��r,�]�=�/�mr7{�d)ʒב�e/4���{{}P����'G����z�~�a���,�� @�a��k��ɩq���/��;�C�B,Sk��7t�[��:����3i��R��k4 c� ����V��9���{������F�op4*���&*砻Q�RWv�r,�����vc3C�HeE%Z!b=G���՘����������Z�v������O�S�  �7����/��-Z$Ƃ
�5�`�j,J��k�Y��R"���$Ly����H��Ӑf�=%N)ĪXl�J��ҊM�qC�  0z()��1�㛧      ��P��V�]��L��[\u);���?4z��6�d�=��j�z�ZM�#�w+<5m�ks�cQ��|�^�r�>��'���_/�6�b,�<� i��شi�D�����Ɲք5�O���B��\#�:x��J���]�����w�
����l��=ao]3=ފR, �� |��5M�K'U�����͏!��'�nlp7
W���t�]�Π��Aw��3�U�v��@%���Gy��U�ʇ ��P��`�G���~��1��9s&�|�ʹl�2z�����_֖-[ ^ �F}}=�s�9"�~�g��B�Ϛl�%/׈�X��)�9VAʩyAi~��M�����TZ��ǘ!��=�n���5|�}Z[�<z�u����   �H���na�gM�ڪr���'      
�g�т�f:�tw�+C�r	�Km*���BØ�U����|B����0�r#hJ�S{����a���<���˧7�e��k�^�x��c��=��Co��&=��s���SGG�B @d��a�=ĳ�>[|-e��5��`|Pa����Q���X�R,��c���J?�l\��g��[	 0�@� ��-�c��g2]1��:H��(��q����Z%%z!w;�J�7~F�ʮ�A#O5�J��9�\�k���ݵ��裏���.��~�iq:t�t�{��Ӹ=f.�luuu�Ķq��Q��?s��(���F���|�ٳx¿�|mߙ��;������������O�o�*_a�׃/İ{P��䣝H�y���v��v�@5����@e��.���*Z�;�6�@  `t��7`{�����>��{�]     ��x�@��UM����Sw���F%�C�;?'�ڗ[�]b�	�x�~���&�>���\�e�Kyi�%��.���������;�T�=�����g��uz>��nz��W�g����z������ �.���"����̻�3Q��S�Z���;��z�r<��w(��Cc��T�e��<��3<C�)��'�s&ҁnx� �Ep dEw��\EW�̢����7G�J��~�C63��gW�b�*��t7�U���
T4r6�6w�5^��W>ǂ��͸�5���x���O�^~�ez���u��aG��^�����G��?����
l���@���5&_���������H}S�/��{�s,,����Z�?���Yg�E^xa�$����)*�|�q
���;4/$��n�v�p���=����IS�U�5���   @�t�8o��OO��H��j     �z�j[-]�\C�������n1V���*Ŋ��ܝB��]�����5׵��B�ϊ�ڝ�#$E��|�����P{�A� ���]�iMUU�(�������z͚5�7d�T�竜)�A�~�3�?�|�3���U����Οk�j1Vex|�N8A4�_|�Ţ��ɧ8�<�\��������X�;>�l<CyTO�In.��8�R �*� �fh�&���bZ<��&�lARS+C�x���7X�6w'���8���t�D���e���Tm�f�ʊ�+��8�m=ʂT>��l�u������#_�җh�ڵB�⦆ݻw  x���8��y%ۦ�s���0��X.,�%�e�T^[۝�)�p{����оP9y��T<|_�q   ��:�r��)�w������	     �B#'Z�ZD�47S���~�g��j<�*�A�r,�������^�v���3����:?c~�������:��p�>�!q�ݻ��{�9Q����;����)���D����a���;��r*��LA��ۛ��;��?{��>����$dS{CC���a�<�B��TF��?��;{�<G`��ҥX�ޡ�g����5���0�A� k����sia�^���$������p|���$b��4�����I��4��a'X���w�-�XP��(����
N�B��@�t�E(�-�]w�Eo���hk���@;w�$  ����^����nk��&hQ�������cVa�(X�ϻ4/$���*�慴Penmw�L��������k[���9� !  dä�U5��W�8��:�W�AX���Y�J      "��<D�4����"L��z��9nis����_�|m��|n*�2�m��G9�o�=L0j��h��O�N˖-������W_aw���3 �0�P��'�L�w��O�:U���#��&����B�{�}���&c�`��R���+<C�+����f�IooŎ�  � ����)�BKf�Pס�����A������,Z�O�f�3�-�w'�*����@2�>��n
���X�*3��t��1��~��;��~�ɟ�惷%\�n���ք� ����?O,^�8���P��5a�[A[Q��E(�,C�r:T[;;�S:�vlE�240TU��+�� * @�|��K����V>�v�?�=������8���dO[���8���v�*����t�gD���     �"���5���ɇ���H�+4iZ���ӥX��{�d�Wt����N^a��,��������_��l�u����9�^y��8|������A�= ]xw��;�Ǻ�:1�0��(�Uc�����=T���P�4�b���w����G��I������� �w @�t��i��
������l��,��U�=����.�IQ*y#�����Nb�Q�2�U�Fw�6�4a�V:׉�Xs��?.Z�H��smٲE�����khk `�_W�9���Ρ��N:)��'���ӹB��Y��u���A�.���J�R�S���N��T�v?���=C��<��:��b�  �����64\VZB?��5�PWC?Z�
勪�2��/^�nw����ᯩ��'�{w/u�7yB5��篥��%ű�	     (L�uѪ��tes���4k]
�0ᢁ��ܭ-�	�Prw
��С͝F��$��}�{�s�c�����xPk��'M�DW]u�8:;;EН��_y�:x�r- `l�;=s����N����Z1���������Y�K����\���s�c�����z��:�v�p��7Lۇ���Xv>��nϩs�AW?��D4��  Hp ���7�i�&:�t7��o�4�����%螾Y��G��C�NbU�1�>����^T�׋�h�� �5��sMMM���멽�]���x��h�޽� ETUU	1�SN���ٳS���ӝ��S�
K�ʅ�%q�\�t��	T���t�=)B9�Ucn߳Ml��C  A��@;]������V�X[�q������/��S�D�8���o��~�w���cf��yfm+}��W����::oQ]{�q���H_��<����#      
�X�hUk1-��L�z�S����_h�o)K�F��3wv
���B��Z���Q���6w�o�v�r�����_�ܰƃ^c=?~�x������Z�[o�Eo��(�z���0�������;<��Sš�ӳ����ڽ�G)خ˕�h�/�2<D]�0p��l�Z����Q<|_v���^iE)  � ���FM��#m�&v�f'�*�6W���������GnO���*�`e���n���hejN�Ƃ��x>��b^x�8>���Ѻu����_ֻ�+�� 
)H�y�"�Ώ�snk��/�*j"V���U���ۍ�Jv���bU��M������������;�Z� � ������k��;s�N�����]E����N�H�����2��v��o��os�1����|�N�?���Or���ϡ����H      2k��h��9t��6���P��R�~n��sFx+tO$��ݟ�~�])�|�� c}-�B�6w/^�D��F�-~aP^��<�Z�(��O}�S�m�6Z�v-���˴f���(�������>��o��3Π���>��:�+�p4�ݳ��S��m�g�`{Bx��p��wK���`���V�UYSK�v������ jp �N[O��o��+Z�i�m[��ʦ�����xOV#��F,}Cg���Tb��R��8�-f����읂��T��_�)(�*�k�\���������M-b���'?I������녀�s�N�z @~�mO:�$:�䓅0�`��@)��$X����`���5Ԯ�|T�ܩqA
SI�*�nn��SB���o-�
��s5�]U�яp;  \tB�W����>���u����4&���h�j�9O�m��!�>����O|�z�[�SYi��<�~��k��/�7m�{�      (dvw���:������2���XV��i�紦��W����X	C9����F��X�%B��0}�j���zr�`�B�^<�(��Aڭ���y~lllǵ�^K���"��ꫯ�cϞ=�
(��3��,wz�R,޽�x�i�۵�<��UO��D�0{����+���+4�=�T���z�LZ����� �A� ��"z���3����v0�M�6��6���4�`�lv����N!��V'��]�2�V�`D+�X����B��r-D��g�vڴit�e�����Ɔ?����/P{{; r��F9��cE���N���]�q���s٬3��x�D�0�)��$R)����TV�ʮy!S�J�S1�s�F�*����� PRI}#-oM��  p�����%��G���Y�5�#߼��������|��v4���Rey�����6�6�������]�8����~�՛�/��:C��      ¦?��K���f*��F���T���چ�-~aiJKK��l�:����Z��C�(}� ݥ���F)���ot��;������z��Z�^r�%��y���b7h>x7莎���o���Zb���X�w�)������F=خ˥w�
���ܼC�p��w��	:��v�_��B����! �� 9�]��{�lZ\�F]���6C��I�rmf�d;��Xelg�[�����G�ж �㪱 �\	Oa	Wٌ�Fu��Z����ؘnl�y뭷��7��wny��G��0�1Gu���?�xѴ0a��0)��A�R~��R��27jaw��$�D*�}�O��^�����TR���n-�$T95��ظ�2�V�H�[	  r��[�C�G�i�Ǿ}����ц��}��$�Χ�����n̏V�Bg;�.;��y�gM��߽����rq�      @����!j��H�*�QoOOJ��BU1�S�=c��%��~�gy���·�$+	?&�K���Q��	����͸���u��y~�?�8���z�����;"��~!7��+ w��0K����X�>��w�P�jf��J���;T�ٝ�C�b���;4������>bEe��J�A 聀;  ����v�ч�k�����U���VN�����[R�R�3X�4ދ�ܭ�u� Lb'V�q
�) u��ׇ5���ds��Z��������O�tg!K�{zz ��w�_[,X@'�x"-\��-ZDS�L1�ѹNX�s%Xy�VX�V�D�`���WW���0
U:���im��V�*B9�/8�c�T3����SC�{n �����I���}�r��o����� �_����]�� =�������q��-�7~�     0�t(F��hɬ�lۧU��S��\#}��a�����0����������?�ҬD�����w�=Ho�mn��:�ֹlϏ7Nj����[������+�П��g����{B� m9��E;;�b�z�TWW�:�?�v>��aB�Q�[ǒ��o����om7z��z�N;>�Q[?��QA](| x w @^JЪ���-4sh�h��ݭ���X��i3�3E+�6wsC�J��υ`���he�E+�^��^ǂ�r�>�qݏ'�s^��9o��m��{�8���>v�����oБ#G �	��ܮ��v�N9�jhhH�"Ю3'���ӹ(S^�FU�"�[
�*�p�}k{�,L�B��ւvq�V�y����&Z�iH܋ @��	���ہ����w��|��W�;ν���i۾���O�E      �:��|S]��L��[3�Es�
嘲��R����7�osOͱ��y�c��w	?U�?&d@^��q\5� {���B������4i]v�e�`<H6lHy�z����_: @
��͛��a�0<�(��a��a]#*c:ޡ|t��!v;���ώ��P{Vޡ�3��"�_��&Z�ʾ!�C �7p �7v�h[�L�`Jui������Ūx�/v���������U���t�J�݋��p����习��̩��?9��?8­�7n�w�}W�X;v쀈��'����������4G�Z�:U�*
!�(�S��,N97/�m+����.NŅ�}����A��
VUц�i�n+��{�� �0�R���77�Ǿ�[��A����?XM?���2�7��rj��F���� ��~   ����-C�2��U���n۠�]���X´t<���p��۷��s'�P�ڶ�����K���9�����1��~��;��:�����B��X�4ݹ �=C.� ��?hg�����C<�3����\'�9�����c<�>���;��B��s��=�y�	G�P�3b�,~�7�P����#��;|�o*�ߊ�v �?p ��C�|k-i��ءm��vyC6�XVVf+V%_������ܓ�U�A�*6�uC�P��h�$S���$Z���B��>��1��s^�5���\�D9r�޽{E�}ӦMb�µk׊�w���h����	nV�����:��ϟ/�k�q�������~<�"�~�]�j+R��m���F�Jݼ`mn7�T:�
�]k��
N�N��^N��  Q$
!w�ہ�����o�@_\v��qe%�󿽉.��Oh��C@.��'/��xǁ(p畧��s    ��M�b�����h�@=vfcY�2�`��?LXK�F|Ä�3T�b�}Cݐ;?:��<|��i$=D�G��̧����|��s����9��Yg�%���W���rA�cmݺ>!3�3f�@;{��%.Z�����Lst�����?��'�͘��wȸ�����q��[۝��=x��b,CȽf�tzt[�"� �� �H�H�c�q:~j3�+�E�}��m�f�k[�ʦ����`���n��vB�HXnr����c2+�/�t ^���8�����^G~�>}�t����c�"�Y,d�����5�+��*477�;�*��p�B����(���DA��&a��ܨ�Svw7�ʋ@�l��1�P�Y�r��乢�"��B���|�  D�|��n�|�7���&�ҳ:��ÿ��e����)��# ��o��p<��f������:z(_p���n������m��8   
��X�Vn,�s����m4�~��k�p*�2y��R����&=���Z}ô?ȸ����������%c�G!�����5t��e���ds͠��ͱ���q7h^��X��G�m�z��E�B���s!�1�C'�|2͝;Wڛ��R���<��e;'�P���\����Gu���g�ޡ����;��ͭ��v�����<D�w8�G�S'��8 @6 � ������i�dv/u�kl��)�*���]���(XI!J�s�tD+��&Ib��|�ڽL~E'/�����:�y�9~�q8���������l�B�7o�;v��u�����!f��!E(�X��@;?�P{]]]�\�k5o�V���̍�8e��bT�Y�2ۍ��@�C�k�K�Bu�xz����mC� P8�#�p;��G|��WS��z:�i��\����7��_�_�Y�����H��k���;^y���3���Aˆ���c� ޽�w_MW�c� �y��z�    P���=F�&̡3�SW��b���_��&d)�˧�܍���oh�
U��/t��9y��1ae"�3A�~^����E��нNkt��g��|6s����,�:�����`���;���*�BY���� D��������(�S����z��s���X5�0W>�j<�P>�O�v�v7��/��=��l��ޡN{�kk{�Dz�`�9� � "Gg������M�Tܱ����f��rÖ�ق��<1"Z鵹;ݽ�ܭm�#��X%1��j�V���:�s^�g3'�y��բ�	��m�6����w�߾}�8@Pȿ�3g���|p��[ZZ���B9�˵���*w���
��G��a��0%���mE*�Pe��┍0elc��<��\D�8 ��C�ܗ�#4i|�ɓol�ۿ�p;�FOߠ���'��N��q�A�sNh�o}�
��& �e(���|�A��.�>w�DZ����-_���mړ������~�77�Y��Α��w"x   �v�Ѫ��ty�x8�ͶKu8�-d�]���cx�����KPU�e�j��l8�X�i/1��{>`X���|�lר�yY���9v�sهY�h�8$��c�ΝbWhnzokk�� �5'NeX��3�+r��w)0�7�;/�/��Q�úF�>cvޡ������;�ʰ��v����C�_��;7y.�ܔ���p @p � �,On��I���� �tv�������F��N�2�2�#���9�n݂�)��[����d��3E*+A�VA�97�q����9?烜���e.�d;���0�mooA�]�v��w��k~�o|� ��f͚�
��s>i��ɦ��|��j^�
V�
�{/�`���^�����N�]'�Ώ�!s[�J�r���i+A�0ŏ|��V�H��  2����?�ӎ��{Ć?g�����ϩ�w��;Bw~����[����>�O��v��~� ���{C]5=�n��{9=��5�iڤZ���?L���A�   ���D��o9N��B�b;D���b,���Z�&ݓ~���ݝB�����ih-];�%&�j3��{e;��sA��fN6�x�]ٌ-aM��A.ǒ!�7m�D}}}@�������T���#��C~��GM�h���	�Y���_3��# ��lwkm7���7�v�ͥ�Z�ћ�  n � �4��h{�$��i��ṑ�N��7��F���Ħ�At7
TR���
W��+����t�=
A���1�e��9����|�s��e;�_�Oǟ|���0���!�����~!l�s~<p� ��c�{2a��3g͞=[ls��]��?01i�$-�@�}������y<��v�/q�I�򶥠�0�(PY�t��s[�ʰ�`m�4zrW%�C� 0:xo�q U�_���u߳����u]L�7綾��J d�NȽ���~�w�����Q��'�
�c9f�n�9y���ہ�	���_���̫�ӏ}�   ���m��IM�ζ���T�a�3LX=ô�!v��{�7��C��;@�#�j#���lƃ^�v��Z��A�Q��2���б�!�����#�����^ܳ5ܼ>o�<��i�ܹ�G��bMM�i�W1b�sƊ�`�jL��T�Ct;����3?�",{�Щ���)j۵���S�]Ut�7F  � "��P�l-��ͣ����'�u��
U���V�DR����A�d;����V��*^Y,w�trnX�A�	z���{���y��~�s�ٺ}!���:tHY|߷o�ٳG��y��#�^x����z!2qco������)S���ܶ�'��u]PAu/����Y���uM�E,�cA�S<]G����m+(��:�l������������n   �%��E:�e:]q��y����O]A|���� v ٣r/-)����4�~<}��?�1,>����on��U�sn*�Ǖ�U���(���  ��C=qZ���>��B�[i�����y�����d)�!����Y�R�b�&w�r�0{�D�;@����1*�`T��0��x�~����ӵTs�ί�����:JF8��^ {���޽;�C4��yx���o�7�?� ������`%�0����<�0���?�u>������!:b%��Ot��Y]�e�f�㳝whjl7z����Vx� �pA� P0��;H�6�MC�spW�H5�f�����-M�j���Πr�G��SU~��޷!�v,�a��Fu��Z?�u���<��~�ۭ)++��S�����z���t��Ajkk��9��Y���w�t��wd�iڴi��ֹ���;��Չ����?W��g��a͏J�=��A��Z�]>�����)��(J�ۇ�x�V�A	T�p{M�$z��x�s�    ��Ɍ�h��zq4N�D��^#<���Φ�4c����������ڄ������G�;'Аyqq]z�QTVZb;�w-��^��  ���S�c4kB#�9�u��,�Rx�v>��3Lq�!=�d)����n~��3T�����=ƨݳ�n6�OX�>o7Gw^�>�j>{M�����:���> {���ݻW��G.�b���=A~��w8��>"��`��"�y������y�0����+��Ϛ\��^�flO>�Ɯ�B'�P'��KU�%w}6z�N�v���� r	� ���/F���:kv5적�e�}�g�{��!�����1)J%���`�ngP�18�ݕBU©��y�5��m��k�^�ϵ������l��5�n����<����Ǐ���f�:�����]Z|�@<������9"��2$��d�L�Ϛ[�u��,6qX]���o�ǡu��5�x�l?����R�ҙ3������`��u��	Tn"U�@������H��J����8e#T�aG���bӐ0�    <k+iѼ��q*5�����@G�j���2�׼纳�S��0X����W�D`l���Կ<0|�8d��ΜsB�nnG�   ��l��ʎ	����۶�6�;5��=C���g�tO��N~�Sݭ�@�[2�a����{�l�u>��΅q^wN6����o��Ǫ����w��A��d����â��[4�Ỻ��	�߭��V��9�.K���ȏf�9����:�|a�/�@���\����G��h'���96>�f�]5��;��<�f��Ss;��E�i�fx� �܁�; � yi� M��AM��C��*KC�j�A��3� 9�B�jB{��-�n��B��qB&�Aw�k����ky=�e���~���ӽ���:��]�~ܸqB a��	���? ��w�X�������uww�G����k�:��|c����9��0:�` �F|��cT�F~]YY)>��dh]պn�~A~�a�Z��B�}�V�
�g
PjQJ>�Sv�J�rn^H
S*��CFN┛X�!NY������j�M��CB�}    @���b��=Wӵ���Ǖ�Љ-�)Nh�No��5�[p��g���x�r�n���n   ��}J"A��&��f:�b?�vw�c<C�b,'��tO�~�ݟ����/t���'�w������Y��u��չ��g3G5/��v��ָ�eo������'�eX���k.������9��x/�h��g͞����G���ȏ�{��<�����񱅱&�"��hy�N�vU������7Tc�J���T!w��m[ە��A����?�N�M�	�!  � � (X��i��J����J;��@���T��M��*^��dh-ns���:�U�@�
���)e;���݃���x�k���|6s���4�n������u�ð�,�� ��F��xX������/������M����O/�S��y�K�����y�?^kC:��s����5, �Z~�ya�7^���Q���WH�U���(۽�.X*'q�*R����[:	S��*q��|h(F�&ϥ՛�?Ʊ   |[�ݿ�2�p{�����;.�~�D��-�rG�    *�;�-��芦��{`��˩���3t�GJ0JD)���w6��N>�*�Ϊ��P��ݑbш՘�����l��s/k�:��|�s���^��~׸�ӽ�g:Y���8 /��dA?�k~Ώ|�\~d����c흃���a�{�Mx޺^���s��s\Iϐ��9B��X�Cz�\�%K�x�]���	
��
�Gr^ء�B��St
���vav��خ
�����_���Yz���X���1��<�Vo.���  @�A� P�<�%F�&̥3�PW�!�wK3�]��Ѹ��%i��*Z���V�*�vϾ�!-RY�a݃���������a�Q��:�i���u:�u���VX���d#@�AX�\�o.��|�)��t.�aS�q�`�v�✟��P�N�1���ܮl�c\y�(�K�6"�   ���	մ���PY�8��N�H[�"0��w��v`d�������T���c?  ��Ѫ�Et��y4�v%���EXr�D_���_(���tC�� �vhh���C!V����~�{ϵ_����=�����\'�yNs�Yc���5t��H���~�?���,̒�w���G>�H���",�\"˲�9�3ң���#9Yv�A~>x�_��~�k��a�ٽ�j�C��a{�z�v�o�s���D/�X1�o����������(m�u�� �� �Q���!Z�QC7M����6���h�r�n;h/Z�W���Z�6�w#|���N�=�k��o.��9�v}���z=��~�;����~��|�sE��l�YH�U���ۜ��=�v��W��M�2�q�l���L�J'�.�C��z�Lzb�8�@�   �B�ނ��q�0��W��v`徧�   `�=��Z>�.��O�v9�����_8����<Y����ٮ�]wh~��;�ɡ+M�Aw/ss�hw���z�A�����<�s��;�q[�{/��sm;d��s#z��Q���X�^��B��z}~���?̗��9�n|�!���zkn���Y��n��M��zb{9u � �/� F�D�~s�fMh�3'�Sב6s3�%��7oeeeC�i�*!�hemrWW��(P��|lCn�]g��k��o��}�nN�Ts���Y��^�^��{E�\�[A�W�Av���t��C�ʧ���j����.�Sn���v�慌-]�����l.�m�Z�    >�w��{�>v������c�\��n   �W:�㴢��Θ5���v���Tm�C�P�z^<Ä��=�3T7�K�Q��8�Hw>(mOct�/rnX�A�	{��|6s��S��3�m��:������~�R�+a}��\7J>b<��j�:��`��[L���j��3[�ݛ�UM�w�;>������ho�\z�!  " � u�l����j:�q�uo���&��Q�hu/f�J�ɽ���n|���]�!����	'���0ƣp���l�d3�i��|�5٬ӹ���e�^����r)\fם�*Z��l�j�nw�2B�6�v��v�(e	�Ũ�~�nk1����
   䚿���hׁv:�e:�n�N?��k �!��������i��ρ#]�W�� �B�    �yeg�*˦Ӓ�C�{p{�Gh|���.)����EX����T��̇�3����aw�9��\d����	Y+MN��=7��ר�yY���9���;�n��:��^���A�g�ȇ��{��N>������=_H�a��&}>��1؞��p清٭ޡ:Ю*Ʋ�=�ۍ��n;>?������ �� �Q��[c4�f6�;��:���*cC|D���Mv�R�J(E���;?�5��s�{��=)^�2�G;��>�n��\�=��a���F���@D�=���7�^"?�G�E��ȅ��{��F>E+V��úFX�v��}۝�!��l�n�i_�[VV��{S�Ϣya� D��2��������c��/��o�F�O���+� �Nl����?|�     �L�`�V��I�[��x/���f��������_(�C�h�'ˮ�7Xl��EYf��vW=�|C"��{&�Aw>g�����ָ��习�g3'�yNs�滭qZ��V�:~��{:a�>��f�>�h�s��c��\����j�����{k{�?��5�C���iO���7  Z��  ��5D˻�����г�L��!��屙�D4�g
V��uI|$��ʐzW�38
V���vB�݃��xPkt��g��|�s���^��nk�Y��ϵ�y��N�F�������&XEM��f��`��5�n=�_���ڮlO=7���ۇ��� U�ϥG�� Z� yd��)��_���*ʨP�?w.��O�Ow�!�w��        D�������tYc���n,�Rce��ʂ,�����]����ZK���aAw�\����x���r��Z��A�Q�j���uNk�\��5�z���+?4���{�0��ss1�a���6�*��mm��S�e-Ʋ��9�ھ���� �	� �1��7TϢ��Pg�>��A���k����^j���A�*IXR��kfP�3�V�\܅'U&�=���e�'~�=�k�\'�k��r���{�N6��:��f��z/���ڣ�0E�|	Wa�VA�Kt�fm��|ە��,����TZ���g���,���}�[��h���  ��ʳ�-�p���E-���>I�|�!z�        ���H���8���K�ͽ����!����Y�Xb�g���k�	3=ôo(�B�2,�mН�a�L��ۍ�������g�%�Y��:N��v���u:ku���Zپ�X"�?�l�1(1����^+W�b �v�q���^)V\x�q�p��_��Z<C���մmp��!r �肀; `�p�;N�7U�y��4�{���������f'�J�?�+u�]������&X����aw
/�n7D ^�:�^��9/k��׽F6��u���:��^����^�eX>*"ZP���x]����X�r���į��v�P�Qx��T[	*ũ�{��vǐ��qA!P�{����zs�bq�� Ѡ���F���w3��ï�������!       }��ѻ�tyc�zns�
u��Lb���$]�e�:�3L���v��_�]�u� ���h��K�z�n�}�l<� ��:�
�=
�\��پG�Av/��C���^���3�>�ڽ��z�X�?O��q��v�R,�r����x̰�3�C @�A� 0����!�X9�.�5H=v��*v763ȃ�(�6��X%�b�kc��]�=�Ҡ����0{F��p�K�=��nܫ��GPMU���a�SA	S^ĉ0Ũ��γ%��G6�-4�j�	V��t�l�	��*;a�*Nŕ�v��v[q�F���0���D�Z��   Z������Ӥ�U4�/U���:c�\��7K��       ���K�6��Σ���Qow��+4���w�]��c�6�!�۔c�����g�{�]!���;e�s� ���:����e{^wN6����o�Fw��z/���=@�N����/�@���B���v�]�7��ΥXv�v��K:�a�?T��Z|Ī�Z���@��; � �$�{�rc	�4}5�ޞ��f�J��n|���`If轘�܋�����@e|W�e��[�=��������ݸW�����`������09��QD����$,!�,0&���:\��e�1��p}1~��t16� ,�BB�&�
	�6�<;;3;������]�U�=�=��<�U����ݙ�>���mC{�Tq����S��+�4� �$�!�%�̨k,�h���v�Z���^��.3���/(��v��JmW	T�k���v|f_��qS�"���f�'��/F7�ԝ����o|�m��c�A!�B!�3��<~����;֠8u K��Z�,���^����X���:_FY/�%e���F�F�;GU\)�B]/n�1�qI�������5�o�Nܵ��f��e~3��c�������v0����f�X���d�g��G�0�4��8{&��{�\��CBHgA�;!dE���~����vL"w�``���T�ҋUA�{:dr�Y�p:�:��,�=���5�W�"�AP��*\�i�=�fN����㌉3N5V6^7G5�d��:Q�L��Dҟs���E��`պ��ϯʟ����{N�خ�D&��P��-x�)_Q���n N9�������8s��j��BړO�� ��S��������΍��q�'F������_�'�� !�B!�t�"p��"6�]�������i�(	�2�f2�]�3�w�齱��I��$�����V���϶��c��/�c:W7�f��k���F��c&��V����n2�]j���f�	e�4���Ac�>��ZS��}>%�]�%�X��G&��;gFpxw�҉��NY����mc�q��4f�Ψ�ڑъU^�{Ɠ��ن0��`"V��M��u��sx�!�'\�m�=�tN�}���#��X��y��6kخ��sڝV�ZI<'���Zi|��*�9I	SBc�����]%L٤.�M�E��]"N9cu�v��� ��p��"|ew���A!��'�~ ��ǿz?>��W��'oю����~�Ÿ��u���*��\&�Bl�����ç�y�����k^�}=~����U95��>t��D!]��s��!<c�*�^:���Ey0VM�Z�e&�t5+S�vk���B](�������jT�BY{+눦�M��yQ�u�G]�v=�X�x��\��&�D]ӆ�6�7�f|Nq׌��(ɱI�[�����L�6�a�z�O�����vQ]�|U�����QR۳==X߁��:�v��	!��R���B�Ƴ.ê���U����D���g�s3�T��p�VoA(>ĦvS�;R�4wS���7�pՌ���ү[?�:��َU���3�k�F���>g����%�Z�$Z��tc�!h��`9q�s�3�#,T��)qJfrڋ�R��$/8�v���~`)�!���053�_�����%xٳ.3���{:��e���Oczn�B�3<Ћ[�������+�?åx�{n�<�'ֺOܺ���g��lZ�
����@!�3��`�}�p��<.�:�Ɗft��ce�C���&��L�T7��B�|5�XFwu V���ͪ��J2�j��q�����ج���V�>�z^�k���۩��R�n��z��nin��u�X�ݞU�C[c{AQ?Z�	w���	�	!�����،7/	E+��@� �5����U�av�&��7��z�mA�2�����o��bV�;�NQ�+*-���*[�i9RLװY/���@+���ψ:��(�q�(XE]���v�0�0�{�f���-�>A��Id�6�����}xl�����yBi>K������ޣg�~�ќg_�_y�����I�>r�B���?�Gs�CO6��{�Kq���:뽏c����J
=!�����b	�}<�K���%}'17;�B�����Za�������3鴴f(JxW�
EFw��V�Z���֕�������؊Za��	[��['�I<�i��g�f��m�'Q4�jS��/���}���ZTG,�$al��ݭB��EiZ��~hR7��XC�8�[����3!�����B��/TD�+7����1��]h��%�"����^7�ׅ�tM�R�V^c�hB����]dr�}BCu�@kJ���B�l�8k���g�jl��9�sMְ]+��q�򱵻8���׮��J����^��w�2��)��=���$�|[

��u$qJ��༎XۉO�w��e� ��N�����[����f�o����5���'p��y#���������$C�?2\�͘�_�_�[xp�QҎ\�k#����+J������G��p�__{�x�SwT�3�_�[�ɡS ��P/��]�ŵO����P?N,͢�x����<��!���<z2����q�I�`i�X��.�cej;?�ꆞݟӁDw�Za��.��ꄲ�Za�SW�5�Wi���^��(곙�?꘸�����k���I=�ShU-2�s��_N3��85����Z?��mRs;�glW݅��ޠ,�k]Qu�u�R��:ar+�����3!�����B<p,��ӫq�4J����(�Fw��r��	T�d�h%JbPA�JezwE�PbC���	W&�����(P%adoq�V0�)Z-F��Yݡ��rW�)ZQ��k�	S�6��]fn�S�Rja�����-�S����<Vo���8��vBYN>�����s���#�}���#��_�w�ӝ��/��q^�����^�K�m���;�ǻ?t�Y$"���;7�s�y=�{*�/.������
��ןǱ33�v.޼���_�+/�To���]x�-�$g�������w�?u�Va���<�S�gnw���V^/���>��B�\�E���El^��M���ٓ�zB�X���탱j;=W±j��tc��t:S�:uÒ�(6��0�;���vqHVR��f��ev��3&�8��(�esL皬e���Y�$����^��6c;����CQ��=G1������R�v(���2�ڄb�r9�N�÷N��n&�B��	!D�+Z�l�s7�p���Ƌ������
ƂU�^��^��i��u��n&Zɶ#T��+S@�
&4�W^�s��[)^�ε�Or�l��zQ�U�1���o�NԵ���f���Z�ώ��r�VI	[� Xٴ���ʟ!a�&q!hn׉RraJ����D���v���T�v�Y5�������P��%��*���=x�;?�y�k�qrT;>�I�O��\r�:�����|��veۺq����I�~��w�'�~�����g���.ϼ|;���^�_z��v��W\���66<�_�ux���H�3�׃���ո��m�����������ٲv�?�7��6B�|O�q�� ��t1��8�/�IC�t�X^c��v�A!]������j�06�7�%e����4�CP+����^�.��$k��#��X�x��\�5l֋�~7��zc��[QG\�b�1�T?tk��ks���6�#z�5��4�Cݎ�E���m���8ݷw�uj�Ԛ	!��b��|�}<�K��ē�`���P�*8i��v�A���v�Ӂ4w��=�ۊ�6����.<"Wbӻ;O'8-gC�s��o�N�q����9����M։�f���T���-�p�ѪU�vݘVVI�	�Q�k� 垅�v�E)���.Om��.Ȅ)�8���ٞ,�l�m�
�ϖ���n<��D%%���z-��u��'Yy�����ƅ&��#�tJї!�DO6#l���w���1z����7����W�˷����Ư���R��N�E�=�����w~�B�������$nڱũXZ
�b	v���EuB�>�螮��ݟӵ���^<µC��=���I�0��@Tt�hM�^�lC{�Zb��Q�Q�wl�9�y�kخu�($Y�l�e�S+��Q�$eV7���N�6�]������v���X��a����vO����܊/���B��	!ĒGN��hjϽhٹ�X\\�T2���hUOe���}�L���c�V1���/�������/��fn���k�g;V5^5G7�d���k&��v��WR�k� e;>I��J�T?c�"���njn���4��S�����;���;�z�:Ѓ��o� ��n�1���|����YO�a4��/����z��=�ĩss �BV����s���Re�V��<\�]�����Ç��n��y�D�8	B!�A��������u�9}�������2��Q0�~UIt���+��42io������U�CY���ae-T+����ܠS�qj����1����	uu�(�E�<��6kE]7�hJ�Ѭ�90�'Y4�I5BU_�����ިz��5C��uĠ�=�`,��a��S��}dr�ur�v3���r���B"P*�pϾ�6���K�?}H��P7�[�V��Zz{��^3��ū���o V��V��(��c|�E,��=(^uj�m�16�Dc���g3_�F���z^7ӌ�A�5�m�o�e2�S+���L�
�	�="�J��nl7���2S�ij�t;A�0���02��yfw���!���[����_��o|���k��\�k#���7�����!��R����#�|��?����~�>�G��h����w|0����7]�?닐I���;��|��q���#���!�t�g
�m�Wm܅��0;��f�Z��ce�i�3��au�g]�Pot7��j���ݩ�ðD&wO���6�����Ю����7g��X����t�mױ]ׄv�Z��fR�n���v|��u��P?tk���`��gh�T���!6s�ga�Г�^Lj�g��}pdGrk�=Nb;k������s�|��vN��U��03uFlt���]Ѫ��P۽}��N�Bp+B_�{����Xw�_�	Xq������+���C��W��:&�$Ǜ�3�o���zI<�i����s�md��*C�ɘv��)���ڤ����8��R�X��*a�4yAgn����ف�𕽎с���iʿk���_��#��_}>���v��uc��{_�W���x��iB!�NoO��x�;�c��������ct
�����/�o��2�h~�_�y5���7�>p!�t����j<�����Vw�ݣ��{��i��d�p�P���EuBU��^3T�
h3Ǽ^���v�c��j|7�k�N�5�~v�ӌ�3Κ�TGl�����=�z��0Kan��
��v������r�3��w{��:�k1y>��<��!��Dhp'���s6��SCx��1L,��¢��.2�{�L���@��$�;/�3&_�J���"C�N�Bɟ�Jw�
Yu��T���iN�{����3&�8�X�xݜ8�Lֈ�^�g�t���R�J��n:n%V��=���@�����f�S!c���]+T�Rڝ1����ԉm��~ W`�!�t:��>�9z���:6ܯ�qr_��o�k��_�Оc �B�����[^���%�o���o���½������;/��'�7��j����{�B��B�T�zrp��qs��C�l����X�za:�������&F�p@�,KV?@#�]P/t��Z��T/����K���u�f�u��(u�8u�n�ju-4��E]c���PC�:7������m�b�j���y;>7�v(Ih��<Wo�=�{q�N_!d�B�;!�$D�����ѓY����P:w��� 2����#Ni��Gu���6���kpw�+q��_��
`�v���J�R�VH�&5x�j|���,P�R�JZ��*�A��K������%Z�����v��=�2����>w����+J�
Tbc{8q�&�����Z�	�8ևS{��N!��7ڋ�����xu%�U��� >�'�����G���� �B���l�����MO�X:��Ǐ���/�S����s�߾�Ȥ������N��/���@!�{9s�������ɝ�j�<�O��E&wQ8�*KT/,�ϕ��t�����[4��YP/��~X�!.s�0�z���g[�z��:a3j���;�+I�[mog��Z�Y��u�V���?	û��n��^4��°LM��@�(�v���X��G���,+���I<<;��vB�� �����0�B	w�.a�+����ų��"U&S9g<��x�3�{��G���+)�{��v抅�F���]eh�ۅ�D�B�>���;w9��Q�u�G]G�Vܱ&s���͏�V��mh�a��ĳ$?��ku�hWpҍi�`e���Kk�S6N�r�('��D���*H�)�HezxS�[	��\.�щI<p~�w;�v��	!��w�,^t�?���r<����}�Ļ^������g@!�t�����x9n��	�1������),,u���N��գ��.ߎ�/݆o?r �B���g
�cWoZ������ka��>���f������F�{�V743��v�.Z�e��RJR/���F�$��~լ�8���c2O5�f���xF'ӊ�c�hE-�Sk�]Q?�=}����=j��ol��G����5�����ކ��w�s�gBq���B�Ĺ�">�;���;p��,f�G��Ne����e�����3��(d���sc+Bw�´O�*
�)�x�No��D�RP��Լ�R�W��̵헍1W�R��:G5�t��ZQ׍B;�ϣ���!�ڝ(Z-�`����~��T"s{]�
�SPS��TC��T%�0��.��m`0�=�8�D"U��ў��s�#L��N!�ι���O>������M/�F;~��0>����uo�B!�»�p3���'J�S���S8~v���~�۸l�z��Y�)ǽ�Ƨ��N!+�����`z7^���#����vۚ��ѽ�F!�c�����eY~�{��,�}�xh]mPD�^��Wͪ&mx�;�d�j��\�5l׊�R%ɯU�k��jh׍i����X`��α�F�
�>c�[O�R;���~�w2&/¿�-"_����M!̀wBi2����Wo��2'1w�|������t����zPbt�$4�[����긆ѽ0��ī��p�%O�{I��,�������(╮�*۔�V�2��ۮc���NHkX.�-����n;����ɘV	V"�{4�W�i��SAs{�^'D�M������h�T�ąb��n+N��$i�nOo/��[��}��S!d%�/��y�?ށ���{���d���;6N`��!���!��l���9o����}��-���x�;1>2 3��B!+�|�koý�p��"rg��Fa��1�v�c��F�U���Z�LwOůF�V��k��M0�m���(�Q��'�u�n��|ӵ�X��iv�1���6�یo'�{�L�?������ZX?Ԙۣ�c�R����n�2c{QQCtk��`,Y�й/��X�	w����"!�����BZ�}Gr�~j�ܶ�G�����j[f���*��=]��F�t�yX���Waӻ(�A$T��#�w\I��P���jv�6���Q�����5]'�I>��h�����6�����_�����e�vq�^���Ku�)���7��D)o_P�%/�D*�[���u(���8��~�B��|�'F��W>K;vx��wB!+�o�`/��G�mL�-�o>{/����@!��]*⋻�#��0{������R��Za�0+����]�tZ�%��hlv��/F��^��Kv�@{ۖ��n�gL�q��Q�����ͷY'���,�Y�]j���en��b��[Y?�ĊR7�����}��'ê�-�۵��ڡ3ndb�sv�/Կ��B���N!-�TJ����]���
�U�!��]�*�
W��z��ճ7��*<�fw�V�A��3���UB��ZD+�`����yY��~]��[�J׿�U3����1���k���I=��i���ĳ���ܢUR�V;�ڽ�2��J��\��E����]����N�!>U���2c�I
���^_�]�z3�u�'vS�"�Re~1g4��� �BV����~�#w~oճ0ĤvB!����^\�v'�<p��S(z�5à���p4�t��^pj�Հ,��銮��
�y�T�p,�к@,i��фe�Bxj���)I��m��Or��8��(�ustsM盬g][��l���|���m�v3���4�~轎U?���jMj�~S�8KV;t昄byw{V�
��à�]XC�axt��V�+{���B�C�;!�,sK�J:�X�V<ws�gU^�z������D�L�$_Oi(��kUE��V���oBC
�t�`��+b��U�6�@)�����&�T�cf�X��~�x�Jן�@�t�B3tsT�L暮e���Zi$�5ie���$+�q�Ni��*W>*<���.�l����H6��*I�ab���.��y�L��}S�ط��!������.U�)�����R��?!��Ng��"�}�_v!�������(��m�K�1a���s=��S3decc5v��xj�ձ��u�X&�wY�[#,���B�{_�U�FX��k���4��g�4��̍2?�:6k��F/�c:W7�t�(��褠��y&��V��U�_��iW?\�ꉡ1�uCy�P����j����Xn1�ecn7�r���!Ln�W:�����ބ�hp'��e��B�۝��n��O�g�b�#RE��9����h��oE�Mh(8�����P��"VY���L�$43�'mv�2�t�8���c2O5�f���xF7�
1+�gD]c9L�-�`e*J�*A*hh���P:a*(R�D)�����S۽T����ctb��M�ѽN:/�)B!�z�w�
�m_/��*���2>��A!���`v~	�B�	�Й�<c�zL.���B=Kdv���[� �]U��Za����Ou�c�±��Bw��Ю������Ix/٦����n�/c:��u�f�Mkw6�I�WjPV3>�kv[(�ɘV�ڽ׉�k��u��9�ebp��ښ�m������4�_�W�+�vH!Q���Bڀc3|v&�ͫv��0w�2�=�1��ݽ�����y�"LW��p�	�ݽ�U�DwU{5L��aP�j$�7�W�%6�&5z0����c3N4�f]��U�L暬a�V�g$��?F�;I~��L_���J1�dL�M� �d�.yAdjW����5�&N�S��V�R�������V��}��=B!�KO6���W�K�I�8�Z������}B!�{��+!�;
�7��ѽ'��ݖB��,..�j���,whC�{#�V3�
����ݠ3��kvO�����p�p��i�P�elx70��k������7g��X�x��<���kخ��ڝV�%�1�f�r�e�QL��Zb�@�(�X*C��nX�����s{�f�����n�U��Ln��SX�Q�]C!$
4�BHqx:_>��5�W�������*����4��E,�V�+Sߎ0lv�OtW	XJs���
V��╍��;V$^U�,�@e*:%�����k��g�f�n��f<ힾ`;�U�v�1I��E����.PA/N��(}ꂙ0��m#�M\T6�	����^qjpx����N���B�d����m/�O_�K:��vB!�{�U��B�=�B	w�-a�w#��������=�0��k�L��Za�Z�s�a��.�Z����ٽ��:}ڀ,Ϙ�x�+�7�;$evO�?��q��I�Wͳ��[#�zI<k���ץյ�f��P,ﵸ~Ni�^�������bi���X��[p��fN��C!��	!��}�P>�����������>�L�G.V�CbU��6����t(��/Z�����u�v�X���̠.�/X�E�� ։U+ĩVSq����⬳�fv�q�����W��\��R�I&�TP�2M\���(#a�.H�)�(�^�Sn�+:��^c{� �$������_^�K�chn'�B��|�wB!�[*������V<gS�g�w����J��*�]�Up�f�J��thY��,ѽh]/��9z��F(���>f�f��S�Mj�ɼ��۬��3��V��#+ʼn��^��~hS;����Xn��&KW/�1���׳r�y��v;Fw�$������Bژ����Fq��Il�I��L#�0�{��A�J.V5��΋wg�\��
P�T���%Kso�W:s��_���	V��aa��A�j�Ѹ���������7Y'κ6����Y4�s[�j9L�E�*J���qE���)[�{0�]lj
S��V����8��J0�䅠0U(���ߏ�ѭ�}����	!��y�n�/�|����vB!�����!���L���)lَ��-b���J U�&�0��±d5Co{�����T�Y�P��Ov�6��4Yh���kVI��^��_˶'���qꋪ�Q׋󌨴����?�V�m�tf(V�OߵI��=�j�qꇪڡ��4���É�ạ���&˙;�z�=ч�;����B��wB� �}(W�sWoZ����1;=-��I�"�J���	Wn:C8��MhHi��Tw[�J�ր�f� ����$*�)iq���6�DY7�g��!t%��8k,w���R��Ȧv�E)�X�JYP%.xSt�viZ���^�T*qJ(X�b�����o ��-���"���!����ů��:i?��B�ʀ	�B���L���b��.<m�fN����u@�]��j�DwQ�Pov�����B_}���)y�!�.��m��b�_߷	�J2�*�8�X�xٜ8�L�ۮg��I=H3?��Ċ2�SB��5�h�C��)&]?��E�<�M�f5Dub{�;>;s�'7�N��n�	!����N!�}G�c�z�jlϜ���s�4�um;B�m��>�nr��W��y�������TwSs{���L��aqJ���k��J����Q�����7Y'�I=�[i���U3��c�ѥ,4�����Ȧv4)��Qڂ���T$�= J��)m�T�j��p���iJ �bƛ_t-���gJ�in�l~꒭+z��r��?B!f,,�A!�4�}g����v���Dw�.вCU3,k�<��y���^ب����UcP�'���uB�k�:�{wl�.X[�cE�6��+��g�n~����mB;�e-w]3����n;���?=��{+S{m����t����^�%��k����}5Ī�ݴf%�bl_��?;�}{��{4�BH����B:���}��0�]}S�9w�BOU�*��v|��4w��cvW�=�n:C]��$4�5)��?��4��F�
�W�������L���֬�i/�*��׼�t2�ɚI=��h����s�-}�fl���{[S{Q�T�R���L�!J'L�M�6�TE�����il'��W��T�ɛ�/���y�s.�+���y�������σ/�=��O��� ~|��z�O@r��BH�9|�P>�ؼj�>��4�g�XYA0��fX�/hk��`,�ٽQ/�	E�B띠�/T�N��ژ݃aX���k�����Ǌ3�t��ZQִa�M孠[�l�%Y4�|(����#��S?���Mj�E;>G	�
cy�����ؾ�1��?3BH����B:���� Fp�q��¬ct�d�[J��u�����Mh���S�i�v��*lz�W֢UL�����,�ݡ�w�ؤǫ���׭e���Y�$�u��^3��6��&0$���^�)�����J�����lA��]������.L��s�@�F����E�4�B���=�/��X��I70>2����yx��n!.�_��닰k�d���w��%>5Bځ�S���cgf0��Դ��d3 �BZ���|��ݯ�\ąSG�N��B��]op�c��I0�,�]�t�/z�Phv�^���(�����V��p�8�t�mױY3�����&����U�3t-�ދ�[ej��AX��D�nϚ��vE0�kl�ޙA���B��	!��g��T�(��*�]w]��3C{�Y�L��^��Fw��]gt�%ZE0��Xa�_�
��t4S�R�Mj��<���kجw�n�BVψ��r�Vq��{��]�� � ��(%J[�Q��R=e!dl�R:a�(��+F)�)�	!����W��?��e��=����[p�3Ǧ5�p��eR�K��3��e��n�j������7��rL�&��7������~�F��A|�?��󝸰�k�s�{Y�#��Z�F�6�ڎk'��Fwg��[�=fwS�{�Z��N���mw�v�]��R3��vh���:8�U��V�	��M暮u�$��h�ע��XQ�td(Vm�I�7&����n����kl����#�B�L��v{.T�;�z#���P]#��.�5�_�i�{�p��)�=�D��#T��EB���^7�=�fFw��]gtOJ��	Wrӻ^�RWĒ��+��g��Q׋�~�a�oW�,ɏ���U�dbT��&��)�Y$L!,P�B��R���onۃm&��+JI���8�����kq����B"s͓��÷�
�=�V��I7�fl�wR������7r�{��I��ן����عq�=�G��h�3��4!�����t�jtێ�O,`���ݟ� -��]ft��ܫ5�zm�`Z/T�dk�&�l���fA}��s4xO�*C{��k���%�c2O5�f�5�zN�Ҫ�rbE���X�{��]gf��Uw�N����i��e�=ۆb9׾�����88�	�9ُ�4�BH[@�;!�t!���>�I��q��fOEڛ����>m(Z5�_R���.Ou/
�դ���e��^;�J�t���U�oU��w[K4.���9q�η]/��QiW3�	�����n��M� 7e�'FI����v��]�� Ml�l%hcp�R���U�8�I�y(W��i�!��˶�ǿ��5�����N��S�x��)BH'����'�!���>W(=X3��m(�p�0��4wQ8VV��n�tu�碸^�	�Y�-?�M�nOY'�uBQ}��0��k��Ú_+�p,��&kDY/�sH�_�Vb��Y�P��g�P,�k�I�eFwۺ��~�6��Ų�r��'7�;�{pl��Ec;!��4�BH��ӹ�ы�c;+[.�9Ry���U������L �Amp�EFw�x%��fv{�*������9��%�9���cM�ę��e�(k7�٭`9Ŷ$��*#��$��{��=x��`.F�V�w#S���]kj�Ra�z�12�?��
t��w�)
քB��k�$>�?�����4��n��o�:�s ���	�BڅSs|q70ҷ7lR3G���X�Jñ,w�6��
���ڢ��]it��5C�w�6C���Vخ�X��6kجw�n����$�oE-��k��dvQ�����6�G���ljl�
����d��l=�[��i�;�۹�3!��4�B�
��А���필�⹪p��nC(Hq���%��kG!�nW�9[6��īD��oM��gub��oKoxwƸ�q�)���sT�L�۬eͤ��-4��mu���<��*�)x��'�IX��ݳV���%��L*�ąVۃ�T�ޙ;�z���NZ;�X�B�m�8>�'��ի���4��n��؃��u?!��ѓ���BH{1�X�����ܰ%�U��1��n0�%�����Xz��xG�X&�`[��_3t��n��
�}���5���g2�d۵��oK+L��V�l�@��s���.Kiw�6f��M}Poj��뇲 ����8�C���?Џ��|� 0��vBighp'�����0Է�ڒBj�(B��.�l�A�*$RL﮹=,`�ܛkvwϦ���3*��-���]8J!dU׷���ʠ�o��͚I?�]i�����Zad7����6�%Oi	Qq�)[c�wKA�%�B�$Ol	T6┱0%Mj�
S�ԁɍ��>��@!�$������^W9�p~O����E|ꞇ@������i�&�b��H!��#Ky��}dRk�S[2X�S�;?�L&[Im/xM�
���t:��!��U0���.�#���}ú2˨Vب��;3K5�t��Zq׎B��ϣ���#���6��Ƌk�Qj��P�����y�P�'6����v��(6��LﶡXEo2��v�0��142�ٵ��@��HS;!�t4�B�
dn��;v�Л]��l͠g��/�V�+�P��sD���-hxw�&�6����H<��*�>~�{H�*�S�e�jbCt���?xWH��0�����5]'�I<o%ь�I��/�'Q[�v�lml�_t
�ۘ�U�vS��q��:S{lc�H�*�����̃BI���A��ǯ�$�����B!^F�@!��3����{:�8�ܰ�����(d{�fv��=_3�g"ݥfw�`,U�0z@��͘P��5�W)j��tw�{g�c���ͷY'���zv+Y�z�rbE�ۑ�Xh�
��q�Q�������2��$�+���`��WM�8&q�\��f(!�t4�B�
�Ih�ko���mO۸���c��I��[����Q����I:C���¦wo:�_�R�uVbIn_������W���V��qL�9&�Tsmְ]3��t:���xN�5�kf���ڃg[�*�������5���{]�
T­���R�c���(�zW��X8Y��A!����	�0<�9�/��;_w#��e���1����vB!�����Svl !��)<p,�0��n�O����'�L��@�����`,}8����R��lk����q��=�����a��c���7Y'κI?�[h��w�V�bk��1I�����Q���ݞm���FvuP�M�0N0V�X���:<va̡���	!�ӡ��BH�MH
���>b��.\9���3G��吕l;4��W�6_2�"��'ZU��)�\�����(����`�m
ux���F��P]����bD\Aj%
PqI�k���(fvQ�J���k�ܳNhR������]-N����%�(��n+L9���$��qW%q��vB�^tݓ�O��
t���V��	!�+:�?���^S��zA!�t��!`��N\3�G~�(�&wY�6+X7��c�$uÔ~hS��C�b�Ѩf(��g��=�i]�O�±L��曮eݤ��δ�6���X&s��Նv�b��.�/F�ǩ°T�X���1�;=[�5D��{��F���>���s �ҹ��N!�Ǿ����h�6<cK
��cXXXP�ӆ�h%Mo�T)���#V�,u������ ﶇΆ����+dU�*q*���%Jp���-`y�)[A����4[�j�p%����P�v�%IV�L41��ۓ2������K>!��KZ(9�Yj�h���@0�;�6&6����س����@!�DO6�w��ft����3��B��u�n��.���ĺ�a��/� B!��9|�P>R�݂�7�'qan��ӳ. +b0V�:F0��f���k�q�����u��|g�ذ�]M�.hj�O"K5�t�n�(�%���H;b�η�#�k��6+C{m�V�b9��&5�j-�����I�j�1�����&|�H��P�B�thp'�"��b	w�.!�Z���҃���9w6dtO7S��4��vW��W�_̒	W�k���!�p�4��g��G�

Yr�Jnz�!(�J��#J%)�,�Y�]�$?;V&@U�۪��4BTm��=Ч�T�]֧�䂔{�
P��D�*�*]b�N�*Z�T}����&�{$���NZ;�)B�D^�`�1tnr;��B���'�)�����!_(���G�x���#��t���%B!���Rw�2�5�r�zl�;���'�v��6fw�v�n/ˬfh��N(4�W/��@����\�W8Vu��Ȋ�n�u��bU���ۣ�U�X��ø�X��p�Q7�٣��,7����l�
��cx�N�'��9*_�!�t4�BQR(�p�A�D8������C�1{�DE�		V5�Ig��m7h-\	D�T$�{X�
�''\i��:�{@�r�t�"ӻ_����-U�C*Ԟ�0���b2O�f~^�I""��Dl
�Uۍ�����>�H%��������.3��)�/(L	)ߘ�Z^*�@%�T&�|>�щI�(M�s(w�JEB�\.Z?�n�5��Js;!���=�6N��%7\*�[���ʹL��x޵OԎ���kB!�E��>��#y܇Al�؅+'1�HE��x��@,�]�ͮ��R�z���ݮf���~]���u5�(�X���	v5�v	�2}F҈>�N�?._ V�O��`}Ѥ���хb�ꋒ�$C�d�2C�I0�p�g���_[l�m���*��;�f~pn?9�ݞ	!�����B�1��!`��N<}CٹX�_���t��]gxo�W�����6��d��^,`9D1�[ޫ7���M��P��$Tɍ��5S����L��щi�%|EKè�i�'2���M���kk
~�)x61�R:a*(H	��KQ��$fv�*$Li�|�g����p���0E!��w9��������4�B!�8��o���U4�?��n0�����o����q�}�`�5!�ҩ�;�/�ڎ�6Q:���v�B�.жuC]0V��(Ʋ����8�w�}�&tv�Hk��;<}�p,����F(C��$��&k%�~3hW3{�?�$�����p{�Ϥ�(5�{��bk�"c{5C�ݻ˳��=�3���^������ݞ�ñ$��j�{}�}�ݞ�s4�3��BV4�B���\��v�#\�+7f���OW�U��$��L�:�*hzO����]���䞄�]kx�VB!�}�h'8��(43�˷5ԭ�Ώb����� ծ�R+��5������r�{���׆��(���ꐛ���T8��+N�)�6�:qJij7L_p�9I?ëVa&;�of�P�"��n��؃�����]����Ӡ��B��1���_|�����'K�u���5?}��-?�5|9�%�燾
B!�p�_��7��j�6�TJ�env����B^3��=s�5C�"Z���������%�7��&�d�f��	�
���K��D6�{�k���X�`,�:���.1�;s���D�j��ݞ�q��<���BV4�B�Lc;�~lىk�*)�d�u�J(b	�+YJ�R�&4H��A�k|O����M�a1�!	�*$by�)Q�J��Yhl[l	Z2�Vc���6�W�Q�Gp�A|j&I[*���/#�t}F�g��Z��
Q2q*	C{�^$FE5�{�R@�
'��|��ȸncn%.�)�(�����þ�a�Y�F��!�t;������!�z:O�Z��q��!�b�cr��?�>����g�I�q�hr��\����a"�|����?B!��������Uy����l6[��j���mS�Cm)O���V�Ɗ��Jw��ܻ����>�ñ<�m�p,d�>��]_wl���8G'��b`�����k�a�����{mSOl^(BuC��]\K���D�����S7��h��*C���.�!gL>_���A��F�w��9�D�bB�J��*��Bڒc3|q��l�u[2X�������f�v�p��.2��S�S�kٖ�jӻ_��9؈X�kibC�F�2�E/�������;#��ޤ�O�hl��O:T��X��]�/�E��Jl�]��'�垛'N���p{��.�����L�R��m�*�@U�D┛�>84���GҘ�˴vBYi?K�8!�����x��?�����O���o��z��/�d�C=��������!��88W()�d6K녢�a�-X3�_7�c����p0V�P���R�{� �{�3���r�Di���F�>	^�n��xm�L�䠬f�@u_�����^�7m�~\�5EUm�=C�̃��;=��%͎϶YZS�4+���1��L��E,�v�BBY���N!$Qr����1)�`��	<u|KSǰ��'3��	vF�t`{BW̒W)��]$b��+�	���n{:{�A��v-Jx]����M8͡*8�����G�7C�5��x;C�h�8󛏍9]=_��L4���^_!���{�2��LM��k[C�J�
����!C{@��T޴���]gl׉UAQJjj�;��\���q�Q����vB!�BY)8&�7��3���{9�w�������4���8z��`���9���?����BV�z���q\1�C~�H�^(�ZV'�ޛ���v�n���B_�Ц^h_+���	�7�6�����z^�Ɍ�*�L�Y�ݩaH�x�J�r�����Ƅ�����͌���tufv������C�t�Cq0V�nhalW��U�DmZ���2����3�4&6��s���!��L!��B�ƞӹ�Aov3�٘�ƞY̜9^IiH��+���+`iīHF���� �\KhxoM��Lī$�J�;�bV��v��F@ਜ਼�K�Q��1�D��2'l���,���.�W{UQ�g�ƈ�ebS�^y]�Wؽ׆fv]�I���]��`bh�R�T��v���I[���j|�hg�0��B!�BV2�|o��O�C��7_��UC����_��O�BY��;�/)�n�������?7��ct��fw�u"�X���XI�ܓ4�k�)�p,�4Kb|��냺ڠ�o��wN���l����cb0���~=q=0�@,��=0�& +JQW+���	�2������K%�UIhl�����k���v��a�����<:>����~���3�B	C�;!����T~r�A��H?֏��ի�Ν���d2Y��}���uaʻ-������n*b9$ep׉Y��ꍱ�]�X�{�7���<�T,2����S�D�Jm�H`=��1V6��05��j�6�*1�='ip�nl��BT�2�{��8�v]�H��R�4��f3���G���#Lk'�B!���1�����������\�t3_��Q�z�C �BV:�KEܵ׹�Ήո|"����X\X��b���@]]P[7ݽF���XqC���Z�c	�M±t�º�����6hRT���z�x��-�h�g$]�F�0,�q��P=Ѡ^(�K����u3C���X��v_���v�nϽ}��ۈG���N���\B�C�;!���r|���g����tmO]���c��s>����=p֙�e�+:�E���=lx��M�+�������,�����{��%}J1�+V��6�������X�3Ë��ϗ����<{q�[�)<_7^g^�iE�ڽi����4�!��]��P��瀹]jl7��+��$�di�θщI�(��;�
ȝv�nL[ �B!��<犝8��?Z�{>yQ�����۴I�́S����7B!�Ϟ���B&�Wn����Y̞=�\.�4��5�[�C�B�N�㻿�'���[���e���u�޸>hXԙ����Ў�|
�Aͩ)FC����m°��e���������D�qk��5����A#�8˭�k�>C���]�ebl�����58Q���;�|�X?$���wB!��#'��#���\�9�u�)�?{&�� ��gK��䨋X�{J%b,�x�>��w0���c��2!+�}�-�iڼ��pl��Peon����U�iV��e�AqI�f|_k3�tF��9I��q��Sz��+PM�r#�IR�L�2��Fv�UOiS�C�H��}��G�9�E)B!�B!z�$���J�|���&��x��?��� �B��B)����q�1>��l �g0;=m����n�h�0��(�=x��
�ꄭHvW���x���*�{���*k�A�g�iM�δn:����x�?.��A�`a�@��u̍���i_�v�@,�0dj�E�DO�дVh\O���C��XX��<���}�ѝ�CB!v��N!d�Y(����~������W�$L_8�s��@��3��|	2�{�6��	�2�{c�_��wHB��1�{���4��{�i�XFm�>����k|�%�vEfN��4����6���BT���>��mL�"A�onOX��U�v���'����3ۏ�����)B!�B!v8&�_�����w�Ͼb��������� �B�S�Eܵ׹Ǯ��x�x��cX\X0�jB�P�%2��j��ڢU�0Z-���NhZ��_���>�z����f�h75�{��R��x�:m�]V}V�������^(�������c��~B3��.�%}R{�ڡ��.2�g2iLl�޹~<pĭ@!�D�wB!mž�|�pD���5���W���u��(�]`z�	X"C�Ѷ�³�ɽ��nfh��٣XqD*��]3&t]m�ߋڂ�y�8o{P3�2n�	
?Q���L�CO�hh��MƘ�EcTb��.6�{�%�(U=�)�e-T�"S�̮��&���|�����0��p�S�W��vB!�B!�XX��������ϼ|;:����wp�� �B���3��B_v��1����={�R�Ig��P,U���쮫z�}ie�P`v��e��t8V�s�ڠ��%m�z�uH���g��]�I�`���	������%;����E3����b�ñԻ=G�!
��5Co�X,T��kq"?��<�������!!�����N!�mqūLj#._����,LG.�'5$`r���Hh���f���=$b�c�X|Xܒ�Y�8۴��f���Mfz�{��k��Dka*e=�:JA8Z%<Iƕ$}Z㺤-��`"@��L�D3�W?S!J6޿e�����F��%7��(YH�Ҙ��BV��qc��#%�NAQ�B!�BH�8&�_z����^����-_=~�4>u�C �BH|�%|㠣Gb��"\�1���fΞ���LC�du����Ʋ�	Znld%���Y٦�Z�a�j�"��M�b����z�st�D��i]QSS��ez��%����P,��]���~���]bv^5�����#��^�	!�$O�*��BV�����@��Vov3�٘ņ��p�x�[:m`vX*K�������^,^5�MM�^�ɤ/h���9�����鬒�#�v�O �Ȅ-�8� �K�z�|eo�`�#듭ob^�]�R����1���Yڂ+DU�eb��ܮ�:0�P%2�������R8���:��B!��9{~�f06��k���s�!�4������A!���b	�T��A���5�W�)̝���
�I�2�{û�v(�JL��Z�����p��k��5CemPV+Ԙ�C�:��F(��ψZS����(�X���<�qB�Lj�&uBU_��<Klb7���&�X6;=��&5D�`,Q�0��chx���w5�?�������"!��fA�{��ߛ�P_z����`_������\�Hta1�Ky��|a@Yٔ��JRC/������13u�&�(�+�uPĊ�����,���6��U�2�L�T}n����cԆwXlU�:Gi�{-����D&Ř�X���s\S���FOQ�=cJ�f3��O%>����T"��>lf�R��F���.3�Wۋ�k�06��S21�����TE��S�1�jz'���4�Q�"�B�
���<��g��C����}���9�w������ �B!���L�q�^�j6����\8�s3�d�Z�{��.	Ȓ��m�����^�Jk���wY8����6���-x-��֢�d����΍�U�1X�3�dV����nږLQ����ܓ�2����fv�`,���P������3Y�;ꦴ3���dʯ��z0��S��ɦ�ߓ��|�r�/������Bd����8�q׍b��1l����ym�m�`Fz�ۓ1Zk~)���05���.�������=>�ss� ���¹���Ϲ���(�\��dzsS'+oڼ��:c{��+`��eFw~�{��4�7D�ƽJ�r�&bAK$d,��JT+�u�{Y��=4�:�z�c{��Z2n����Q���T�k��LV�ڃFv�����AA�.D�M�k� ����*��=dbטۇFW!�7���bߡ<��&E)B!��\���}����u�n��3���{+��i7>x�����1��=GςB!��Oʇs���ۀ�GQ�;���B�d&wI@���nS+L+j��0,Q8V��Nh��uAXfAY��m_��&��v��}��,��RT���P��b3��k3��OnX����5E(�d��j{�P,�Z�i��6kphZ���������<!�S��V��[�c�Xճ�xxǇ�*;�:�&��?���-bf~	'��^��Ss8vv�N����J�5i4�7�գ�t�.�:�'n�EkG1T��q��V��I�'B�S�������#�ǁӘ[�BH��$5�S1��c��"\�!���pa����aKez�km�fw��]ix�	RRӻG��Z~�J�.��4����"aKvW�j���� �Ldb�����zc{�J*@�Ũ��]����mJjl�'-D1�+�T�vs��q\��N�p�kf�kFB!���ǧ*!�����B!�BH��ȕ�t�j-vMfp�x��Ә�'��-1�'�<���~�{�>TL��B�cnxW��eF��L�Q�u}��&��FUC�jf�5�vhcf�^�r����ݿvx��`��[7����:�A�0r�0B0V0�}`p��I��Ã�r�g9��Y?$��?��4��i�n��;7���k� [~�51�_9�����E�?y������O��Cgq��,H2��� ��\�s��x��x-6�-�������Z[9�L{�M�{�����x���c����犸�`�|Ջ��<mcz/`~�$r��\��������e#\)M�A㻯-�Ԡ2�;��-��Zntw��}ɧ.�ڣ��M�4�f��EmI	Vb�r%ik���E&v�}H|��I�>1�#^I��Q���hWR���:�j�bj��X
�:��"!�B!�B!��nd��B�p�Vc�u�t����fΝ���D�0��=�V3�7���&�c�j�~3��6(�O>�=ʽM�M�9�z`�9I�
u�Qj����Ѽrj�mk��6QV��.6�B��E�n�I��M�����A~`5;׃=�r����޾���B�_�;׏ᚋ���'��%[&�ͤ��c�ɦq�Ʊ��]Ti;7������>v��>Y�'Ѡ�="�ϸd#�}�f<m���?�v�y��~���O��B���1|���+�<��M���f����ރ��^�e���l蹀�󧰰� �D���he*V����߰�Ml�S����CFw�hezV]G���n;&)L�,՘VT�s�O�Yeh�Nac�8�AlbW'���Cfw�%�d��&���0����(��;[�3��K������#�B!�B!���88](��*l^5��Lѷ4���)��]V#���5���FwQ�P��r�8ؘ�eFwy�����F���]�n��J���e�Q녪>��=x���fv���Ԏ�Y=hf��	C�C} ��NhSC4Ik�������\���f����	!�=q~�:��_�Y�n���~�+cC}���͕��}���S���W<���/��C���������W_�k/^߶�v��=��+�V���\������cG��2!��Y̗�f�Lj3��&���y�,Ma��tE�Ɉ�(���R��1��S��	�"1Kjl�E�;�yU�
l/4�7�+W!�J�fs	Y�>յm�I�͘����U�Lĩ`[T3�x����8�(QJgb��GQ6���M�Q*�!2�����A�����|?�?Z��ch/�B!�B!�B!���|�p���.�(a�0��sN�{�W+�d���~��=��=X?T�E�w��]w ^�{�Ψ^(���񪳹�=ʽ�M�n��
�������+*���X�Zb��$KQGT��XI��uDU8�&���M`6�
��u�\s;!��/'�*��7]�kW��p^{9	���k/x
9xw|�𾘣�C������Q�F��o#=x�5�+��G������W<�oBȊ�P~S���|�p�ƱfhOY��dzΝ��RQiv�z�L�*�*���4�*Y���^�����yϦ}b��:(0�����6��L��^ӹ�^�'�V���mz#�(�]-Fy�.�ٽ"Z}�A�)	�{��+:9��Iu��ڇW�B�w�g��Jǝ��!�B!�B!���5���zGq����. 7��	:���n��nW+Tރ�((+�����ʕE}���n�e[lg�{Ts��OdX�]����EuD��]V��{�EE�Pdh������^�4�G�
�S{OoW�ƙ��;Z��)�kƝ�	!��D}�%��s�n�;��w��t���)�&+�{�Sq��������S3 bhpW�y�0^���xo���p��1��%W�-�
�� >��Ǹ!dEqj��{�9W���n�e��:����i,�ϋ��&"�+,Y
X�fw����R��bUX��o\��^iX@<Ѫ:_צ���ٴ��%GC3*)�K�6ս͵�,j��nh��Ae��(���b�F�j��=���
��'ë&1��C'S8q��ω���;��B!�B!�B!�dn��	:�Lj�o'���iy����R��^/����~ӻ�(2��{�x��r��nۧ��c���hr�5��k��uD}Qox����=u@O�0\W��Ek��M�jC���!c���><2���$����cy�O9_9��B:���,n�|3^q��e�0����,^��x�;��ޓ��w�໏�xr�����~�<���Za!��e��ċ�������o<���EB�Jb!�w$���)�X�K��T���y�N�Ep{Ba��J�
W&��M���]D�@JCX�
��������
R���8�uc��>8^5.ܯc���jI3��l7����'��Į>����u��&4�������dr��^*����(Jc8t��!��(b�!�B!�B!��8����NUt{��=�f����N���Y^?T�	E���
�ҙ�m녺Zbr�j��>���qofn�^�c���uA�����v���j�g�Za�����nXO���02>���*��dG��;<s�gBHg�ߛ�Kj'^y�0:؋���⪝k+Ǐ�Ň��#ܷ�H�=l�Ư�t	�u٦��� *�=���]x�5�+� |��af>BYi�J)��5���1\�6�-9���a��4���-�"V*lv��X�"�0�]��0�#�'4�{���
V���н�����o��)�_{��[��6��ɡ��c�}zs{p��ϟ�P���E'wl��afكb����1���-�p��t�Ts{P��R!J�_KX���l8�A<|*�c��t�#�B!�B!�BZ�w'�ޭx�,��/ �0;3c��nb|�mM�~�{�@�@�PT�E)�vY�구.������}��ă�*-�1��R�킱Bf��C�aX�Zb����n['�bnW�ڣ�bUR�GGP����><x���s���=!���ɦ+)�y�16ԇ�Γ�L�}ox>p�t�#���thpGuk�W�pq����!�z2x�3�����"|���/|w
E�@Y��犸�H����Ć'�IcM���Oaaa!$b�j��R�r�����njt�U���av���'j������@�L[���^�n��Za����?V&h����{��]|��j��5m!�/@����$�uƚ�m��&"�N��m'�����c�ό���,=�C���b!�B!�B!��.�-���CNM�|�ƚ��x�Dk��͜�
e!X���, +n V4��:ˬV(	��d낦aX"�{cL�O��oS��Z���X��`��?.z0���kV����cIk��:���hr���I�ۍ�6�X�=�P��N��a��B��랴o��˱qb��S���_�����c��7�� Ǧ�RY�w���چ7?�)X�¶6�ed�����W_�����%B!����ί�Lj#��&��9�g0;=U~#�lQ�7���Fw�uRF���U@�
���Mg�P�B�=`x��i�aa˗����}��{Y[m��R)�ar#{h����+�"Su���~�5���New��⓻���.����o��m��Q�^1����v�����02:�|�(����y�ܿ'G�JR�$�B!�B!�BH3��
��غ*�'���
�?{��Vy���-Y�{e/�w	a��B��R�h���Bi��Z��(�m)�z[n�C�-���=BȀ �vl�{H���#ǉlK�lI�����p�y�<r�ǒ�<_�N��6���=R���s�0Q�=��a*k�Z��Za�����q��kzI�����>������m}�������-Y5���K-���| Űz��'X?���3��(�.=�S)�����@�-�5��X[j��U���84�.p�7VΗ��}[2�LL,����Vy��-����p/�ˑkV.�����_��/>F��~������� @����M5AeS��b6�ej�Y�z"∶K{�>	:�޻&�����8N|��P��米�]�w�1�%'�R�K\�=Q�=�~��{�?�y��TnK]|��m-�<����=ں��S��O4%��
��������CކZ�=��dS_A�>�������J��}A�l��Hî�|        ;��ʦ��<N�XdTN��M���(C?a���Á�jtҚ��WO~����6~�Y�Gؽ�}
����#�<̞��`*wMdOt�h���������� �I��Y?�c=�`�}��}�r�����h
��z�!�ܹ�yd��&�C�ѭ( LF��\2I�|�L�[M��X-&�`�4�̜��'ߕ�>���d���_W-�,�8Sl~PC}O�7V�O,��?�����Z  ����XR6��.&�(��o��ިx��k��`GG�2���{'�'��5	5�
��{�<�u�����Uj�/���}�u�%>N~��(N�;�S{!ѭ�g��	O�	N{�;R
��?�`:�:�P{�ɦ��u������6U�Ď�;5�`{J����d�	���"ǭ�s�&`���#���hg2
       �C�?$���ȍQ���i͗�E&)w��i����غJ°{_A�T�x��t�v��N��=�x}��5Ã�ۺ_\�=�5������L"�D�n���7A��h������{��P(+>��|1q��ۺ� ��Z�&�Ǉ�5X;LV���46���(��ФU���E2�,W08�
\򳋎��^�&w��}	��j�#*���ɷV-�%SKCW�˭_X&ϼ�]���z�� �\8j����ʦ�uާ�e�7,NiK������L,�O\%���#���D�P'�Tڄ��;�Mb%�wݯ�4�m}8��<���a����6$���&	��ݒ�-�� nB�`{��	���N��C뉂�]������M�ɩ�����ړLJu�7~S?�����䖪6�l�I���;D�       ���-���t���nv��"��r��n����ؚC�Za�uB��c��^�U�]��m��cG���ܧP$+�~��$X/�uҽhV���}��ِ� V�A϶�����>
`�O� �ą���[G�8��놩Vp�V�s�p����k���ϑ�啈�#�|��:$~���[����+�R�Z��sg.�(&�-��)[+�P7b��w�,��&Ў�"�b�x�>:O~���ew]�  RV�a�e_P��3���K��$��)��l�����@J!�>����hKGeU*�}�':Nm����7$������{�(ڐ@*�U�>��I��G�8?\Ov�;��T'���5	��]�ɪ�ǉ�����s�N�9s�M�٭i3�5a	�G�w��        }S+��[�wcg.���2��$��a��[���A�@�����궦�O[:6�@�����?q��T���w�jH�=�h�u�h�ۺ�F��|��b*{=����-�:a��Þ��Yr�y�3�dO�I6XCT��`���X��5�d�a����"������~ ��������K��:L�|���/�H���^�󫟑�=����q�  goKX��#�=�+�W+4�XOD◈�EZ[�c���Ǉ��	��tO%���p[϶����{����J������$>,��~��{��֨��gx=���SZ'���s�)Q�`&�������or����
��O@�:��l���A���f�؝�Xe���E6�F����rO��        ����n�wu�5��\�\s@��Vikn��a�8V�����5О��a����W[l�y�Gہ����zvo�}��:LL)���`K��R*����~`1A[*k��Ǚ\7Li1��a�}|��۝.�i����&�l��HxE� �lS�s���K�4/G��Q�8u���/?�m��r(:��96�\w��tZ� �����s���{~���ܦ�A; ��#"kBʦ�Y��@J��2�k�B�Z�U|�M
�zOd%���U���ڵ��0� {���P�Γ���x�~�0�޳-Qp=�q�!���2A��-��3Ğ`"�@���`{�I���(�{�r{$bsKc�&�Չ��H]׳�D        Ȍ�MaeS�L��rZs���:;�c�����=��X���n8��{϶���Ֆh�_[��Άnߓ�`|�����H�z��5%.���8�uî�@�S9J�=�:b�������b����Εc��̲�6*�{��� �I����g���$H��sF���\��W���M5�l���㐛�_�42G�E���ɘ"���ț� h�{�wwl+u�d�� ֐�"��I{[���='�MZ�0qeL�&C�':�~0�}���>���ݓ��S���٦U����DP݂��ݖ �?��m�ǤTgev�8\�Z��.V�i3ʦڰt4v=/��'\       ������I-�U"��L�X:�j_K��B݋cůfr�0հ{_����6���:a���E�k�}���n��-��YOLV+�zb� {�uD�8�^��s�>h��D*k�����g��X O}����r�����}�P��^�\nx�5ٰc�Jɀ��R���eR��㘙���m����� ���л*'��9Jd|��@���EZ[Z�OX�q�k�*���@'�DR
��w<�}m��'k�z�dP��j��| !�T���4���V�9ի��`{l��"��Dm.iYeg�ȶ���뺞��PY        7��!eS��J�	�cE��h�֖��k����ɂ�����ZO�*�ߞ�8�����O�8�y��D��_�k�];��8پ�x0����!�!�8V�:a�`{���0�ͮVf�H؜s`���D뺾g���/f�Q��j��0o� ;<9V��EG�-��)/n�#��C.�>ut������
�k�������w�Ij�} Ȭ_$�uR��c+��f)���i�9�_{�t�}�'�����$U�aw��m=�Ed����z':O֖�m��k�j0���㡆�S��u/}OLI���&�������X�bW���M�}&���ڦ��:��       ���{q,{l�u˄\Á�Xa_����ű$y�} �CY3Lp�/�>�uC-���\3T�s�0�x�놉�h�'��k]1ɚa�0{4fw�s�Ø#u�|T�����îc�@*,f����r��rAvY���9G��O�#ϼ�]�T�}��b��%����?�����`�/j
þP$��D[B�H�����$�٘k1�s�c��b�x�E^�2��wc��򋋏�o�ϋR��. ��j��;���g���+��:L2�m�gT���X�>	�����&�?ލ�&�zNf�:1�j�]$��{|{W[��z�w�$��S�$���b��g[*�Pݎ{���%���'�"�BOj���p����X�!`�]MQٵ/�ܧ��BUv         U�/,��M�Y�e-�q�F)sE�m
�9엠�E|����k�n�a�u�������s�輿v-�c�0�x�����}�t�0ٕ��%v�#��9�1�]2:�)l��v�lkI[���5]� ��`(Ԝ�.X*s'�p���Ե�C�M�F_G�)��i���Ñhk8m����f��e2��V��e1�^�-�؛�t�-����Q�
�Y�@lf�<��'2��$x
N.���[*V�I�����^Ӳs_�����ۑp䅊����`����~��B����1N�uA�ǱpR��Xy���Qy�S~��c��������@��	�F���ؙ�V��r�%2!�$Ŏ�䘂b��%�K{kKlr�8�J=��Ez��y�&2��+�*2�r{�dRIo�?����q���T�DS*ǉ&�����Y	'��`��s�ɖ#a�MڣV��ewsT������5��_�  @���f)�Zēc��(&���:BQ�D��-${�����\�IJs-��1��j�����3��QeklI�2F[����$ϥ���ƨIlfe���1�T�hD���J��+t'�-!c��5,{��z^G �ε"��F��3��3Gl�(�����r�Ar�!�E��h�֖�ߓ�5\7�-�%�>\��q�%kK����~��d�d�4���a?k�Z�Jh�����՝��i[��g��ui�uug�� Zʱ��'%3����^��TYߺ��5�v[G�s�����W5��k��iv����eq�˶hl�kJi��":��
r�isc��~i�g�D�}��B�Ig�v�:��{��4�^nl������?Pq�_�=��QC��=��:֖�6*7�h��q��!�}��ƽ�Km�O  �C�?"�Vu��_M����%ϡNj�@9��C␀D���oo�`G��dS�Ė���`�I���$�K����Ie/7qߖ�8�y��$�H��z��������������6��<��T�ۺ&�ԉOu��bWC�v�P~=m���%*����O*� p�Pm�Rf��csd��L(��M��/4�4?����]>yw[��k
�cb�Mf�ct�C&���a;?uя_X�V���>ٰ�M*�z2I���9�������:�#�u��=,Uu�����]�2FuC}�W_;g��|U_S���4M���M���{�{}Mc  �pT>�+[W�=�9,E21�(��%��(�߄|���;|Ov%h��&���*�5��{W[�}�����o�;��O��DfВ��`O�n�3���z�t_7�/�>�`{��]�="6{�؝959�C,�4Iu��*����� �f��|�R݅�wֶ�+����:�hln��m�:w������5[��������;:<�麸�k?~��	n�~&�.9y��ay�Oe���i��c?,6���_�>�ll�����:��]�bo&�����\w���Jr�S�sOS�rH�����O/:J���il� �����Ķ����\)r�b��|GD����s4(��_:�>e�Ht�>./�W���z�w{�}?Ǳ]��dmɨ��J
�&��(�j�=�C��>���{lf�Y����v�m������7J�Zͬ9,ц��� �P�Vi?~�W���B����2�"�S\���/VV���MM���V	�S��s;L�9����<�^�8��X0����B�to����Y^��"� �٠V����in)e�Ʈ��h�+�]��\������8y��J��剽�{���������}�8���1ڬ�׷Į�  0��������<b5��:MR�4H�-"nSPLa���������h8�OR+Y�=��¤�����%�'�s�4+�/�uÞ�IlOe��W��}��)����Y�]=�Z-bw�%juJG�� V�2l�7���������D ���(7��T�N(=��������-���ʵ�g��|�9o*;u�����]��o���\<�<o\�v���|���������hX�$�*p�-,�=����-��{��>W�����Vn�b�{��L�����<{t��{�'ϵ[��m[�V�gG�տ{A:�\� U�m��v�y��~�*O���(�Y��\�������K$�!Ae����'��WzIp��T�����R�}�yl�����N��z�������;����j?p[�@��sױ�b��!&�U���$�|}���R���ְ4w��rS��/8�* 0y�r��|9z�[L&��Q��6���,-�g�i�g�7I��[F�68cQ�,����1��Z�ybi����ѿ���|�3!�e��ϗ�f���h2���m͑����(c���{Fx̲R���t�����������m͑���{=�   ��@HdgSXٺZ�P�+�Y���;D�֨�L�� |���������',��J�]�n�(����}�ǵ8��(�������
�S�'YK�3ܞ�PVך�2 �*�&�C"&���f�M��Xu��T�F$ج��nuv	��ިos�Y�P�R�կC-D�~[��5Ϳ
O���sO�śF�E���7��7��R�����
֌*pٳ�5�W��֪����7>�h�nMۀ�'�*?��H�:mY�j�}��?����֋o�fm��؍��|D�=����<���w��c\���M�'7�s�\��W� �@~�W�O�{�~��Z�ڿu�s� � n���AxsD,�Nx��	H4�p�#V�A�Iz�c��G���e{�����v���Q��rOi��B
�L&�����&��l����%(Fi��C�%��ף�Ҕ(�^  #��(r��\�ܑb#4�2���y��	s�����{���a2�y^9{I�8l��r���FY�4_N�㕇^��De�/-���^}�s�
�$�u���\����z�_{d��-��T����9�PN��'���1
  yj�}[}H�uk�*�匝yl)v�(� KT즰X�1FC	$���U�Pq��*���|[l�ߓ����?���n8���Ű��\W���v1[�b4�$b4(���a�}��T�FzT`�" 7~f�?wL�?���O�}�qe�7_���c�]y�ewAEE�ֱO�p昂oL,��$�9��?�X������Q��ap���S����ml��q���v�~お��2��|ٚ��������R�����KNp;�_a^2�T.��l՞bR  U�IDAT��o �d|eKtKׄ�Aꤗ�n��(9��8,"sT����e�I�e� !�F�$K(�����Z�H��S�����&��'�dT��������:p�ߍ��4��h4vN"){��"�Y��D&�o�l��F	��V��HkG$Zo�+�KT��}5��  @jFX��2J�cpJ����e���fy`]-^5V�(c�D&�f�xʰ�V����9|�K��g���Y�֒���JeBq���w���1:�S�S�h{��j�<O�e2�����R�Π��9��?�U�/�{=  �ԫ7w����V��-�@�Z +_�ԵA�%*9��������DC!	���!	�u���������.}ȒԊb%]74 ��d�0��^!�~�{����:6�Lb�Z�d���d��5F	�Y:�Fi�%h�F�{U׶�J�	sr� ����c���Ӳ���pD���v��*�z�k2�TT�	������=uݬ1��5�����בc3��,�+�\'u-�'�<,�W��#��f�q����������W��,�؏.?}��;��w?4il^ޣGL+�k4d6�f����Y��� `��&��O���o��}��GtZ�b7D-:�Ĩ�=�ay�r`6E�}T�qT��m2t_ 7�)n�)�-6�Y����j#Q����n�	D�����*����JiD%��զ�Պ��`������9��*  ��Q������J�vM;�#�K�r��{��! ���r�)%�"�&Nr�-珑_>U%�j:C�h�S.;����9b�+�A�ە1�s��ZX2�%_9����9r�2FK����=u�Q  ��t�J�._ �}��f6����wYE&�r7�)[�Se%,�HH�:Z4��Q#�	c�C��D"j�,�
ս��������MZ+yQ,��X�hP`�cՍfuo���iPW,1�%��R�`E�W���z�f���kT�:±J��Q F��e�r��Yy�U���}Z{ፗ�~R�����[��-����/��5��^�5�kE�T��$V�=���.�~��1r���v�U��f͏�X��Bn���O�ݼ�y��œJ�W�vf��q�|�to�l�^�>  ��I�@H�_��J�<  �0s�\���B1�mהZ	��猒�=Q%[��Ou=:z�;�T/�	���r������+뷷	�e�^��\��"?8g���齲aG�`�N��/W�{������u��'���J�   @��Ԇ�R�����/������j�� j&M-������n�Rh3�����u����{��tDcű�����I�u @������%b5g��Ac[G��-{�k߾��+�#���k/>�o�����Z\�d�S��/��2[~��2�����|s�>f�����w��{��Na7^��V�����J=zF��Sf^����?�X.���#$     `�:��9�<Az8�&��Y���G+	�����Y��3Jc���F�}0N]�+������j��o�Q&�=UE�}��X�'�[V H��(�]].?}�R6�&�  �G�Օ�$���<  �u���Ii^NF����n���.?}��n���n��w=~�Q�K�+�w�2�ث�LR~�6��6w��(מ}xF?	�����͵����ޖ�������P��7c�K&wT�K�<m���ѷ     O'��n� 5�����r��{dgm� uK��	�g��d��N+�}�
��l�[�=�p{�Y����2���=|Xh����%ܞ�؇����?��5��    ��X�t�,>�4c�����~�o�{��W�q�e��x�/~f����O)���ǽ���yW�T7�Ȱ	�_r�,�T���cE�QymK���G���U����Z�=|����>����	�c2�'�+on�+�����B     @w�'8��	2#�j�Uɾ��]��ZX*&����	�g�U�,S��N�k檍��6�.�2F3F_}�2F��S����#~���Lqؔ����1��c�    ��_⑋O�����^��{ss���\���0�_��^�����{��Q�ح�u;mf���Er�}/H$*�5,��'˪��3�X���?�����/^u��`��**��k[���gf�>ݘ�����>_�o�'�-T�    `�(p�	efA��"��Dn{�J�:�|���(W�R�,��qٍ����Ç�H8� ��n��~V�F�h&ysLr�2Foyd��q�@}����hf�Lrթ%r�c��Q     �1f�A�]�H�fcFﭏ����޲�ƫW7���O�􆻞�˱3�-�ͱ���f�+�5˦��/m��}�]�!���yY$ml�<�ޮ�o�l՟RQaPK��q��<����/�Ŕ��s;,r効r�C�     .�l��o��� 1�r�q�<�nC� �?S,E^�O��&����������]|b�x��0}�CV,̕���kg���IŒ��>f�͑��y���6	     @&�=�0�\����zus���M'-؟U�n��̧����,�U���b�#ݏw��3�M�RY�&z��Ys�	U�J���4���oϩ#����Kg|7t��'����9�58v�(Y6�\^�\)     @ߖNu��1i�_C>T���q���ަ�v(�4�s�H���y�ڇ�R��6{\�,��ͦ�K
�Տ�d_sP�ۢI����=k���[ۤ�5$      �4��%7-��F��v���z���[������}r�/�8}t~A:�f1�7�\ ߺ�E]^-X��	%�X	�t�^��{������$t�WV���������aI�'�v�\y��j�X�    @�,f��wLZ�Ր��$k�̗���t�^��e�ʐH�l2�9G���O�tgT���
��jQ��Q�g�=�W���8���a3��er�?�      ���r�X-齒_(�����^t����n����_=31o�;�hT:k��"�̜1���]�7��_v�l1ӻ���-���=�n���M�>�xɪ?D�z��E��Lc%�"�C�9z�<��     ��Y�s�zji�8n�G�|�^�[)��I.]`d�.[d������LuIYcT�8�%��j�����;j�[
=A�9�-��V'�MTq     �qԌr�?�(���Vn�ݝ�n�_�U�6�]��D���m����t>�%'ϖ�7W�(�nW!�M/�E�K�������[�w�U��Su�e�����5+N�=�����ч����.Ս�     �E�Gp��\�>��OY�'��Op���z�V�?��\��3T�w��<�>���ϓ{�Y#��ܮX�/����i�kWl     �`6�+'�J��<�ޮ'�s��_�䑊��ѿxx��j�6�<ד��)��uY�Z�w�j�%�M�Ks{ ���=�n���Wr�WV�2灿���`�w�i�Ƴ�l�/�0Sn��     �e�8']u昙y��:	���qE6�Xb����.q�k���L.�Ǫ�C?��?��V|^GU�F9�<��z=Y6�->�O!�(     �֙K&��BWZ�ō��\��g
��k��{�|��f�<������(�_��&��}����8o��.H�K �g��~ɍ_=�i��|�����?�u��Z������1���[dgm�      �8j�[�/.�Q�ˑw?m0F��d2��).���fcT���,��71�:jz�
Ba�6�,���>j      �8�f��1S��o}\��f�IG��Uۿ{�Cǜ�`ҫ�.�)���V��������f�A�_>-���n��?U|���Cr�+>����-\8�xR:�W/���g�M�.     @�F����Q+dp�x
cT�'��^���魆��9��{L���:F	�     -�Z:Ir�����}�����/�����=���W�����^�r��{�FcZ�����/}$Ս�����p���o�m�;�����h�}���
�;���t���r_��5,|    �J���3s�C R�5K��"Пi�X%�p8*#YY�Ur�i)��!�>�+��CT���ig���e��@���1
     ��Vo?{ٔ������n�:��k���L-���3k��3��t�o6uVq��S��*�Nʭ9rr���iln�ްL��[����p��:b�c6���FeP�}���co     Ⱦ�	Q�U��,�^��4e$�>�1�WV�A&���J��d�G���c5����j:d$�6�1�W���ʷ�      �)ǉ''-��c��`ϝ7^��Y�f^���(�^W9{|Aq:�?y�X���7ICk��Hup_2�L����w0��l�}�O�:k�@S?����s��?~v������	s�����$��}     �ktA�&:1t����H��)LߥT1t�k�H��)`����B���:�o��(w     0T�W�� �[�?��O�B��G֮O����U�� ߭�e����x���ߛ%�tp?{Y�~X^�p�k7}����E۶_�Z��iS�rs��[����#&���(      ���-�*ϳ�>.�=�Q}+��C2�Q}+g�2Fu��Q     ��e3FIY�3-}7��#�ZO�ŭ_[��{�S�^�h�7����%��O/~$�`X�I7�1�.�3�(-}�k��>�ٶR�6��w=v��f�Q��OY8^~��&	E�     ���C�Mϊ�|
�<zV�e��\�W7�&Y��7�(     ���'���W���W��K�6߽茫'<���3��jݷ7�*G�(���g�[��Y���(Cz�~es��~���5�����O�=��7��^v��}�lr��rya�     ��j��vh����x��nM�$�0��7;���Q�c�    ��*�ˑy�S�zkUS��iW	�n�u�N)���b6i���E�	���&��8lZ�޼���{��N��w�=�roe�7G�S�#�    @���<�T=#�<ƨ�1F�1�s�g|Dlf^G�,��Q     0D+Mc*R�yo[�y7V"�������?�����9z��}ϝP$c�ܲ��E�E�%SKc%��F�]�	2�o�f����.���hJ���R��     �y&����H�h$��g|HF�<�6�ǨQ�뛌#�9�;3�!     `�\�	��S�����n�t�_�}�o����*w*w?g����&�]ܗ���~7l���K�m�\���wA�ǡ��R�ԏ�9J�              @�f�-�b�C�~C�����r� �~���5����玝5�D��>n��p�YLr��Ҵ��aU㵂�����ۧ�ᯏ�8o�Z��>v6w              ��:vVz
R��i�֛.?�eA�U5/j��r�̚^�ot�K&����U��Y�/>�TV�M;�ko�l�YѼ/piC�M�ˮ�e�O��R��               ��`9zf���F�Q����JAV��������o/;k�QZ�}�2^Fn�}JIZ��pO�����zUc��<s��1�iٯQy�=\3g�               �K�R�qh���u�n���
�foSۗ���Gv���E���_�$�p_���{e}k����K�U����E"����q'�              0 �KOA�O�#Ȫ�/[�u��޶`R�-��\�+n�Ե�%Ӳp�X�b���ټ��?����kk������WP�e�'��Ѡ^�B               Џ��4�S���1��n羦{L*�E�>��B���BQ���M,Ҽ�H4*��?����5��-�t;,�O�|T�(               H�b6ʌ�����yW���\zrP�u��c~^�⿩�m7i���	E#/�>sl��}~�����+׼.�����큫=9V����W@�              ��F��B�Z�����.�s���������勵�w�X�?��,ܵ�Ko�izB�W�m�ؿ>Z<�d����W(����                �t��Q����5dvu����se���}�*pI��&��IY�y�Mk��mw	t����e�m�=K�              Nf�!s����}����x����H�Ӧi��c
��͕�IY�O.�ռϪ�����8�M����wF�ѫ��f}���:m�Ԗ�O�               '�˴���k�xJ�+������?�x���N.󎜀��R��}�i�X�;7_�f��^�)t۵�w|�G�o�               ��[�؛�i��pD�C�	t�������@�>'�x$ӲpO�_v_��]�YۺyL�{��}N*%�              �������������^]#Н����y�]�����Z�}t�K�>�Z��
t����we�i�}L�[               �X:�{�[��ҍW�\���7�I�>�\b6%�H�d-�^���Ls{ r�Uk7	t��C�Uv�j�gi�S               �Xin��}���o	t���W_�qi՟� R�uHe}�dJV�n�E�6m����"Э͵/�a�Z4�@HZ^t              e��nD_�V}k�ne�Y�]��>��騼]���+ЭG*��t�+��6��TǑ� �
               z(�uh�_4����u�j��(��Z�Y��٢�Y	��95�8��l�ZCk�nt��k՟�l��Y�:B              ���]vM��k�n�ֹ���F�Tv�ײ�|���?Y	��s�������ZS{�Ne�Y�]�ɱp              H��qfw_��I�k�`�?Z��qh���KV��4TpB�t�#ޫu��U��               ��qٵ&����]�RݱQ�>=9# ��[4�3,F.w�s�`�Q�>3��              ���i����m��p�]�k�T�����bҬO�H��n��	��k��D���b6
               ��������6��u��ŤY�֖��w_�p75�8��oW	t-kp���              �dNC�2
�
t��=9V��٤}���Ǔ,���!u��]�uZ����              0�Y����Qi�^{ Rv���d� uV�&�+�G�Qy��"�@ע�日03��              ������e8,݋D�a-�3G@�=�hڟ�`���ϭ�zU�@��&s��}B���              B!m�*�����dԬz�*�~,�%+�t�%;��ReG�]��F)к�P8*               �.�����l�t�n5���/0��4|"�d6��-�2�!�3�              0�� ��h���0�u�=
K&e%���4�S�6t�l2�jݧ?��X              �ґ׵��N��٭&����:2���J����C�>QC�@�,�W�>�1�               �����C5��Y�6�)G�kW���|�Q�﹪�= ����{�/�y�v�q�@לV�x����              �p��H�ۮY^�%O�k��2��l	�tT�v;m3��粕iݧ��              ���B�Z܋s�Tp�9�ըy�}DTp���׼O��:N�k��G���:b��               @o��>�P�]|3�f6\��?Ϲ�k���f��u��8ʤ�ܫ�%���`Ь���P�[�����<�ͤe�{�               ��#k��1-Wv�u*7�6I�>�6�K&e%�
Gd_�_����T��W�[g�X�<$�S�w�A�4�2��              0��#k�[�V��V�u��.J�����J��jp�ZL���,���	tǛc[�u���Tp              H�*Y�����N��wO�G��Z������ɤ�ܷ�m���5�3/��y!�K�^�QZ����I               �X:���=��
_d��4�s{M�D��Q��W7k�gi~���TTD���)׺�O�j?�               {�Z�#-C�E^��{w<|ԏ�X��@W�<��Z�������Z�=�Ie��V�o��"�@7"eO��vL4j�g(��ʋ.               �D;+pO��i��N痔w�]���u��(jޟ�ܫ�$��Ԙ���tX͆����*��#Ѝ|��\���T�aQC�               Hnke����\�r��|�g��+v{��W?�����?�O����)�ؾ,�uel��8��ܰ}�               �ow��i�Oд�)��q�z�Sqթ�/�
,߱����E��=�iY��6��<�>cL��u��˗�YWq�GN*��j��Ɲ�              ��}��N�>������r�_][�>O�>7ﮗP8"��Հ�;�e����Y�q�M����rx� �
\����`�              �SY�&u-~)p�5�w|��!��<vش1y�Z��1�HEV��|R-���Q���肜˅��.6:����V�{�              @����FN�7V�>���+S�����H�U��Gf�Q�~���F�!��_P6望�c4�W�o�7���}�\�|g��z��<�U�~��Z-               H�Ukp����q�nR?'Ȫ)e��h�g{GH6���UjXY뀻�j6���V9\+Ț	�����7�              �L��F�"F����_��슇��T���⷏^<���Ժ�w?��P8"ِ����[�ʅ��м��
WW��⊵�����7��8wb�8��m�e�v
�              ����U�=Nۢ�%�9����?yD�jAV�_xK:�}uK�dK��W5���[�ִ�B���r��F9�P�qFy�04����ō�Y�4              �p���4��f�/���"�͊
����??mt^����"Qyi���^ظG�?n���ΟXt��~�̥����A�\�cK�M(������`�               ``^�X)W��'F���-t;֏}���5mT��i(H����X��l�E�}݆�i	���X�xj�^*Ș�ŞߙMF��mjȻ��               ���/�?�����5�{���oV�[wS���!AF�p��g��_�����!��up�^�,�w���1����tZ��߻㉛tř�i��;�`��������ww�.y               ����;;�p_�u~�Ύ���iWQ5����4Too���H6�"���[��p�uڌ�s�R�Ҫb�:������aQ=��v     �
t.�8@8V !=�S� cT�ᨘ��Q�
�G�U_B��QcT���      ŋ�*���êy�GN/�B�=��Rq��i���{+�MG��zo�t��0����Z���Sf��nѼ�#��λ���ι���	�ƹ����u���v�Ɏ�f     ٣��p��L�M�|Bo�@X\v�@���s�E7S����0*N��z���a     �����;e���5����z�T��滿}t�i������ �nf�}����i��Q+�/�R|Oźu�X�<$�ܵ���e�K?����     �����l�S{�2���t���pl��::���U?���A!��B     @O�񩜹tR,_��������'��KV�+H��Ş��KZ&�6��'[+%�tpW����e�Ii�����{�]�(�'	4UQ5N���:��7��oC���q�     ��m
�7���^�4e��i
��B�/�
m�4Q�V��y�_�ڨi�uT}�/t�j�q�     @���ʫ[�d��r��VC�GM/��;�z�o?���M������������>=��eucg���٣���1�F�������w/:���ɛ���f�]��������%�    @�U�er�]�O{�U)cT&	tjoC��t{�1:w�@�*2�U�d�h�@�*y�     y䥏�pW��X��E9+��w~���������zԲ��U^�R%z�����?�cg��t<��B�N+����}��7u퇂!���ǿ|����꿱�C���v     ���N����k�̝�P��Nƨ�c����<z���9     ��;�)[��W����L(s�����o~a�y�!���~���ʟ���ғnW���%�GAj�ܷV6ʋ���13G���|��4g|ɋ�֕W,_��p���w?4i��Qw��ƴ=Ɵ^�P���      }ؼ�'Ч���Ե2ݵicT���^M0s�.�@���ò��p�&��u��5��Z     �����&�ŗ�N[���u�w?�č��|D0$Kf�Z7���IW����ʳ����]�]��o��f��*����1�EMV���J���ΙP�v�ב�1T�◧��&     @?��tH�?,N�I�/�;5����> ��V��lQ�hD�_���)(���R��EvG���P��4��{��l��.      ZZ��V���F�O*NK�V�I��S�'�o�U�ճ^�O���#��.I�c�����$�.�۫����w�	�Ƥ�1�L-����y��z�`@ήx�z�伍Sʼ�t>���� ��    �5����mrܬ��� ��Q���[���#���k�����Ey}y�1��׿��EN��+���    @:��_����%M5�%�e71��?߿���7_z�'����'+N^0�2C��A�m�Ͳ��]�'�����̮�N��/��If�{�%�$���Z�RPauW_�(�e�(AX\��R�f@B�&�!!!���3��{�eqeW�����|>��ɄDN����s���N��䷸w/n�!�{��]w׵g|��/o������޻ޒ��.r�g�    ����r�{b�V4��U6�����eq�?�|��w���9��2x͓���k�YK���������1�,7�   ��7�xx��]J=r`�nF�xƅ�����Olޖs��������-���e����X��7���MO,�/~dB��#���#������~�}�o钛�v�C�i����RR�:    �ۂ�ձzs]�`Cv*�S�J�o���+�9?�$H��Wʣ��)xͪ�s袵51vX� O�\u�H_�d]m,]_����܌6x   ZHk,��mh��5�L�t��I���Vuo�+n=�#���}��M���_�/Nd���i�w�a�z��9�������^s����/����]�w}h�!�=������U1���,   �k��#�xnk|��!A��6c?0{{�FSgl�'"�����o4�٭qƉÂ��E��������k�7�������3
   ��l)���_��-z�	;�ܥ�ˊ��v�^�������W��gԕ�J�[tu{]CS\vϜHQҁ{���h�q��ע�.,(�c��K�o�gط��c�7�t��5ŏ�=d�Н[�\���{^
    mO/����C�m�Yۢ��1x�9˫l�NĴ������ы�*c���u��m��e���!x��+�w�-m��9e���k=   в����x��#b��-z��#��+-.\��7�'�⛧��༫�������'݊Zn���{x^��Z)J:pϼ�dc<0ky|���m��t��g��WN���5���t����9����ߥ��v0�5�w�}s�W   iklj�k������l�h�;f����\���s>3*
Zt�	o���)&O��o��0�~xC���Q-���7WY��<eF��lF����Y'�4�mh{Uc���   Z^��ϯ��|��_}���JK���b�%�}��'?���.�����-�niK�m�[�/�T%�g.�oN8fp���>t��}_Z�q��_r�a�q��,�N�Ko;�	C��ثU�\�zuC�3si    �C�!�مq��=�����6EM}S�-]_��߯e������ͱ��.��gɺ�xtnY|h��A۸�����&^Y]����&�
��Ol��Z��   @�X�jk>z>刱-~�A}J�>v�n^y��~��/�N����~Ȅ�6n�?ti�m�M��۞����HU��˪�����?x��_�>�>|@�Ž������z�U�	���ר/�V�*{Y*j��S^�o�   ڏ����=�[�]�����s�*�7wӓ�c܈��yP��u���2��=xs�?�17��cx��u�X\�.��]���=,7���ַ�gT����   К�~��8`��3�����Q\p�!�]8t���}jޚC���Ś�d���;������&�k���l�����=���q�S�Ƨ�*�ػ����w������m���M�ԥS�ǘ��)}��(},�dߚ����Y�a[U    �KeMS\z�8�Sãk�V�N��k�G7o���9.�g}��QQRlF[˦���Z�������O?=*���ֲ~{}\u���ew
��=���E�f����RW=hF  ��W��?��\\��E���-~�lcy֬�[�v�eS?����0+:����sď{���/-���-�Ե��=����޻�=F�k��u-��g����=��'����sN?����ιjʷ�}�����l�uVw�X��Y   @��pMu����q��C����m�h���Xu��+�/�cM|��Q�B�WQ�ܶ&�#o��Mٌ���8��B���:�<:eMTՙѷk�������;��vB��V�LY���    �-��X���R��	���9���wh�3{]{��Uˎ�ZG^L}�巎�uP�;&�2�K+~����6~>yF4�����U��]r�����}8�����Z'��?p�}9����W~�3?ѡVf��?o�g���M9`��ݺ����Wn�=	�   �}{fAE�*���� �{*�j��o[���wf����F�o=D�ق�k��?���_T�;3wEU\���8��!aD[NenF9%7�[�wf֒ʸ����Z߂^�Hhul*3�   @ۺ���1nD�8�]Z휽J�
�>p��,6픳.���=퓷F2iRsA�.w_vĄ�_��[[�܍M�񳛟�Me5����=�q{u���/��U��/,(��a���U���z��t����w��+)�����Tڭ��+���6~zӳ�   �����GUMS|��C��Uߒ�6no�����[����3+��ා%���m{Uc\x��X��6xw��R��M����B3��e[��{]�ь�[��-�=�6���RdFw�����gwu    H�o�����=F�k��޷��C��2�O���pS���v��h�~|����?f�e�ٹg[�������e���hw�{f֒��܃����m�s�SRt�������i��«��׿��[N9�1ڑ�\O�L��3�������7��o,�   ����̲��8��!ѫ�k�c�_U��{]> �ɶd��ϫ�[�����ۣIZ��6~}׺ذ�����W+s3�&N?vH�iFw�W��įsϣ����\\��ڌ��aFw��k^{��R�   HG���ᙸ��#c`��z��n��O~����w���+�U~�?�8e^�3�]s��F�y�����ui�[#�?kE�:}q�'����)ϼ����O6�Mο��>���۫7W�:�ڻ�0o��o];�I��?�������}G���=���'�����B�]�9   ��g�����+�G��#K�w��9b�-q��[�_�cd��nX_���8pt������{h�����M��hHw�,t��������W3�^d3z߬mqӴ��hFw����s��+��G��w.޽lF�z~[�2}s�6�    ����i�}0ztk�츴[a���Ě�/�1���K�V}��o��|$������C��d��i�?�����_�������C�����ٟaĀ��s�W3�K����u���=��O���4���`��SG��y��;�{ri�{��������v�   �Md�G~��8b|�����ޥ���SK���5�l�%�j����1.�cm�[����^����6�fk}\���l+>;^yuc\t�k3��#�����|cm\�Ȧ��x�]Eοm�k3��A�8�.,]���G7��I�O   �e��ܛ���}�(,h��{qa:~���m�����^�������M:픊H�/������~:vdߏ�4�W�o����~|������M�~����9Ν<#~�����1����2�OI���<<���V�xmٽ��T�{޷?�R[�y~r��c�.>s�Q�6���H��O.�   @Ǘm$}r^y���2>��8j�>ѣ������T�?�%f,��iY�r�9oeU|d�>q́}�o�v��i�X��>�xnkL�_n�p+�ft����h�9����`�mX��.?��s3jD[^6��������7�޿O�*1�oe���Z�^�   h?f,Z�:3~p��(h�U�E�]c�]��?(�����[��zK�%s��^wˤS�Z���o��>jpi���:��?��`A�6�C��zsE|��iQY��Q������)~|������20R���>=s�ɹ/O�ȴ�K7�-ް��ʆ���=�S�Z��U��u�?�������c��>3��%q��s   �\*k�⶧�Ľ�o�����������J"����PW�3_��'�ŜUb�VV�������x`��8t����b��R3�W�cֲ��.Z�ͪh�u��7ŝ�m��gm�����#���q#<��������,��<ں�k�b�[���f�W~F��݌���܌f�M�����(   �>=���(*,�3N: R�{����}r_^yL}������[*��\^{c�u'�8iR����;O�߯w�{�7�σG�ӿ�kA�dcYu|��i�����90��ݨ�o̯�?�s��^;���SR�;�������#{�vsYu��+r���U���64>��[ɲ+�v����wү���)�ۣ���K���YR<�_��Q����M1h�kw�\��5;   �Ϋ��9zi{�ػ(�ک$�U����Fׂ�#��d�j�ax�ژ��*��9�g��,�}b^y��ۣk�siL��蘡�bH���ڵ��hb�ݚ�hM�[Q/���_�B���^�[�?���{e3:�4F�ftp��(L�3��]��f��U�9��3�m-�`��9e�����{���k}I�64{��\3�}/�����h6����    �w���<����	m8�^Ե˸���玣s?=��z�u{�����k˫�U��=__W0��8��OX�f��I����yt��.{�ҳ{�޽K�wЫd�~����Tm�^g^�d��Z�Y�Q�;QYS߻nZ��_�F�e�zv��s?͎CrǗ_��Sg��u�͵��Uu���CqQ��®��
���U'�N_����m$   �_l*����fGY��Y�6�OQ�v�%�Qڭcp���E�5�QV��+��� ;�m���M�ّ�.�ػ0z�׌��f�}�]�7eٳ�*w�U5�g��yi�R�O�\�?2ٌf���1g�17�5u���^�[��h겿��_.���>��{t/��E�;��g4{��^ݘ��   �4����O��/�URT�kD�~�/�cB�8��_�̜9QQS�\S��T���P���Xڭ����k�nE݋��~��ެ�\g^3-�ok�q{�������OǏO����MvEG���E�u�{�=2?��;    �LCSĚ�����R������z3J��]�y��e��ٝ!    ���"j���:(����zv/�;�U��c��/��];-6��DGС�L]}c�}�3�c������Ô���b�*          :��箊�۫���}J���1k��8��������U����v���5;�l����wtI��TU�򳛟���          Ӽ�[����_|��9�gк".��|4d�t�!������X��<~x�?D������T�nz&��/          :�l!��^�X���1q쐠�565���7?�0:��g�-�_������c�������5q��3;�-          xseUu�?L�:b�������.]���=���ٟfĬW7DG���̆mU��?��o{�.��UW�W=07�<�j4w�;          �6di�Q|ن���'�>�������q��g�����:E����o��o!��[g�t@���=x�o(��n���n          :�g��/���8��!{޻����W⏏�M�`u�	�_7c�8�w��7��/��0<xws�[�/������          �m��q��O��w��|l��ѽ(xw��My!����E��3�Z��o|&7,����Š�%�ۗmk���Y�          �O٢�;f,����������sD����7����-������:e����_Ys�m��9.N<tLt	��������yqg�ɦ�=P          x���?���8|��8��cx���{l���9�~[UtF�:p�T���e�Ή��[���ǰ�����g������          �D��}Ƣu��C��?`��ѽ(x�Ek�ťwώ9�7Gg���׭�T?���1aT���G���w�]Sss<�����cU��          �V}CS���¸{��ġ�㓇����X7=� zqE45G�'p���g\�d>p����~�0t�6�?�Ҫ������          v��꺸��1��%������k�v�|Y�eq��⑗V�S��7	oӬ%�ǘa}�S���#��]�#��m��^X�L_�U          ��m��q��s��̏��%N>lL�[�����Y�6t�����-,^�-οuf\u����~;űw���{DG�pͶ�kƒxtΪ|�          �%�Wo{jq�����o��q��]�	ãkZN]QS��]S�y5^]�=���o�������-�=pŇ����*)��h���|��Ћ+b���          �����«�Ǡ>%����kD��7ڣ��Ƙ�h}<��ʘ��ڨoh
ޚ��jjn���?����w�s��-Y�=� �6oM��j�[          ���۫���䏑z����>4&�4 R^�^^]�/�O��6���vz���{����,X�?2�����20��=x���֦�5[*c����Ҳ��ܢ����&          �=Y���/�{���8`���w�A���b�!���K��Y�>喘�bs�\�>������D�-�P�?n��8���j�=F��݆��Y �[�s���[+�յ�b���X��,��[��          t��������#ӣ[a�5 ����C{�N{EQa�?����|��tCY�ǅ����]A��%poA��"�����g�E]ch��گG�S���޻�(z�v�n�_ˮ*���®�����M�M��u��+<ʪjc{U]l����۫c���TV���         �3��m������e��*���JcH���׳[�)��K��WIq��-.,���.�=�uu]�k�����khʷ�Y�����WǺ���~[U��iy�VVW�+6��          `�jn���옻|sо�          H��          �$�          H��          �$�          H��          �$�          H��          �$�          H��          �$�          H��          �$�          H��          �$�          HBᆩgw	    h'.���v����HPCCC����ۃN/7�����"=��8㌱A�w�E}?��/"=r3:.��rϣ�rϣgGb���g�y�    h16�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��۵c   �A����Q-�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,,�ъ\�    IEND�B`�PK
     )u�[����C   C   /   images/ba153158-cccd-4fb1-9320-38bebad1b7f9.png�PNG

   IHDR   d   4   |l��   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  �IDATx��|yx����=[2�=dOHB6H���Ȧ�
����R��jk{�t���zi۷������R�*b�V@TY!@����=��d��=�L&$di����I~�[���g��9Ϡ�Y�����b�x�Ǉ���'NwC�R�j.�s��u�B��Z�?q�'-jJj��c��c¡�v9�v�w,��G�O{5:L�	}xߋ�mgI34�o��RB��h-��%C����v��:as�q5��Q89O�2{{Z|؟����,{r��
�:6B�U������B̞1}�������N���*�Z��Mya�������\.}2��Á��V��P+ZL�o5M`�����3�)++3(o۾� ={�ɖ�j,tOrL�_�:��E�]�����������S�qy��Mʰ:7�-Σ	��my.�cA�	Ĭ��Q�Oar�e^�3<C��Y�e��w���k�5|���Pw-��X�'V翐�����mGOgZ�.��e����@�� B�@t�Q�֪eR6��f�賸au)}~\���e��^\���RM�����FNz2�:��i'���G���E+�AH �F�9D��59�X��5;e��DJ�V*����8~z�ɷ&'�{%8P�����V6w@�V*���j4t<5!6�ʖ^�4t�	Wx\HU� c�MN����H��BhH04�h��h�Z��׏��v�jơ�N�t�`�0|=0,�H�����c0(*�I�t@���p{!���1==�s�0-k<�b���@Q@���fC���ӭ�8^݂/��Q�a�٥5�"96�/k���7O�}s[��*��,�AV豿��������7�"�X[�������i!��T�wAI㓑7m*V,�A�ށ�GK�i%���p��Ac������D�.h�k�W�I����~�(��f�c�iț<������zss�`�utuu�HI����k���U���� �m���Q�D������*�
n��Wb�j�3�
��	hii��`�
!�������T���a���������CxsW��c��'�e�A�ų"`�*Fŧ�jZpOON�����W"V>/y�%!xx��#8�h)���D{{;��܌��^!:�����0aRRRI�187%%a��|��{��8��.�O��9��zΚ��-�I6���+������������ݻ�u�V�<yR�Ɏ�d�J�PZHFF�.]�U�V!++	I����k�?�8�����e�U�5Rg�w7Y�ƣ��	�"'#���?�>���
M&�yY�F�҅�����~I��r~pЌ#G�࣏>�W_}%��K��S	�������E��zsss1.:wݴy�����wa{�����I�ya0R¼x��B,_�� X�"�oߎW_}� 5�e��F=:G��Y,�8q���X�~=��<��Cb=�����"�����r�Pغ�f^��һ1))ڀK�C����}&|Yg@u�Opc#X��S7��{�,CHX�X;�?�	��n���3�*��+��y}�x���
Q�w�yG@�я~���Lg*��X$��ފGڅ���9���T<YƳ�Q��Y"q�������q�F�8�d�PrK� MVE���dF?i�iP����_��_�w���ϟ�I�&�?P��ڇ�]k�83g-2���Rf���$���g)�C.L�g�ñ�%y�B4�9ߣvS�䖟X���X)q�l6�7���/��Ʉ Zg�&�ؙ��
^/���t�J�`��[��o�>��7��ʕ+����_~�k�-��q6&�&�f���ibFSS~������iub��� L�LG�����F&Ǉ�h���@{[�O���|�V�Eyy9x����X�b2H{��ף�孨��H�c0��`4ۄy�"#)
��:8u�A+ٍ͋9�0c�x�t�CK|>6"�m��n��¼t4wP\݊�-2�G�����߂x�n�Y8��r��100�g�y���D��`�൦f�#�,��(��C`��Bz��q���vY�^�Ǐ�cqs=� b���Խˡ7��%6ӛ
�(f\+��������i30uz��G1�?%��9-@�]\,�f��T)�ع��� �F#�q����Ǵi����v<��ð�Ւf���z�"��ff�AO���!� ���us�VbޔT��eAv2��}�
'cJZJj�x`�l�,vܺx�\s��E��?�Q���o]���q��>��h7��C��&�!o�L�Q�~v��1�x ���D\�R���܂S�J`"p���{N�����GJ�<~�BԾ����HLF��G*��U� <"2;v/~0xL��M$���?�ȄU�O9����Y�/Qdm�������(!�_�BX���������n�K�Y�y�t2o/lD���l�l[��SR����퇫�EI
rRĪq�dQZa0�SSq����Z�;<XK�ha�9d^��5��ƙ4�	���� Afdgaz�,YӅT�����dM�QQ(:p]�bM,K&9�/F��<ܽ��o�aG|�y�z�Ǎ��fbJN���mۆM�6[��=u
M�-�����u ��i���iBPp%N��I#<����7^}�>�P��^HB(������=�P0W�jw���G���0g��N
�UL{�	�����ാs&���6��d塺@Y���:|t����Š�!�E����)QX4o�ģS�Nᥗ^b�H����s|5�`��
�u�'H�3���%2��x!����=��)S� �<����`��F�u��s�a@8�'�����>�'6,(�C�I���IS'K��+X�J�H۬V�\32�
$���<AC~ۋd���q;�|��K��c�	|7�p�fcav�QL�B};�,Y�6�-���pk5h�6�bs�����(�m��RJ�0�,�&�<��M[(����u�`�,C���f�x1��^{}}}$�-��ř��ȝn�:���!�ޡШ��{Y�V���B��OwJLe��Ĉ�����3SQ�I�0À���ɈFf��{׮]�Y[8�O�1]bSvO+�&8�%��vv��7�L>�4-��$��T,�����g���Ѽ6��P޲���֓� ���LEc��fsbDPf+9R�$����Ҙ���51|o߀e�^!I:̜�-��4~�Ν�r)S��|!*~ː�@8]kHl!�TС$r��x�?b\$&Q��x�����vYI�����{��c�Q}���B�<2����l��ux|�NԖՊ���\��`�X�� �W�J@#Ka��Қ3o.N/����~]]�$Ry�iH
/BC����$^�)J���tW94'���G�+Z׬�����?���az�������n��p�.X��;�e����jQ���Z	�LKANB�֛I�J l�Q:%rғ��B�؟2�<A~�
[�m�B�g���_�j����3y���db$��u��=zT ���AV\��p�5��C�ʃ܌DZ_ �/��R\1��#צ䎥�u1��3� �:>�aוH�My�S�$�˗/��w���}>�bB4�����\��:O��:�؂�'Iʔ��-�27���ޞ^�EF�ű��H21���Zy?+ ��MYc�WjpHP"5!F��K�O�<)w`e.���\�^��5)\^���K�Gme����Sl���'FQ���k��R�@}ȣ��U\	�I����Sc�p�e�����5(�
����v��V�K<A.Nr�NK~;n\���Tx�еJD���ߜk��b�j��Q��� W
�m���?}����}��a �{�A�/TK=����%�`���ݗ��QA���6��5�`.E(����X	t�@J��[׉����!-�r�w�}�af5�!����u��Ā��:8V���rrhw�`YBۆ�����-�@��O�Juق��:���pY��D����|_�0z� p9}�Kz��{����0 V
B,,h�����5ea-%��;i�<h|��XK�W�9�:����؛�{����8씧8�\���������/!��'��i�)��}���X9q1��N�P_�jw�)��Ff�qXOLL���o0צ���M�R��C��;)	�Sk~'�D�tW��p|%��D����c6L}�UV�v��a�U�*�4�r��^�N�db�M.ޚ-�=Oo�	z>��D��ϻMNt�(�NEzz:"�]q,��%ם8��=�)����b�F��Q¦PKi�=�շ����p�qM�,\��O6�=h�����ڒ(q�0V�F~���+>�
	̸��� ��2q����;?��w�."8��}p�)��B��Yݨi�cf�4����P6�EEF���q��#�&�G�'�����)��mX`���K��]�b���={�\�Mϭ�0�J��݃�is)P~�+Ic�����L���66 ��U��O%�����
�`W�J����A��FC*�{x����%��l�����cٲeؿ��.q.\ ~����,#-3�Cp�|��٘��.�x�:�a�:�;l�-s� ;;��@Em#�\���"�c�� &6Nji����F�]u8y	�q|��[Ɍ�uaP���rD��$���5��g���Ȁ�hjmC��$uAëf����Pd�p����E*��z=v~�V�^��d)D�R3ӥc&�+Ŷ��S���N>��gS���r
g����K��j1c��Z��\Y<�&V�6���:,��EAA�Ν+JȊT^r
�/
���J�Z��ű�<W9X�آ��J��bs��Sb�L�V�^����1v��
mnz�Y�E��6�����Id��3�>� ~��_I�ݻ{�⑛7��Cu����}Z#�`4�IBg�Х�D����<!+e��Ipsб`��N���{�;G5�.u\l�$nڦ�����;3O�G��?���Ue����c�C�x).(�P�������ix,�_�B+[���>�2��6l/��-QC���C��6��wO#3+w�y����U�-��$�͞�#����W��9Fh�>6�4�Y��Ox���C�슷�<���B���Al�u�F�9E�1�s=�� V�E�z��'۱�D��?Gv��{��K�PY�I!.ܐ��s"t.~��G^/ˢ��hnh����~&ۣ�7>���hTg��(��M��N6l;���(�췿���5������o���� �����~�Q�P=�'�A���ȧ)~�q�z֬Y"ރG����U4g��gh���k��i�F������T7wK�W��C���h7+�����JCTL,�|�I���ٳG@9q�X����dS��!~|p:QT���&���>�(n��f�7����]�{U���O� ��=Ԅ�̃X{�R��*6皚i��۵ՕU�6#_�V���=C�Tu�:�(^�46����@��׿���.�����K���::v�ă�CT��6�GZ�	Q����'���'�s��[��C� k�	ύ[�g��rf|�?�{�R���?����,�RGk�loGVN��Wt�[T@�(���O���N6=�e0�������\<����l�C��<��[������,B\T8
��A^^�~�mq/���İ�(���>��01��p�0P�����8@ԸG,�����yO[�ڵk��v=^ܰ���"�Q�F��I��w
{,r���zS'QgàPU7�E�E�D�t��}=s/2T�%��9<\�4�����<��|V��ؽX�l)�������f�͛7����?�*O�b%u�Q�E����k��$����o�y��`��!�¥eЄ�l܁��]R�:{��e�u��y����4�ysfc�ĉX�n� ��[o�����4�Y1BQFm��I�֬Y�'�xBr�yԞ_�16��WFvC\�	"vc���[G��99�������ơ��$J %%�|�ь� -��c��/�)��{_ɽ7^����b)LO�Cp��˙<����ԐG�[��pn�.�c�op��u?�+;��R��A�%��_�T�O��9�6�K
%���?�Nז-[�^__/%��2È�[/��-K���1�PQQ����������B�������;��/��~�_����za�!.2f��p�NO�����X	yK��y�K���ݶ�Z��p�s�=���k����QUU%���lο^�e����[n�E�8qŃ�b�{}�gX��	6������l�A�����QZ���+"%5E��2[`Z����R<�dq��� צ�<����38�I�~v(�+[�q���ۊ:ƻ���Ĩ0vj�x^;opX<=Av��� ��w�fwbRJ�����A��]a,���a��M�J�U�g6�@9=��51ib��0�w�}����K����if%c�c�p	�����j���'��������_���a@������_5�l��48�x���+����9�v�t$%&H �5�_$���|�� ��t�xi%���>/�ɥ�(z[�ԉ)�@	[��9��e��_Cy��ٽ���k �}/r)��˚?Nb̠��[�җ������݂�da�5��?$#<<LX!���-eT]�<��4�ʚz|��m�~з�y�9��^8�zd�λ��b�hQ!8�a��`��|/=�X�D�{%��]�ES1wj2SE����el#�V}'J���T3�6a�+d��X��c�E�/˛�*\�m%Ƽ�dG��J�|qEjE�r�d���dF�]�p��ε���PX9�����wV���X89��i������Hى��N�fqb�lFGW�j�e7塚��<�Ϯ<��c�u�J�@g���>���|7?����#!2hgC����R<�X]�(Px��0<���r���F\�I�:y8o�d����g���`���@�����[�NKV#9�E��`�-=�PJ��`j��A%v�:�r<�	� .�W<�8�M\���fŹ1>�Lא�����o�i��&��A��V��e��w�8�#tDE��0�[o���n�[j��x��Mf�iSR���-�NLJ���k��yǩ�>:� uTh �Z4���`Ɗ���<K�y��w�ԩ��D����~��a㲒��v��>3M|P�r�eu e�
�����H*q��Eh������]]������J5���Պ�+gG��Iy#=6 �fD�q?]�U	8F�ێ���]|%YV*&�����h����[���/?����K�&N�uw,�ؿ|IMs�|�����������j��AZM�[[v{fg���{7��o �H�_��,�T(��v����C�!\��\�s�s,a0�w��3x�3�Yj�(R~�C��/������"|H;[��7����gz�� 3;X�_��܇c#?i��~�����m�o����H+I�3�B�:m"�v����T+�7�"W��T�Y�(��}��A2��6#5bQ���+�g�صٝ�-mM��]��ܜ�����`���5��&���ge��>����-eM=A��4{�+�D���9{&��Ӷ�4J��:<^���N;~��YAnS�pzݬ��%>�ʀ�NE�t���*��m�C�V���xlN�W��f����֣�)�u=1##�a
A[�N�?q�&�+f�5��A�/��z=Qĸ�o~c���m�OuSN��F�w˺"˟c�U����������[�m�[�Z��
u��m}�0�@�b�k_Y��)5d8y�Փ�w�=/�s��~l�R��dl$��q7�G�����M��/�&D�vI�T���Q��؊�E��	
E��A�۫�X���w2�f��3m����h$P��� H�4��e�+K�.yF�sq�6�i���kv��q5���qa�e�;m�>zW����/3tJ����UM�Uc��s����+�A�fqZ ���tKcZ� 5 |���MF���P���__�%��q��ߎK�r��o��Ʒ�\e�[@�����lS��?�    IEND�B`�PK
     )u�[	��} } /   images/bbfae99c-8036-4c5e-89fd-a87441410720.png�PNG

   IHDR  �  �   ��ߊ   gAMA  ���a    cHRM  z&  ��  �   ��  u0  �`  :�  p��Q<   bKGD      �C�   	pHYs     ��   tIME�#Պ�  � IDATx���{�m[���Ƙs����8��GսU���袍�i�4��A�("�q�6'9�Dq��E�HEVd��HX�d���&�Н��g=��n�}����ךs��?Ɯs����{����f�J������k�5�x��p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8��}�𵂪 ʳwQʄRZ����k��{�Lǁ�%O�h	*T�J�`011@��#�QD
*B)�@ FI�"4"L�Db4��L[�>T	
4AU0����11��*��J���N�L� ��m��l@�(`\m.@aW��7W�G�|������%���<�Ç?���p8��h��@K�J���s�H��K���EFi��_j��R�kh�,A	P@	`   �jQb���!f(PA�U{�B8��W? � �FE}E��z�T�0b��P�t�>��1�yPr�P)[��7���I�����>P�+��T�hT ��ۻL���J��ui� ��5%Nd?#��z�vH
U�w�[��}��rV)R�""�%' ��f�v�U!�bs�!lJ���x�/.��Σ�~�S�����G����7 xD������%b~�]  A�=��~l�,!	"bz���
�*�E �
$S�
t�Nb�Z�L�WaEM����DՀ�Ĭ
�h�AU���!7�(���?��˯���1(��a��%�۽�����]���$���}i8���U�5�ժ��T�[T�GE�C-�J��eC�����	d�VE�RM��F���dQ�liO~M�?'0�w^d^�b�Op�x<��L�$����3x� T"��q���/@%B���w���w��ڄ����k��3o������k�q����:Eӯӳ� e�n|�Z��	U�M"�7h�Yr��((W���� D��@U�����y��䟽��� �6� ���X��D%"H�T�(�R��0+���	|KLO�x��8L����m.��>��m.@aa�]�%����P��/  �Sm/�J��eM�7h.�SD��J�$_+t�RM��
 ن^X�f��@�aJ��QS�t��k��纽o>c8y�l�BqĻx<������{MH��sF����J�v�������U�v�+��K�������]^\��^��������ԟ��|�^�/�-�p����; t�0�>]=����_.���FD�[%���P�)	R
b�K)PUÀq� ̦���2���_�+t�;������2{��W�~N�D�DF���k��q( �fB8�g���90��2�d�����q��o}a�X	�@�>�G�ᗍ�VU����n�./��'�����/%�n���Z�K*%��Pɦ�T d�ά��H��Du�Z�9��yeӕ�����}N�]�v�W-�~��;?��c|���	s)(���QJA�fB�C`036�`6q��F��,��j�@�.�q�}�_o��v�y�~���g��W~Ƌ��Ǉ��q�`ڿ�_�o~��-������<�Β�o�o��V�|����D2��\!���!F\]_#�(Q�W�Y7ƽ˧3]oqǕ�\`S���"ZM"�� J�jTM1+���y����M`��P���ϙ�gƟ��~�Ke�q�1^\!��1��,���;�������/b�]�����U��HI�Z2 ��"	���`^yۨ�j���l&��mH:��@��l�
^P]���u�{	@��9��s��{<��s�7��.���L@��i��%c��؍6���1b�<b�#��E�0�+l����U�_�������b|�_n���7^^���, "���~����g~�G_�2��W����O�����%�v��7�i��|8n��[���R@*��PJC��`�!9���E��^z�U쮯�(��RU����� p� )�z�5���5ki_2����&�5���5�Ye.1WEO�����9
�'����e~������3������1ݾ��}�������o����!����?��9�.��T��9���I�"')�
�慢�B{�g�Z{�^IU��mt�Y�8��ieٮ����$��qԮ�0Q���.~a�9|*���ÌL���9�((#cF�P��BDĆFly����.�<`Ѐ�p��Kx��|}��[����/�~���T�O@)������W�������~�ǿ��y��/a�yʘ��b�]���o�Ͼ��2r�~��p��3,����4�P) ./v�$ bLsƓ�^z��x�ʫ��
� "���ӅA<�t����<���])U��kH��Wy��P��]��� �r��G��C�U�/J?�!�(��#���,o�M���#���#��p}�����u�П���|�G�|���������e��_�|+��*�Z��BHU��(t�ͧg}	yK���*3
�U](y%@hM߯��@���a�y��`��s����N_�8�@IAA���`F �!�b�
��1�6<"P t�J@���p�勏��W�`xTv���8?I<��ƿ�H���4��.��C   �7��+��4�i�p�x�xx<D
�:�ߖ�߭i��A��8o���� � �3��Md�H���#��9g�./����g�N	�^~��������Č@=Q�z�I��;:_���LV6�^�l��H���_׾6	�<vQ q�P��@���Y���q�� �o�D7x�c����@�P���/�*��A_�����폐����_�^�����Ayz�� � �J�h�V���c��S�w�Vν~I5!�)t�j�/%]š� 뤸��P���x=@B"��%Ct��@Q2��j�H1�Z��JI#2fd8!% `@�� 	!d��������F��:��?����R/�t�{C�o���6=~��v��o�~�qw����AU�RP��Bd�p�:s)�ó�?V4��9�ߍi���p��·m)�I��{H:@JB �%�'H�(iF>�Q�H4(�>�@cA�	�M7�i��;()D �%oz����q�9t�:W�dg�o�;��#����u��I�%�X�a���|����(�߮y�#!���@o}���8~vs���[_�N
��~$�}�y��޲,� �Q*��9�%��kXӀ2A҄��4�z�P���oYY����aJ�E�*��j_�*�cYXk�PN��l-(/4;��.�S*7����S�����	��IZ
� H�H�.� K-��"
5�d0�6؅+\�x�W.���xix	�0"`Ѡa��4���g���e��2���x��p����-!����n��K�u����9��3 �����͗���o�*2��O�\~_��o���O�i��N��y"�3Ho�Z 2!�#JN`"��9!��r�0�nn )!��8D��r��E@q���5~�۰���FFV3#R0Yc���Q�.DW��ޛĉ�~��P3	j��6��*s{ͪ���O�u�y�T�����UM�0(�X
�'a:��C�i�ݏ�{|����Ȓp������/	_W��/}�!l>���(�Z��-��D'@Dg�(D$��I�\��%�-h�Ӿ_|�U�v7Zy��1o��B������״}��;��"�ܴMȋ�iT�b B$�j�,�JBT�[J�A�X���B� �غ �H ��`@)B�6(��3o��4��4 �	�kL�c�O��g���8�0��s�Ͱ�~i������w1lw��t-����@��m�$�9���M<|囯5��۫W?6�~�j���K���U��n�O!�-�dYfhI�r��-E��	I,^.9!oq�y
��0n�u����3�4�c��ͣ�-bܘ�#��a�K�J��J�S���$�U�ng9��޳�R_T�9�h�EƂ�@�����OՒ�J�I9D����)㯕0��D�ߺ�<�����~������������O|�ʬ����O�ւ�Z��!�㿡e�(�)G�r�j2[���T�<s��qن�R�T;�Ψ*t���F��9��z�Z&'銢jT�4*���-���9��ւ�Y�]D@PD
�H%�&����Q�VC��H*�b�#Ka�]"�Lϰ��pF��~ʀ(
�y�&��M��7s���Y���t��1�� ~!����g_�t�3�C ¸�Ї��43�3���/�ٳ=��
WWeh���u0����#��̀�rP@b-}�j%A���BH�L@mX����D���Iָ���Z�X�K���jZ����1�}��p�b��`@IJ�A��AT0� Ί�2f�vD���q����Q��0E�t�c���
����v���}����;�y�%��j`���A����o��I_�"��>z=ݾ��*�E�'E��Z�5D8���h�C��	�@��|DIGS� H.ȹ@0�	ДQ�#�t � C���05���uw��"_? �&[T$K||�7�ӄ@������u�{��KoΏ9\����%/D��=����f_tN��;EJ�֛R7J_#�@uF)�e��{�O�����~����~�w~�w�����V���u��o��|���W�|��K�H���"G�L�2�lJ�%ͫn��1F��Ϊ
��w�yL��M����E)��z�ž6^O�:��׾�aU �Z"@�lB��;��,O�@����z!�$(J��ށ ���l���p0R�Ť���3bQ\L��-�����A� ��RB�v������5���������3S��8��"z�oso!�o�?�O?���q(1��%��f�tv"�w��T�Բk�a � J�s�a�q���	L#�iF�G�M3�:Z2r���<�������}��ʟ���G�q���D��2LE��FG�b�c`��B���L��	, )�M��`bb��Y��I ��H�tr��7�>½�
�����_R�U�Fji����P��
U"����V!�K��R]
E� n�b#��:�Ah�t�����p!P �����^������ 8>y��h
n�S� xh+�Q
�60C�~a�.�J�s�JB��g�o��}�f�g��]4b��� )�����/�9^
�Hy@�!��H�q���7��oW�߂r|]U^*%_�f�P�W�Vb�%��@�y�e>"�(ǣy���-e���'@b��%c:� D�4�e����!�@nn��gL9B9X)Z) ��oN��%�T��G�ÛR&��!��Xe�$��nғ�A+��.R�m�e���Ξ-�K��%�i3 c)lT�D@��H��)�''�o.����nz���O��#���a_+|���f-�a�0o����5_)�R�Ũ'�H-+SA˃T]�oQ�a���g�8M�X�jU�X�6ֹ-���s��2�kѩ
Z)�wR��G�؅["D�Ь(�0A� 6A�(g(B��g��#B�dU*`Q����)^C�
�hA��43��A�!��A�^�^"���{�BxF����D�%����ox� �q����ՌF��� r�0��N����N3�W��z���y `_��"����.
D>����d�"ø9��IidC�qP�AJ� �1�C��n�	1��R؍X�S�4A ��(TsE��*7�\5s���C��L꒮oZP�7�7T�/IAbJ]�i*UΩ�Y�(DETUE��Q��q��THJ	�E��,Y@9�EU���PJ�&*��"���T�\��-�˂�-Ƃq,�~�_�9�B�R����٫Z��*���l��r�^�3=��C�<�������`�hH�޽P�E�#��HyՇy��\i�;���9�ΐ־Y�'ת
J� �(%[-�<��#��M	�fS�R ()4%d�ӌ4O��0#猔R�P#�b�R��0����f�� sg8툩9�M�5[���Kύ& ���K�{}��$ԭ����ԍ�ƪ��ηváv�_=]��p�b� �d�I�oU%��w�VDE�n��2��ܼ�i\����zV��*�ӻ�'{�q�M���/i�sH�G(gh��V�V2���>���@��L�QSƴl�N�t^~��۷}JQ{]/1��Q�&�v���^N� ���M^[�f��FR�`l8��#v�E�2CHl�Q��I�d���I�zp�`��DDe	 &&��Tn��u�b@s���\KE2�L��  03�Ja$#��� V�P�C��8&���(4�(QS&��L���U���(I��+���� ����k����v
�<;��T�i�����a���2���(��r�BsR��H�L��HDL̡*_��i`Bd!��͆i�/]1^}i
�U�K��q�u�V�����û��|Խ�6L+MD$���Ｔ}L_՚����R/n�7o+%Y6qVe) e0���([�DDC9BDTPP�([P�P	[`���P���VG��"�%�HI��R��Ǵ���V�!T�T�c֜7�������Z�̌�{5Z�v<UHUI�����V��b��*K� RX�0����b^}�P�*��g��S�Ħ�i�q	e>�oQ��d�Ϥ-�Rl��������
���cJ8���%��ْ�b b4�:M{H� �S�-iM�@cS���YS���3=]<4e�L��&��7��D]Q�2<f-��w�n.�~��G5�,"�mb%S� ����Cx5���k���n��4r�x��O��Z����~��C\~��雟�m�������'PI֛Xg@��=��F"�j��V��w~" O��~M��S4����z�}�,���歯�f͆��ڇ�d��fc5/{TƆ��BϬPeX�2��Q�D��p���� +#h@�!����!?E. �ƂѕD���huRTC��� �"�z��`G�� ��o�����Z�&�Qz�w��y��CUf�<eL���O�xrTd,�X2B����$b�:
�xf�<�3{�D*}K1�ĀAB���0!h��̀a�������D!�����жt����M޻��o�[}����F�,��'����ͻć��ď*A���Rt�-^V��$��%b�p��[HA<a�`� ���tܢ�K��щ�P��-!l*1AF��lbM����l�=Y���
{?�x�=Y��k�
h1o��Ĭυ4�C(�"E���T{OT�ԩf])tj��u{#I���|����) �֬�~��j��|D"R��<�8���8D���M�l"B$��ʼ� ��7S�(�i>�϶լ^�n�ﲹ�l]���{��*���F��* �:�et�볰<+2O�b芚���ĕ(�Q	Py���P��}������ȳ�O��)<x�[�aǇV��~����@���4���n��*�
��5Ͻy�B���4��*���{����z73׍ghq������K������������E1[���
2�P��  ���
��b,�F:� E�Rz�A+0p(��\`��y
(]Yk5����C#��jV��!�׃V�q���#�g*w�ξ(�/pW�j���1�$I @�3n�7�`�@����D�;WDP�@T0�	%[�b)&l+8�b76RT�	��U�h�\�	~'��}����N�25�6��~��	Z�"�	"]��l�
�{��)T��!@��t��i��#Xf��`�
@cy��4@C��-hs�v�n�p�{_�U=4�¼(��8�2�M�[S�XN?�m�(s�5	x.�5>�3��j�I�z�K���O�,=f�{���'��=@5�\�]q�P�#����JNV]R�0��V�V�3BP�t�����^_B&3��R�t ������ߢ��h��t%��2�O����T��^/�k �Tma��0�����?{�J�KM�CϷ��r�若�E�� ������������'���{�	�|�Sx��oy�g���R��޾�gሇ�UM���K:��G�̖"�f�Ve^�~	��!7�l�n[��%�ӂ�-J����ן�)z�+��O7�J�wLZ{Rj���5�X���ʜ �2�H
��N
S�\@�M�Aњ�7Ȥ"(�}ge5�t�@��r�1�A��`�8T��湒V:��}�*�%j�ΐ�E���m�"H���:��`�ύjڽ���D[̀�� �#O�,RD�l1gV�@��5r.�sF))���!R�e�0�-."a`���UjhדX�3���=(*x>V���-LY��u�� ��=�u4� pT&�NвM7
SX��0���vL3(O�<�'j���J�TD  <��:o �%�`�ov ���^rZ�U��Ր�5-mMZ�ЪL�p��Mq��g�n��[Bz��֥��m�h͏��_H}F�Xy�-��׽�O�}��)��a��$	��L77fP��
�����mă�s��2w�v�n��Q&���	6�U�!��o�N�Jj�u5��]�r���5[��ht�ʘj\���AlD���^�Q�2�~�*��~`�L3�j�Q���`���69W`{��$
�����O�G�+����`��e|X�S�
���ޔ|�'$�T�<hIF�kF��PG��r�V�V�̓v.+ֶ�Im���'V���wS�k�ܳ[�u�z�<��/[�]ey�)��ԪI�l���w&�v�@m��d0g(�*��%����6�%P�Q����4`�r�$3����л���ٵ��^&*�W�*ШUi��P�,lM�����Oj��w��(W�kJc�͆ ���Cf�"(U�81B��� �\��{�V0P�Zl��-×a��|Ļ���u��
H��O��T�C��]�rQ�͋�=����v��(��b�.�`���.��9�ƺrD��L��Ϫ	(
� �	�� %�����T "0,��T�2�)��!� V�._�� ���M�	b��GX6�+��:ٻ��5m�*��Z7�6���S�|��β(������h�Z={ċqQ=z�RKK�2��,Dl}�I��,N���9�!0(0r��b��#f�-V"I���`I��7�f���ۍ�<�?`:$�3dN����z��
�:٫��{�����5��x�M�wơ1w"+�[��`�G�����\�3���}4̌��OU�#֌�z�a	J�������9=���G���'�����q��gq�!m@�S�7��T���%����%�XӒ�e��l-=�]����+���f�����j��$��Ic�٬R:�컀&+D�F�¼��,����*�C5Fd@i�DA����2�b�'�f5+�Փ-( R$�FիoP��(2�5��Q��/#c/��2n�G�A���vo����Rf�;2\@� ���l�r�@�Ӣś����O�\ʲ2wj���k=1�B�l@R0b�u��	9<�f(P�le�2Z�p$F(&���d����Lur�Ֆ�R��
�12�����x0(X'�&�-���.���[����J	P�o�Jm�tU�띪�ꋵQz��-g�R�N_Dd���	:�V#���Wg��
��`L�,IrU�TD���*
���n!�-�b��PF 5�����B���O#�-�e	^�@lFT���<'�6N�5׵Z�ֈ��贌����3�L�Z�ZmHͣ�&�+����o�
o��vT((�e!OG�)a�8B�`�7�W�����O�<��֔��|�s�LG��"6q�V�K����YyY�nJ����^��:��*p���T���85�~�4�3�<�ET_������J *5�*˥�v3���k�$9�/!��O����ç�K/�>T
}z�H��'�|�Ki>|���:!�)	��lJڒF�4�Tzh���Bk1�"[�R��tE�uO��V+�����oS�M6,}�[}d}��x��
��!PH=�k%�����(��`�)�X��>6�	!��MHP��D	3� �z�,G� ݮ����,c�f-�|q�5�u*���m�cB��5���+/H� �������Ѽ��x-$R�9�T���9�Br�� 8��ԗ	`A���
)3�
���2z��@�R���RlT-�R0� S��`?r��y�]>�k���ݵߴ=q�e6�Z���<�~��{j��mˡV���Ȧ�+���6*����D���̥� %�L�3�c�j�V��?GS�f`�	 {!*��C@k¤�A��^I2&��0)jߘ�%le�w2�K�C<�<볳ؿ���[;�K<[����V���.��*!��m+��Y0�*aD
D[WHE)���h��!"�3?~�9M�\I�a`!������./���/DH�1����iF�%3�焠-n^�U(��Da��O7_Ջ���׶6'������ڴ��pL��idJ��.o��oK�]�����M��`�Ř��>��9zB� ��o�7_��v����[��/�>����Q誊��/!�Ã��͟+����<�J2�\l�o+�`�D¢Z�E� 5~��$�d�F�-�k�}+v]�D7VX2�W^�J�T����i{�	�槣�!U2�bk��Z'��`�[v��kw�~�%2� n�>�{�8ҌIf$(PM�#�f0pD�4� &�����܎$t��Q^)iՓ�5������Z�t�i�a=�R�P.��	�2$)����<!���JѶ��1FcD@�hID)�T��"P��{�Rޥ*-�K�=�z������(�^�VN��BJ�F�<�u��'5�AD�O���[�q[y{FEP������PB������ws�fԁ��B$���0K56YH� P��8��1�8�ᵕAB�~i��s^���^'���w��DO�ZU��_�.��B^����!��?tf�����0*~=DJ%�>���Ŝ��[�yBN	77Oq�&�֫���k��/�q��BDPR��`���'����'8�(s��4M� ��j�����@M�yW������BS��o���3�(���Bn����\������nșaѪs �_Z��%�ތ\�1�������O��;�����]|v�o5�&|(����������9������<�ђ[R�1b��%�Y\1KY-~�g�7ũ?���@��y��Q�%�ף�(zvh���3!��n�;�@�����7b�線�F���J�Lv�"@z�0{�v@Ĕe��$�P�g5�V"w(3&9b�	%�`W�}��j�����#@JFN�QJ�`��P��r �լ����h�"�(�F�׷�>k��F��Z%�2 �)f��~5\��@�i&���y�R�#�1 F�u����"�!�keA�sQ�T�Ů?FFL� �ϧ�q'˵�H盡��]��8`�ce���4�e��1&K�9��
϶΀e��ʘ��a�:im�|ʼP�T��R7��{U�x ��h� T�ʆ�5T�/D@f�<IP	�o�������c)��%~�i�n�/K��C��nG�V`(j������k�gM�=�S���I�Z:o�v�TK�<"BQ��������equ��d�>}�y*H�#R�8�v�ǓgO��l0������)%��<�\
�	����Gf��%l���7u�,,�%�ô$�َ'9K�@�r����:�җ�3Q��6�h5Z�:;-����)z�LY�u�2]�r=� ��2�������Q��|y���ǃ�+>,����"����]|�o��S����<}ea6��՚��I
�-~���Xr1�doz~d�z���������j-a�3�W��X��L�L��1*#��e���5_]p��aM�5�A{G&�L`����Q2a�#2f�Z
 B�� ;$��5�02�x��F��x����0F�U����W��r�%	���,KZ�v���߮�sk�c	�F�.��j��S�-	�Z7S��pn}�T�JAI�s.AB�H� �(IPf+�4`�ڎA�%F����m��J�5o�HWR��{�'�����e�`�t��S^�g���JʟP��fL'��d��`��ք�Z��e��["�P5LXZ�F��s�X�n{E������9ke+��u�v�1��Q^+�sZ:A��.9�gJ�mW��E�����]��wj���/	5����p���J�Q����R�tx�iNl//��G^�~������ FJO�1��r��a�ʌ�xDJ	Zex�)�sO}���a]���㥯�k�;"��Ȩ��\^c��V��$����z�S�W����I�z�^#3$��6B���?���/������}��O��cߌ>p��������7�v�돤��?U���J:�%�D!ɐ�{2��R��s��r�~��K&o#�j�2 �z-6Ӕ���9x�ڼ�x�h���z�,����|�r-be(b����q,��2n�P��0}��S��j�6���%aFƬ3�L�2c���l�!�pG�C�ц�l ��xF�R���,�z!��OX])t�$����x�,�{_�V��1w�J�
��� �1a@ҌP
B�Z��X )c.Y3rJ��>�gD�F���E)+R*`hQ�ڞ�4�*������S_���5��[h�y��������0+����e"��Q�EiA��iz�7&2Mlg�$��0��T#+t���Ĭ-�ь 5�Ό.!K�5�l�n.�����ڪ�_)�x�ٛAsj ��v��
���F��I�7���W�S_��("]�o���9\Փ�����QE�d�C q@*�<g�R.8'l6#�FpQ�qy}��|�u���x�����}�� �i�8L38D[����	i^�,����3��s���Qp�F��$c���oxnI���J�\�{j5�:+��8n=1L�����\�e ��L	N��
I>�����0=}��}o���x�o��T���%���ax���(��G�|T&�Z��6�	4Z��K?�Lړ��k��S�Qd�� K���Xka���Xv�2?��Kq��/8��V�t��=ʿ%C�6��"F���������ѫޓ�:oAT�X�M��Fւ$3�L]�[�j��z�bε�e�vW���8>@���:C9#�Yp�����S6���εRWt��}�L��n��lb1�w `�)،f�
��֖��c{(KY�KR��X�%�eA��`�C�hQxUkKlԟ�n�?m��
��;Վr���G-�g�hԽ�h�*���! %,^��>FcQ�GҌ[��5-�7�޲��%���q�8�&�ڡ�@�Pڹm
�Ң���[(Gc+Dj��T���E�:/����K�����װ��Y{R�H���3��(��#pzx{�W���2o�C7ԛ���3*�[�@ss@�qq�4g\]]���#���8N3�d#T_{�%�~�d)x��cd���T0�qs{���{�a
��rFN�ĠYd��lRks��t���8Y�;����K���:�������H#���ۺ�I�Z���~���B[�f	�"��A(vn�:m?rI b��t�^��/��>���;�>��ۿ|`
]U������_���{~����h>��2A$�g#����	�j<]!@� �Z��&&�-�D;�5i:��d�V�D�P������e��k���y�H�b:������;�[Љ
;�Ӈ:�KA1��0b[�Q��)����ژT�@�2*�n�aP����lY�(�R$HP䈩�"˄P�B	�C�Ad��$A�%=����!�xe�j�!<d�Bt���&a�1)���u��{+���E��qq���ŦTJ�BEj��"�pE�����焒	4bX:X��Ա�@$BΊTj�
� I	b`��`?�΄cV0�d=�j��P�h�0�e:��I��v% +ͣ�̖��R
��.���?ۗllPh	�U�	`LK)(Z :!ȡ6	1!�4����$"����JMk_]�F&k-j]�
��l����������4�����	����E�֑ �)YIT��ֹ'���ւ����v�m[v�,�Ѣc"]�-L�:�gevF~�>5�n�Y��+;��i�����w�l/����ݣ+l6�4�����f��^������	�b��<���,'�x8����r�m�{5M���#'
�}y���vΔ�q����L���g'���t9 �o�u]����C뫯'��Z~�U�؜�j�$��I~�������������߂����|�o�-�������=���I���t� 5���,Ѥ��-q2B�Y�u�A��ن�W]j��.�`��O(������W5��w�Z���|�$윾�Y��\� ���7}A���[�U-.W։)�M�b���,����f9X'�b���-CY��?:���@��:C���L��E��������� $�Z�o����,ٺ
�nNUa��ߝ%�����D�c�E���m$"d�q��fQ2�T�p HY�&�D"D��`���5z*�\�X7-����o=S<>�K대dzZ�*ζ:XNH�ԖF��=��c��Z9���a��\�Jw�)Ag��^"E! J1_�,fK����rWB����Lw��(�Evk76Hm?��[	(��a����e�`�|v�������a�Ӄ�&�E�5�Q��f��J. �}�j� h�H�S�f8�Q��q����z�-sga�Z�jkKZR��i\ (6�t6`ETPJF�'����#����a�-B���RJ��v��	2�9c�#a�ݠd`;��n�SB��)8��)M�P%�J�!�,,sKe��{�x>I�<Y�;G�����z���c��3���Fw�c/_���>
����:�	l���a.�24-�D"�%A�d��_���y�}+�>�<.}>0�>=~��똏��W��GJ:��Ɇ���#���T�]J��Z��5�^��K�.ٱ���ߟv�[���`
y�1�f�)�=v}rg_��(],����p
�u� m�.�bD`
��jrגd�(�H�ſ�P���EfZj�U�u���Z�EY��U�	a�#�	*���H�,�ea������DKM�Z���0Е!Ж��0�H(�\=j�GV@R��j�s�&��J�zܘ�$"g˼�LP@����Aр���@V�����L���18��ߺ�qCN�����CS>��;���@Kz����q��ǵ�U ���mF�V�3C�2їw_�Gv^�a}�hM;��Ty���"���d"Y�Bɦ���-=y���=�P��� ��"+O�5�i}�W�\=c�)�O�w�V���*I֝�t�m?\��f1�g��i��[_��&@5A���^�j� ˄i>b�#�`�MeZ.���߁����A�f3"��'X�RPJ�dWǨRs�Ob�f��f��}u�V�ק�)�ޟ��q�峽�����Ým��xr�r"_t]]�Ƽ
 *���=.�2�1���O�g���?|�����	�������UzH4g�o�B��$�w�:9M{)Z������dP9��E���U��Xj?������[��7�*rfMU���ݤ����sZ�Z2%���0%�Ɇ���&�B7Nl���i$��5��דs��SR˜O��:#�D��#����<�;ͳ5��d�&�N�������`j�nBAd�z��^/�s�B*�lXw[k�o����[���L�o�m��a� �%�Υ�Bd����T���U��CR׮������x��w��?���Q�]� �����s��vJe�X������֙��������J�+b�!��i��[+�:e��#v-���K^Rm���/�ql�^�:U�
ъ�4/{CZ��v����7BNAulks�AK|v	�-�	�>9�X��*��_���-�R\
3n��|#����)��A�@ ������vLs�������^sr��@���%��n�#�<M�ӌ� ��<�w��u��{KM}ϟ�����-���'��:z�*���V�ja=TÔ5�Xȥ�L�Kӌ m��@Hy�.�����|��o���>�m��'�s5�Z��+���m��_o�������_]�[HI`d�f����j����ZG�5;�ex/����<I����4�y1)�S\��� X�t3=�=i^�T�S+���,�co* fD�  �)b��V��h�,nZM�B��Ų�u� ��h%p�Ե� �p�������.j��[^i��*Beu�u`E�ʢ�O̵%[M�6/}I$�,N�K���B�;��R{����-�c[d��[+������S"�4|���#�\[̮"��;�t��[������?������$��0��.m?�?R2�5F�0��ތ%$cЪ"E����wژ����v��[��Z��z��+��y5"[0j=^�ʹ��\vHK<����-4�ʭA�'�����{=�=w�2p���i���-	�˂f�BK��?`�����
�,(*8LGp B`\^^ ���W^�v�E%<~�m�\����`��y��B����0�RrgS�ڷ�Y�b��������c0���g�wΤ.N���Z�ʥ��yYRs:Bw3��X�s�:��BbslFg")��ռ��o��o���o������k?��k��U��x>���%M�?O7����3�N��*(���-RȐ�@��̵��	�^�J/�ܵ�[��?>�b����+�6}�y��^�:n�ĈȨ��C��3O3í�zS�l� ˀ��	܇*�c��=%Q�
q%q�����-��X&�e�D�D��Źև�d4X��Xe|��D ���1ĥ�nsS�G��.����C-�8�d,��;�a�z)W{L�Q�	c�"r1ee��Z��h�t�0* �Y�S2�z���kAk�[�"YF<�g��E"��J���&,���������/��+�۶��B'�*��w  c7
�MR�#@�+t4���|)�Z�6��3.�	]_Ok'[g�3B���@\�z[�$�W+O\rmM���8Y�t��Pܺ2R�`�$���s󱭳�X��'�:�V�^-�g�>���������c%�|�*/8\�v�~� ���<ς)%�ĸ���؁'�����g��O{1c�6O�@a{�E�)'�4W�_��C�Z5rNo����؋��9�876ϙ���`w����l�K 3�E�V����$����R��UWC� (׮}���Q�ux�J�v�q��l/���n_�D'���B�����7��ø���i>��r�}%�#4Y	���敷6��(T4O�� n
�y|� �y��Y�Ve�R�W`�Cz�����5�� ,�Ks����l�1�����W2���X�dS�T[��hͺm��)�*���R�[Y��,�)��/��QɹR��h��z��&|c뭬�<J[(,Bz�G6���F;wA�9�VZ��m;��aE�v؍�0�=�f^�Q�1Ty��̵N�j[��yW  �lSڄ�����Ҟ�W�z%(��g�M4N=��/ܞ�#�t��m��z3��Q��5��S�}��Gh��"���޻��u���mQ`�z�5'$�RCkW�/� i�EW��]�=��]W���q�qzv��\�h1&{:�?�x��P#��7��|�|��[v�H�3�[~Ƹ����
yP�h�x�q������~}�5��?���/ �#^}p���#��<��^��ZA�5\rz�~�Ej���ߝ������P����R.w���@��3�)úGl7q����rv��kc�'
f�5�3�}T� %!���a�o�0�Dz�~��e�5S臧ORP��g���%~MI�������l�W�7��׺W�H��@��Z��N�u�,�RA����thZl�5����l���n�s����A�6V�Z�VJ{%,�W)� L�1�ujS���K�w�w��ʭ�����ɖo�;��PK��("�4�Ig3@�Y8KD�h-t#��m=�ﴇ�1���N)���)���Ӻb4*�F��V��J��Xp9L8@��c�
e�D��@�mp,�[IlP2PR3�IUPuN5��L3�d�T��($`�`+�w�����0B5Ygi����fw��oE�'��(�n�Q��P��3�����H#Ѯ��	j#F{�{�F;��]��(� /���L��Uᮜ��̴�s7Lq�����3��{�~qB�.�C��������j��ɯs/�u��G�!+����f�� ���BHHl@#A�`�[�������px���$�ݸA�{��b�C�#J�� l��jr�����ս�By����֖na@�y�����V��v�Ӭ��X[1�?YJӈ��p�����}��Xߤ��æ��bU�(/}Z�	P������c�~7��I��;�<��0��(<��>���|��5Q���u°�����u)�H�H������*����Zfh>2[-�m�:�eQ*�x�zB��E�%l�\����B�8�N�z�Խ�J*�+�2j��Qq�Sl[��*��6��D�m0{O��^��%~�5	.��` #x�R���Q�����:g�!����@T�"KX�?��Go�-�K��R�Ӟ-k�z��ۮ�e>].��ϻNAl��Vf�c7������B�,(��deL9)��W<+��	`%���[��U�)[׳8 � �8��J�t�h����Fo�z摟����t�N֮�&
W	E�=����Pq[Z��,K�0X�����ӸI� k����:�KkV��C����b{4��L{H:�,���،anSW^]���Ӕ岎��:�O��w�W�N��W�ѕ�������w� �_�aդ��$3���1[\<��������C�Y�%!�'�4c�8N�l���W��%A4��f�1s�5gِ�ߵQW}~}�Y�����%�@ݘ��,]1w&�Wj7��g��T�ڛX�j�3����Y��^e;�A*����*� +7���v�B�)�؆�گ���|��)��@��^y�o�q��%��5��o��<6��o�<���飒k�m��j׷�k���R'��X�;��V��إkTU�k�z��O�6�Z#�v�Z���i��}��鲉��>��%�K�����]���,�@K2�G�&\5���}f2�N�Ϙ�-s�T�ր���5���T D�jMD�D!��p�~w
�a�?|qo��{�j��Y��H�Q?���Fp10v0�i2Y��P̛��i
���y��6 �8@UpLq����p�/8f9)�i���%�4å��N�d���{��('��>�xH��H�ɇ(D`܁�(���6aX>�=}�gs�tc5	�v��s�d �$�#���k%p7��ޡ������<�O��\��rg/6#K�u-�2Al��-$�%�k��� :b��@�C��ѣGH�Ʃn�4l��KW`:������n/A���� F#�	�!C�#(
R��l�6|�:7AOBF����������٭r�� �JݘlFX1,�\�����������e�q`�`��T��7VT���h����*P��º��dk�L o?��~����Z���/��e�_<��
������݃������2���{h�!�6��%n��NK��gh��в��j	�Mi��ePb��\��i�ƾ^�u�d���4[B�	��%|��՜�����z]����k�n�[fk��V�<@1#�����(�ڶj��f

F��P{OB*1E��K��`���TP`�Ig���JR��
}�ث�Lt�+N�c��8�/����}5�̓�{	�:����� l��e�P�eEfE��."@jMgH��z%���ƪ.���v�EF�r�1)��8j�mfP�j�m�.}��#��X�-�Uo��;���:�?�A�ڞj� l�@�:?��,�5Ԩ�F)������ޒ�t.X��G��ZjY��[��^��<מּ��x��~�2�p��Wn�]3��\x�;�|�pژeG<x� ���%n���"l������C�f����K��n�!�	"2vW��!�"H���'dN���?S�11���0��+-gq���e�/���sMm]U̵��-9	�6/�tG�ܕw�k�P�=��Q�8��hg;�:TZ"rc�V%���ԉ����\�N�8|'��C��m�����l�^�없��B�g�0I�0>�L���H�o���x�2ی�>AMڈ�6��&ĕ�g=)���5����qIu%�Esr��k�[8�5��m�C�(��,�f=��]b�+�e��fP�JԖ����J���&�{9ࠊLmrي�V�uB����{�p���
��5�A�x��*�gɘ5�:�f8����X�_U��_.�"er�'���5w
�<gZ�S_k���F&l�a�@
�-KKQ�e�}�51�~����$dp����VZmÀY��8�Šh~Z��}�g����*��S��5�{���ݤ��"��q�\B�K����[-�b�-����PY���áf���
S�\2�B�%������?�~nD�oX�W*u���~��>C����j>G�{�'L�z��\X��J������D�,(qD^~����n��G�o�b�靈2=����T���C#�w[d��Y�g���m��3k�b�D�]������O����,���o!�u.��"�sQ�зOO�[Bx����)�X���S\�?�(�t���"��4B�� ��5F�Ǘ���7��}�ZP�_5�>��BJ���K8<��o,i����$iߕ���iu�r���k/�}k����uV�=	�	��X��!%SoJ6p�=X۸U(�,�T�=x�K���o_�����}Z��OX+ۯڶ�)��H�FU�����7$��r���y�@���Ba ���Y�� k��V!K�5#iFAO��I�{�}z�=كϫ�~�8����s]�ks�{��%[3cc L�T�Ú�D���ux�kB�5����\p��E�ՆZЀ��'2���:L��Lh���{���#i,Meb�yu��)����yU�H�-�hIo��b��kyd7.�g ��n%�������8�`�a883D��?/��ד�֊�q��z�מ\_Wk���dS��l�nF��>�C��@`_\�2n1l6@P� ��S��)��裯���o�`�nno1nF���ţ�݀I "�AD"�.���ah�0->��$�{�_�7� ��쒯�N�a��5��h7TE\�n�hj]	V��8yԶ��O��%(������%�K�@��&�|/1m~p����p��?��oc�|���ܗ���B ��c�� ��b��$y��(�CoʼNX+���1��&��zPa�g}��[�����"��,曶f&]!0�r&S�= S�ש`X��d������s]����ZJ�h���*��Uk+1����
BU��YۖZ��x֚1\=�6���X�u�9���O��{�a���4�}_hd�F�5,z�d����)��\yX�@dB�̢�@�Z�E,�Z`��52�PJ�V�!�E0e ��1�Y��S�SO�z� ��;��4�b��e�W��,���홝@�?�ٸϓz/���{T ��/B����?�`=�{�����sK�wu�"	$O 1Y�hZ�]E{�}���Yb��Q0gk�x��_��c�gk���nh�`�M�ٰfCjb�x����5�,	�c�2� 
�0"�$�#nC5�6dG2 	��&"F�$[��Z����dDkBk{�������p����z�¼(L'��u�Z���O�A���`H}_����'_�F3��'Y����%((BMn��Xcm➅�*�,5\l�ܯ1��Ç��t����돽�0ח���BWU��\\}�r�n��L��'���a+���^k2�f�t'J�@$V:C���VZ���,�'��j։F � ���0�u%���RK�L�4�ܼ�:I�Jg�0[BA���xemC�pk����}!V�$d9�G0cF�Q3�9"R 	!"`����j��q�mR�5�4'c=����6�cD�@(A�����&ݽ0s�Ծ�OA�o`Z��+V5�R4����Z����i糖}]�{u�g�"JA$j�����Y�P�9 Z]�%"�ጉ9�D;a�`�)����% ��CY��`T�� A��#H��~�U�6�	�V�mF��%��y ���3�z���r��� #�*tp�B��z� �<�(�V�&��P&�Z��ԉc rM�C#* �� ]���s�#{ُm���yl���r֦���L��lu���̩:�C���+�w�-���ۀ"�kC)1bă��\\���"4���1�@1�Z����e����K��x�Ÿ�8Z`�a�NV����8��3�pY2қ��
;��3��c=F��e���;�����`�:dy��B��UUPX��"�Vm/"�*�ɺ8�8�"A+%���t!՜$�Z�.3�$3q��C������O���ӗ~�����*
���~W�����=�]%�L:<�(y��r�^ �6 D{��� Wk�Q�2WS���|AM�iZ���[�7�
��8��h�!��$'��ڗR��A�4�
z�u8���\���r�%�ED�D���w��/h�}{r���D ͘e��r�Q2
8�0�e����5bĀ�G�&h<b�J@Q!��Y����g^��	E%��xe��ŗ	R�ss��	oX��~��PX�˒���c�e\k˺�V�96�U�����z(�,� jT��J�c%��b@!b ⚓`�������u�<Z��XM�"��"��rPeD(�3D�?=�w_H�%*�)�a��Kg�Seֽ��Y���������z�L�X��ژH	��^�P�Ӥ I�f@�w&K�$������Z�bN��źr5���^���0�:H�e��/��JB�7w�m��%����q�PhZj�@5 lPK�^c��lm	ow�QA����T��@�݈a�S����4^��� �(GP�QR@�;�������؎#<��	�no���*y���"jȤU�gW׫�yzX��	�ȩˡ&W��'x[����T��4�~I��Ő��˸Vjlom���.h�5"V��fК|�0Y*
�ĕ2���s5H �BTg�#�y�
�����r�����_�;���W\�����{x��s�����XJGk	ZR��[�[�c�;G��z�z��S�;H14���_8�R ��;�0��и��j�se�`od��^3����B�fL�ק���>�s�qO~L���(�tƭp[�أ`��ܺYu@��D	�D4��:�qd2CI�oy��b��TD�K��^V	'[��B��E+[)��z�p���K_���Z.D����] �!�ZՆ�T&�ƃZwd�gE2@���])g 38k�ôE��|���bh�s6���j]�kr't�}�֛�t�\���3�Z�J�`�� ,OČ�Z�ީ*To�NU�������Z޵<1õ4�.�y����~��>��A{ц��W�%�� ^ga!��Ujg��h���w`����Tp�zߵ�'x܀���K�p	�> o^�#�� (yh���ƈ;��+\\^�ٓ'�}�� ��K����MYS6��K'>c�*=}O2kk-ߜx�]v/����J�tMO�֏^k9�Z澨"��Кoo�**�(R�b���~�"�4!�J"�+��_�������S�W���WT��G�X�����9O�ߓ��<�!+���;ݞk��ORU�u��������2��շ�w�P� o.�����6h�(J��4C�h�1�t�f}��)���iC��{a�k�
^_�П�Da����(Gܔ=����q`%�8D� REfhIȚ��l�ݣM��楪��4%�C;�;UL9Cj�j�*],]�5���-1���Ig����)�JǞ��1^��� _'0�L��4�U�}e-H%#e���U)G˒堰��R�X��@#�1I�X��Z��R�ʓu���eo�m_����^+��{>�*�v���'B�y��������u�_3��R�Pb�W>�>	�<�F����a�6��ySpP� +��0ԻE�9�痽z����w��R���=I���ܫ��*����,�oz�Gݓ��e�}ev5.�1��L�#����+���a�h���T	2�@܀��|IO1�Y0O���x)���4(h,z�S�����yt槷���|�3���n��$Z���uiy5�_���NX��<|[1���;_�c��٠�Y�͗0���7��O���>���q�_1����SF�8���������f�t i2��+�d��9�ǘ$ϐ2e�t�tK��BO�@�h�vYy�-M
��+��)��#��5#�($g��OG��4�=lИ.4N�bP�^�꽓Y�}zS������ϧzn%�I�*�t­�q�G H<`�������b;4��	�6 rDd�Ԋ�l�e�pT�̄X�F$��5 �U��V�є����Z��J��=����B����C������.���w���B.�Bj�C��:u�fl���DB� .@V "
d��ÚpX����ө�J�4s�=�(���N���k�^����-9HWR���s�k[Ә��\�V(��a؀���J�Mj�j���Lm�*z,ݘ35j3XܝZ<^�|tB)�� ���л��y��e]Ob_��M��g�<ɰ31g�l�K��^}�RW�R;.y �2��'T
�9ˠ��_�x�1��'`�,Pw����Y&��$=��^B9c�#�e�=�JB:�.�V�Z�~v�C��qT��z_6gf����	�� z��I��>��UC�-����K�Ӛ'�T�75���H�U;(J���}�*4e>��0����DM����-�_����W�C߿��=x���������%�oAe����$��s��o�&�U�O�&��*o֚�~7��lr٩��#�C�\!lV�����!
P)�$h��!�(M}-�q�����z=,�)��qy�����zs����Տ��3-(:c�#�2#�BÀ�6���l�Y��1R �`3�À!Z����AҌY�L(�P 
F�ȴ�J�QB˕^c��~n} �IF�fdQ�tv�������U�]Z�)���Ϭ����j�DȢcғ[k�{3��%bY|��]�	<%F��5k�����QVh�R�GPb;�3�=�q�J?�<���kUg	�M�4�5�EkExn?�ӪҀB	d�(�:�������KfhJ�N�#k�ޛB��5]f�E!�*�v�5E�l_��l�������-�sf��8��טr�js����]�������,4�;P+�ۂ�0����q}C�a7� UwU����C[ JI��.��2c���&Y&��ץ5��2��ē>�,T�hw?�51�^�W��./a�u�%��yF�������-��@��Z(Hebdɛ��[������ H�Q�ï`
�V�^�?�O�=��)�_�B����8N{\���w���������&+��Q�g˾�t�J�ݞ34�2]��iյ�Y�ź��5����r31B��a�!l.��%4n!a Q��>���9� T9+d>��	����#\����k3�վ��ž]Ss��5�B�����[րH��k0('CDd�h#�`cgE��9?E){�F����2�L���Y�g��%wn�<�~�p����ڳo������[T����]^�b���]�;Yͧn�{�� � �ܛk����GjR����5-��W�ք�TC>R�q��ޠR�M��I�{��ŕ[� ��b���:ɮӎ�ۭQ���]�֞�B������?��Ѫ�[��t�0��V+�D����JR�&{N�l��➽��*O�>�}}/jvr���E�S����k٥%��=.�8�J�a��3�1���6�1 V�j��"(lL�ǫ���3��"Z7B�2mP;�Ae���sv��D�%gD&%����F������,t9����(xj�?�:t��e��慷�������M�6My��n{��1�Y����s��4MD��)���n�W���_�2�_�BWUdI@�1���y:��<��|�A��%X��kY��i�h��"ٲ�A�M�W)>���8n+{Yh��z��F4��<���ф	�fٚ`�Ƹ;h������o�iM����~����Yg`V�������"�!�k؁,V��\l/�9���`���l��aB� � �
�"b�V�"������_�Ji�j�D��/�a���]K�[ؖ�O:/�Y�%؅:*%��߮��b���9UO* !�1�����b�T���꺔�\2rQ�"(mR��b� ��L�G�����Ę���ݧ��#��#�sݱ2 @�HW��"�7Cc���<�P_*j�[hآ�����j]>���d�G{MO�%@�헚cCdm��(4[��h���P����FX]�6ñ�Uܹ��ʭ�n�2wd���㉫�iL��]�ڶ�&��!�(�J���lz7��IA��C �<nA�N�Bk������9��:T2(^��^EH�1�e�˴ǜ�eo3!<`��,��S�ķ��K�9u%V��ͳ���sWKN����������約7��-��>�X����{c�qҦ��\��������;_5�znB��f����V�,����VAdά�iSb��4�G����o�q���)�W I��V��e�ovWy������曧Q�[��7ŝk�j����(e�JsՄD+eVyh�����e�}�Mp�	���r��X�h#)����-��@ PV�6\�BW"ê�4�C^�U��v��-T�]���x�)9ka��D3ـ�Y
�*�H�L) "��1�כ+��Z�Y�(�ՃHFQgt� �8��8\#�g9���r�� �.h,V��8�u���������i��M��s�r�u��)�u��B�s���ֽ9=m��H՛�'f��1D(e#��"�6�Yj�W��fBa+��`i�f$)Hj�4	V�:q�3!�ơw�Y0���,�}X��߹�3%�ZW����YR���^�Zk_�uS}J�]�/��ј��Lа��B�(ı
��.(����~�����`D�Y�+26�(�Y�Hd�"A	��4�D�n�P�0��)�n0��n�>��A"X���X�qbʀk���3w�n�E�6",|��MX�e�i�����j1j)ku��Y�#t��$_�>���J�0@e5݂�����e�x�3G��̆IB�	Dl��f�۾0z`�נG�`Kl�:WC!U�W�pe7�$T�~&]��Y([މ�0�DK����ʊ��� �XS�
@3��ٝ����@ �t�[q��O�`X���B��d����������)�L)a��t��������r� �Ǐ�}��|�
}~�E�+��G������?7n���g��%[bKk�
IPI�bY�Z2T��shy��q�U��r��P�%��	}��Y���� �n�2o�e�j��P��נkņ���Uٮ�
��̛'Z�O(�R��;��VoN#v���K�-��H�1�#]C�D��4�0!)��_���+�m_B
�y�})O�*�*��vTkg�zl������2��̚Ʊ�&���)��J̖g�;_�xO�[���iĉ{���m"]^�ȇ���rm�	�m�������)@(� ��qS!LaNQFD0���ϋ�G﹧��:���Ӽ�j������`�7���E!ZZU�R'd������F]��~�c���X7�hQ��/˯�gY�+z���;m��RkힻS���J�8�ľ�Y�<�U�~lʼ��6j9��Q��֫�]�(Ue(G�q x@� �@���!8�`b���Ⱥ@��ҥ僄Z�Z�PH�t�q���3Ó�ȼU����=+�?���KP���u=4���Ժ$�M̀�Ϲ(��%���Ͱ.�i�槳]R���s�:�ψ
Y��]�"�&�3*6���QUf,g��p������Ӛn~��/�J��
}�]��K���_�y�w���7��3Hڃ�T��%���uQS/K+y�d��*%���%��[u��q����H�$7��uh{��(Ѿ3M�1� �q���Jn���@WnX�]��Z���(,_?�C[2C�J�Tj�oD���n_��h�<*
���K&<����.no'���\?|�_}#.����� '��|��6�*���v���=��(��4;���"��k��=�y_g����w~�_Ӄ�R��֫-{?hM>
dT;,���0ԟ�q����T�dƜ2b�՟�Q�(mV dUL	��!�J��w/�ݽ,E݇�����z�!uo�����ĝf֚�@�lUzS�zl�җ��t�^K3i[\�ACj65$ؠU�J�����ݙ�:�]IS�R��T��\���� �'o��f�/k~���)@��~�ү�gu2{��ٶ\�
��A�`D�&0���İ}�x�b[{T��=�pUv� ����GFjܾ��}]��F-�Z+\��x9�kw�m�5]��J�z;d{�b8Y�~�Mw*�a����re�Ȫ$�WA��q����J���n�递 &0��������2t������N�� ^��U3@�f���F�=@��䧆���Fn�z��O���|����R���q�3v����p��N�gߕ�O��(�M��*	A������ټ�R�I���.�G/�g4V�T�@�p(�d.�����Z�0�!��oISJ�8�������3쯵�
zO��[6����rP�
2	�����#<ܼ��p�Q�\;d�FTk3aƭF 3T"Bq��^��F���8�|���̄��;�ᖷP�w����F0��֔�gZi��͗��ti�Y���^ѕ����E6N����D�Y��"�����ǫ�^��+��	�h�~�t��l��by����y�\����\`C5�ص[��%����	�j|ϻV�^[&/���U:aIN�����2j�T�r9@C=w
H�B[�)�ɮ �	a�h���@��|���ߡ�K�]IQ�aս�~�������wQ�m��{�-���yv��:�FS���/����:QD�׀�Ge�F�x����h�
;h�����zK�[�ZC)�0hI	AG`�BV�sҜ��,�\�z���sسW�궩
ͼ\BAf�h�R`/Iu}�I�f q �h�kA<Խc��@����e�䄒&n߂Nπ�4�b����W{�$ɲ5j3��,���Ԝ��᎚@K���%���Ų�e��
�2�Oo��_÷��4߼���_������� ����r���|�����c.�H2��V�-3��+b�:�w��@b��J�B����_� Ӿ��M�8ڃo��Ą1T���E,YAD�5�ɳ�ʣu���E��J��hu�����hy�f��UA�bY� L�_p5<�[����%!��X���v�c|�Ww����#\�+��I¨#F��[ڢ �uU�4���Վ%���{͞Nծb����ђ8W��~Ч8�{O`���g/	;m� �j���r�C@���`�b��U1P��f�_a�Y�<�T � ��c�8��V�����������|ߟ�ö�jm,.�=��ژ����<����51l9�`�6�7 �y#��U�������ː�u.�c--,�(o �ސ�V�s�2u�x��ܗ5X��֧1�u�.mq�uX��?S����o�K����q�����Vi�26P���%(l���=�$l��^�kv�ld�ʭM�D�\�`�ɘ��Ҫ�5����Z�l��ץ�b��Y����R��A��� Es]s{��֗�r`�#�"�:G����aD/�h��1g����h�Q(���q@>��!T���ٺ���:���ۜ�����v��ԫ�o!HR��9�����h�%���̓7�EP?�(�����蛦�����x�}6�t ��h�2�4�Ħ�I��<uz]d��X -����i�G�g���V�ڽ/��@Sb��K�U��%�X�\����6-�5���Ք�)NsG���P;�u��N��^p,��#(J�]�jз��x�6@���C��t�`�M�Q�q��f�!��������!���f��y�m� Q�Y�8n�[�[�6(�,m]e�����bG��:�tM��d �~��R{�B�?gs�ΠR��ɠ�E��Da�Ը_�m�U@����ݰ��fkS��(C�"� ��%P����F��_|��9��l�Q�N;�R���r�˄���ӳ|Oּ�Gܼ���^Ŧ�	��b��[� 6��8L�o�PZ-��&ݨ�S&���04^@ɼR�r3�J)h��E�V�v��N��Z�Į��t�f����l��R3�z�0��%?�Nd�赗,	�=L�.���aİ����#4�P
�!�#��5��Fѿ��u韮r��[P�@����� g�L�4��^r5hN��b�-�ag,t��Ka�g�*���#Bl7�@W��}1#�!� !4A�#�a�8n7W���:����� �`	�*�<bsU�RP@&�t��@Q��Ȼ����/���;ZbvԚ#im*ղ����9 
K�.f(���_�a���?���Gt�D��!~�x_
}��	Ⰳ����r��J�?������2=��E5j}�>EU���)�˽%�L�[)��˼���baXL�y�Mq.Y�V+�F1J�#Y	g(U��S�U�Cj̿��!e���ZXh=���R�²��O�V��)�ZA�����Z�
-�&�0���1Dly�_`�[l8b3�@6A��#X(%Ϙ��WyM2C��pa`/�ܦg�ϏqC��q�0\a`�:<Q� �ڍ* {BU�m�(P��yH��@�x)O��noc�f՛����/��Oz&�:F�|�r2u�,Gf��:8F
�d޷���B!P�ҡ�	�)��4� b����YB�Bkˤ�D�ʬeX��
�T&�d��=��߶>ն��WyZ�׽G���'Dj����� 3ۭ�0��]j�3�P)6@f�!\>��	�fH�}N��@���Qfh$�m���k�w'�)�0�(K�s����,��:�ê�
y5�r=��i�Z�/#E��K��&�j��=I �U��.  � IDAT`,�� l�4����/!k�����Xe׋CN�qX��j����,G�t��'h`Pe/�2��i�M,`)uݖ��+c��������^�ꥶ��v�\x9@����7����h?0���/@�7V��e��h��[�TD���9Ȅ0[h�ە�Z�v�?�q�on�<�,)��ͩN�@���Z���T��#���4��B���*�..�'e��R���/�S��|�"���'�V�?�e���� y�"	H��֞C���tD�G���$V�2�)9Z	�����ĨEi��]-�q�J��"�ʹ%d�B�tDψS��ob%��>���j�Y�f^oՅ�0gT�ԕ�m�R���=�6`D넮��{�'#CsDF� ���]���-�a��.0� bE��(e`vd�DŁn0KKƠ���%�7�P��K��n�4���F1�0"���W1n_�̚.jG+dj�H�VE_U�H�P��-�V��BJ�}�P���dZ��b����P�X�ݩ6����C�f �Q1cGT0�3�K���)�H��Tg~�	(e��q�3�9C4"�F�b����{X��b��rY!ZVa��K��y�E�/J̨��T@)ٌm4��~�51��lS5�T ���v��
� ��I�#�8_����j��@a��Q��Q��ٔ�0�6��G�}�1`��R�ڌ���՝���?�����@o�K溶��'�;�P��,��W�Yz�=�:>��$&؋f�����y@�=; lA�L���
 c��V��{Й�׺N\@�Vהn���5:���hA��4�\�"�%!���o��CK�DN��� ���PB�E�uJ�v�0�Ȕ7x��6�6���ot0�Zg��/�Za@V�Ҟuի!@�����yzѣ�Ij��Ѝ2"��n��2�L�T���\�Zե���J���FD���nC
�P �L�8�/y��u���cl���� ��e�|�. ���4>��k����_ȇ�����2�@��!%��y�טۺ,=zƘs����|��jwUu���v����F�b�8a"% K��A�� +	�eǎYF� �KE
v�H�\b.����۷v�ۮKWWWW����{�5���9���=_Uu���|�m_֚s�qy�ϰH+
�T�����v�Ik��#��#�8�O��9����|��yR�*脶^���?!��P�IoN$3��G�Y���Pܔ��ω�?���^�D�M���u������3���'*`%4]q�O��Nt��`)x��>��z��b�{]�����U}��5���N(���5N?�	w�.��_.攈Dy��oƙ�=ݢ>M�7��K�X����At1�~'��ȕy�g�>��
X��+�T���dI�*�ԂR
��
X���P債	.�a���Ѻ�cC��l�[�L5����d]�Fn�A����@�r��
=#x���y�Y�5�ܨI!0J9A��`x�@]l��W��c:{!-`-@i����<~��~���}�����*�\��r�K�<2�?䱯���'I����F����)�k?�����hj����R����N�M����S���9l+�F��H}��8�L�R�(�W�z�l�`Hc";�~ݔ7��'2�W��+�\�i�����@�D[�u3�dl{����3��1�z-V���p�YUp�%��@�dj�U^;����p~@_ΐ� }�н�]:&�n�Yٞ����$Qs�qꌲtD�l�ҧ���gk���Z^��S�7���o~�~���(o���zk����_���x�3��B�+>����{~�>{�������m}����cP��ڞ]_����h�
i�'Y�WF�(��U��m:��c�8L�o�`S�>~�YD�P���"�?S
�Ջ�ċ>�<8����sl&�Go�8�Ǣ/�]��W�F��v(���0��$0�**���k{�����-�3

�r� ��� R+XTi(� *�V�Vp���k����QO�Q�/��e$����y�e�3>[߀���v�"ɨ�� ��+Я��l���T��aN�l���X�`��T�v�'}:_9Yf}6�T�sQT%q+F�z��өb�\±#��B�k\y��Uj�o���1YM��d �z$�4�;53��7��ʹSߡ���y������@�,�k�xq�
�g�j���	�ɯ����b���f
��=��� �s�	�}?	@��@_����c+G��m�Q���ki3���=��$\~/	�AB(����]z��_�x�y��7e~b�J�Vh�B�3Y�l� �D�_��'�t7:d���gg��+P�\�(�-��R���y7�i8�#]�'9r����bD(*)tKgٮ����ݧ3R=jq:�����s.���R� �6ݭ��9�����b;����#o0Іw�x�@���^���{2��z.}���(��Q�|<��Vl D��E��(��S[�����_[�?����G������b{����_no?zC�\�oQޠ�G_����}����z���������mO_�L~�>�����iޮ&�="����}p�>�h�xi�B��!L�f��3Y%���!w؄��Yu�a�/�x�<��!FL5����C�������^�Ƶ�u
:�P����C٢h�q�
��q�.�l\�S�C%,�ONjF�����l VT�(�g��	��8-�V<���'c*�>�ؐ�uW�����]��q��mX����3����"���ZO7>o��G"���C��ۺ�p��,X¹*^UE��]�5�鼸1�>�a0�T��X�������D0�*�p�B�5�ucT�j���QDy�����1�a`���N�Rw9����G�M,�JJ���:Z[Bm��nV��c�:W@�@���i���>�y������ ���v���A�R��@�6ɻ����&�:N�i�t�T�s{���<����á��u!C�
iF&%,��|��j���޷�(�>��@���$K�V�/Nhå�������<�@#u���P	=���+4��ܩr�~G%	¸,8���(�.�֝K���
��d8�B���+�Ā�[�:�_|Ljj�<9}L�#�iԳ N'�,
�t �k���j��- 䱫���������|������!�з_���;_��7�x��[����vy�ej�_|x�/���?���/�?��U����7~���Y���j����vA߬��*�;�wHo�	X��f��.aT�O���?-��yzꇈ�5�no��:��C!,���\y��|��=<
��B���S�N�\8��D��1w�����oq�����N�)�.T˩����j���
����	[��, �"��(u�¦^��k*��,1��R\�:[r�PyK�U���T�T�6��9��P<mh��ޣ�RQEK!J�Z�-%�v���kx���qQp�h:�g�F.���лL����غ�IW1?bEaB!E�B���^�)�`���(�Ƙ�����ķ�U-�B��x��h~A�Y�$�{ 1��4蝬����
�#�9W�� �T��Q3��D+��"V�|��d�� �+*���;�A �C4$Ip3*�G���|��v"BQ��݃�ŏ����Ӓd��X�ݠ[o�BG+�Re����A����/<�L�"�"@{�^ߠ���-����O�iUE���	Z6_���0E�z=�s'�ȓ�2�"3%�rwh��Yg�^X}It�qW��f����NP�է̙~�I�	��5�P�N6�7"t���� .[�hD���}R�1נ��S�D���P�h���������S�.��?[ϯ�����,^zԧ��sr��W��-Z��]�ٷ�K�<�}{�E^���ڟ�m�+z_����B�jB�F�!�iJ� !�α0{���� �yM%yH�U �=?���f�J��U �H�����T6Po`�J��ny�~LQ@���ï���L�=�*V��	�����ͪɹ��&�����L(�����<��S�����v@q�o/Ox{���U.P^��g�͊�z�sa��/c�*�Q[K�p(��Z�	`:�+�@�9?�����쫥H��6��A�1���G��ɣ+���X
^?0F��3"h�
R��3�R��pm �Tl1�\ԩ_G4@Xj� �;ZS�n���HV���1�?8e�<R����L��t�FGEj��܀��+Sqv7�uq�n/1�>=؜t�|�B�����%�w3�_�hӣ)}=;������8}��|!�(�o�����rҕ�H)��ie��������̍NKz�N=�
��������uȋ-%{:
�A���3X�TـM@�t��i��>$�hϠ�-�]��[��d�-3�Pj�8�O�zE�f�E�����I��2yd�n_<���J9�Q�
݌��r�K��!o��y��p�v*d[	U̹��Es9�2���r�t�����
�N�0(�h@�����;h GsjFwN�X�H��a�=9�*5Eӭ@�?�^�~n�G����7r����|�>����ǅ�PW\���7��K���|zD)�ԧ? @�'H��Z��v���f�U��l�8����~3�Pv0W�~��K�1�/�̣K��M�y��H�)mt�x���SRoW#�F*�F6	���+��񏾧D#Ű_�P&,���wҨ�Y�DVi
Ewv�M�6<h��g������9�#l�.�1�D7@7+(%2��ޮ|�UW�z�U.h�rmD���R@'0�<�e�`DE���M>�P�L����f�5�
��٫��<x�Zn6h���5�@�&HY#lq��P��2�
����6�B���{�s+��������G���	��
ҫ� �^�'���$.w"�tTu؍d�:<>$��+�O�x��&GA�k6�tre�� ��٠`/�R��|Z ��O��y3��VK�vg�}{��Q��-���|h��R-�B>���G��#�6շx��<p(��&+���ɍ�ʒF4Y\L?���m�t�`�Qg$$�v�d�]BP��q*S��B$�в��o㍻��o��Z������V]�b+��+П����'k�9�B
�.�ֆ��f��r����q��M�hJIL�H��(ȓ��BE_�~Q�lЭ���ë�q�aNw��`��
ft�X�����LK�68!2� �X^}�V;	���(���Ay"�!I&��&� %S��(�Q�t���v��m=E��`��p}���T~b9���?/��~��X�y��ׯB�!�l��v��_�"��_Ƨ>�Y�+DXW`{F��]�_[6���@�8,���10o����(���BD���5u�a�H�d0vB�1hͪ�IɊ�8f�GH�j�$�Z	Ee��5i�4s!\��%��$�yq�,�6�,L�����U�ʨ^ ˂^*6U4o���x8-hz��
\����9ٮcE��\�[,�!6UlҰ����EE����S��&`w\�v��-9!r����Q8-ֶB��
�E �cU��j��@B ��H�;�Ժ�dC�M�8�ՙ�xR,��Ʋ��]	�z�e�@W�R�h��;���@A\�PϠEAm�\Vh/Xj�b�z��6ԥ�C7�W�mw�MC~4!�(�DH�8���0�h�8!y1�.(w��j7���xP�ttS�tk� CB�-�0PJ�/�yO�����#X���ryB�P��j�_���1��yd��G�R��ܣ�(f[2sVd�c�]l�FW��2&��\����ȟcgB�{���Hq�s
�21D����m�mC����z��S�p�J��[�R��j���ؖ��2������?X.֍kueU�����l��:W@����'$�d��,7Q�A)��(
u�\T)�5��2G�: �a|񔎢A���Д���Rn�F&�Q'� 1C��RP��&}�ٺ^A�
��J�K�b�������罭��e#`r�4�v�b����j��D=��T/�44R�Z�:$��u]��"��g�]��<���6-˟���oy֟��F����}�����2-ݮX�~��7~	�w��c}�Lܝ�]�p�{qlD_� %�KDgn�)����/�!�8 �)�����G�Kǟ�s�=a#F�nހ:j�4�����{�O�}mx�/�����~�4�{ ��;�'�|D]6���+���Sõ_qٞPE����	B�k��k���䊭=cӆ�b��.���(Y�Ђ�Ū޵����W��A��2��n4��>��0JF=r����rS�JT��`�TL4�,c@��٪@��P� ټ�ETr8�Q��t��(l~�L̌�i��E
����BN�NaWb,Ո~X?@W�ed�(���T�z9��D8ג
[I�����FT:�!�v(W,4C��9�62�:F-�XM�@���P~Ƅ2Ph�f
��9�>���w���ޕ� ��զ���d�(8^
z��`Q�|���o�.��g����@�[]���zG�BA�8��>�Z�k!���]�Y�i�&��w�B�1��9�cLg8���N�XJɌ��v(+:YMJ�s�^a��:�#VT�i�n��E;��aݮ�v�yfݩJ1���3�H�<���5VR�+0X!r�&��g�U:��#3=�f�
��kp��qj�@A 
�O��A���f��,�z��CF�;�����5�1r��Ό���M��7�<�v�_[١=Q�n<}��R~h�$��7o��@9�����{������������Q��c��
���;�	��y�m}�~y�����*�p�$._�9�0����c�`��1��&)�o��;fJ�#���o�;�J�Lč�i4�7Qls���~��{�AO�}��_�!� t]��36y�ϸ�g�L�=�\�X��*&�mõ]\�+D��M$5�q�V1��F��`�����
 �] �B��c��(�{����ChV8I^deժ>瘼5���[4t��i*`W+�"hm��r�N��
:Tx��Y��$��	�d[΋1�5�iw�
���h�lmk�O�����(^=���%ИXd�y Y����=�2��0�AK�����A��D ��o���Fa���EUS��C�+h��=��8�+�Π�ЭB�g��{-ZP��gm[�T�
�~t���)��5t)��������	{
&:J��$�P�Ls�3�>:�{W�Y8��]�r��(�E�C9�����a�^���wb*G�f��*�u5�V�|��i����jzK7k�m+�]���]ѯ�6U���M �{�'r=GzpvZf��ᨧ�:Q��2n)	�ӥI���j��r���C�B��zq�9�V?eN���+TZo�����~|�&��χb��lz0.z�?�պE͖{��4�ϵ�	�i����LIa����W���t��S���?-��O�����˫�!���J����:��a���O�_�~|0:�S��F�2�˳:�M���ѻ��m�nu����bFr��LO�/Y��x��$#7!<�8\�Ccj��o9�o���q�Ј�.h�T�;y�&,M*"<`�} �L]]����z��p�J�x�x�+<���k������s��+.�	�>� v�%��Q����̆"+dSl]P��6���	Qṩ�f=: �L�:ds�85� ��ә�@6w#_��y�v�P\Q�l�l�n%JP�jGS��Bj6�����X7l�Fѝ��7lm6`[����	}[�[�R��x�N,`uR*�x�1s���(�J%��K��a*<e��.���9蚽�(@�y
n��[9|��5���<X�Y�n ��H zs�+tmЧ��7_G9 �؀B�ӌ���pxzKT�"�Ha�g�{^�o�L'�����_��g��)E5���Nۥ����hZuؙ=%Aݘ���/��>F�rF^,��`��͸B�o�����zIG!+�%7L����BXN�4(�]8a�w�<Ń&���"�>	���5�T���0j�/�U��08�UBV2tթ�3C�*��qdH���/�kV����ޝ%��9����H$�`����slZ�q�X?��~𖾜�� J>k��������g��������K9����0�z�[o(�	��4.X��'�	''��= ��:q?K�aO���4�&�Q�	H�`(���w�����v�~Sseo�	� ��Ͳg}xD#J�8����c��=]0AX#Hl�`�c��Z���D��bECG�R���i�z�0:z���]m6��1�i�ł��7���+?㹿�S{�k�"׬���x6�f���\��).�D�Oq��ϱ���A6#5'�����`|�$��B�G��m-#2�Rs�T*�&u�֛o�=���E���s!�����K�"��o���n#�\)غ`�����x,��FDUlr�S ��ȳ����i0�|�ff<�N�5�E3�1�<��|5�{BdU�������.gT4`�B�	R��d��-��7C\�+��
m@��Q��).!�e��}��:�T(N���Q(����h\T!2ڙ�ԁ@Gwzt�|�	�TU7��|r��L�թ���q���<�Q9�Ե+:72�aB�\�׷~@��TG>��P_�=���\?�^>�\?���z[����[G[;.��u����� UΕ��n��w��@V����Jwƴ�#�G��m��)o�\!A"dd. G��@�D� yoŃ�pܠ��!����T�����]�@��K>�������Ǫؚ�{��i�z�g��m$��sFJe]�lo��#��Ղӫ�^y!ccr�׷X����V��C���'��:�sB��Ob�(���&k!��6�`�Ɓ�ӚE?쯔�@��m�C�ǔl�X.�`F��C�Q_��wK1��;d�a�v�т��;�Q�:ǻ.غ�/��s����PX��$�njк�k�nxӁ�����{���y�e|Ծ��훸�7`�Xѣv���UZSM ꄾF�����e��  Q�ut�D="Wl~��Q������]�`���r�a��8�0gP�	��h�hM��P���L�BY*�+���P+�'��J�V'S�1ùsAg���a� 8��&̚�YD�ٌ�$0dDd|<���ߴB�:IED�H�n��vf�b�+��YA�`���J�@؜�� /�,'��ڊ�r�"�b�B�3z�,��~��P�+t}��BsZO7WN��<z4Ek�K�Ѡ!O�8���3��[�w�	��
a�ς��fj#��x����"�D���Z����)E�t��z�^���,��xOm�6���<}������_�-�!��IQln�ۺ���:G�r���N�"�R&F����i2��Uy�
{����@�ϵ�N�S�$*T���^(�f�l((��s�[Nei��{J/�3e]F��82qWLޝ.�Ƕ���j����]�\̝p�%�^�J����P�9�n[��ޒl���rap%+n���_���_C��W���HcC���s+��ibˑ�����tSp��{ĳ70����vp���O�Zk��l�2���ߘ74�'2��]�t�˛K)�%�h�t#!���G�	]�C��JX�к�����&�d���
��N6�h�hҽ�Ԕ��/��|z���o�'\�W�b��sW5�Vچ���u�t%)N��iЅ�OQ�2r���s|�Y��#�ɠ�n����hE�J�qL!	��g����~�i������o���� ����4T&�P��X!�n��X�^�:���NU�rfs��N�P������9��t2m@hL�r�����y-�M�M�)��Z*�m�oP�L����ؼj�O2ť�����[����� 0Y�NZ��>~�I��q%���������\&%�8􈤁�Y�&u��mhP�E94�w�z�� �H3z=G��D�Ll�g��'X�@�؞P�[$7A������,*m}���u�� �o�/^Z��ۊ�:�)����s��������m�>H�kBZ�e=�Oq�?W������R�ѻo^�G��!�NX�OT�g)x�_�-��� �ڞз7��Ջ��ta��7��4���#f�T����3n���1��/%QT��@���[��|Ӂ���1C{��.�UI_y�	� �گ��~EU��kk��2�c/R ��z���%�8����ɥ��*9�u���P(1���!sZ@T�Z�����
�9L�^Sю7��P_�(�	SN1�����7����>
�f5ցgB�|y�5���A�����'W���0o���Tl�*�����}�t�mo�XW,� �pU�"�UmD��Y���*!�F �^�D�Ԋᰏ��� �%�h_/0j[��"Y�N�DE��`9��;z߻������=�5��FWkœmZg��j~�J��ֳ���U�z�支��V�b��k3(z��J~�ݨ5� ,rX0z�:H0%�Fp��N+F�="�ؽfa��C�ʚ�*�6(��cR��R���Ũ �~�� �0Zˏ��@V��M�������
*����庁zGc�d�AB'��ijhHk@5+jjT�Ng�9�t�����N9,��u@b�"�������u��8KF�dϑn�!���sC�J	w���q�C��P�Ů ���Ӗ���U6P{���/�П��X�'�j��-����7X�>�N��>w�U�}�X���s�7�8I��S�}��U=�:8�^�z��)W���J
)�*�6%徏��{K�=�ih��M�x�{��R"ڡ�f�t�v�����}��}�� �W��͂T8\ng�F��u� (ڡZA�H�ϐ��6���^W2�,�hc�à�)-ÎhJ3�e���eQk{]��3��a����+�Ӓ�i�S?���RR;F|9�p��0��*��d�`�:`���FN�y��Ë�@�x���y���B�+��]�e�d���!�}NP ���8��"=[��u���u�<9{qQa�@дa���@���5zF��du�Hq��¯p�U��t��64����gT� �8c���[{��dR�vs�:�)>*��d��! ��׾yk�5&�����+�y�F/���+�(�q:�3"�����7��+x�,�o�n[S���������Z��)s'�7)ˬ��H�$��A��ۉ?�<�M%��pBU��]��
Ō��W�h�
�iA� zD�oW�l�A��A�|�z��N�/b�$ h[Q�'�u����xOV��a���1Q����`T#i���B=��G��@%��d��Tq$-ȵ8�S��*2OӨ��GQ��k�:UD�ӹ6��~��QHgU�$�������|hV�.�<?���[�4h��}���� ]��+�nX#�g;����0��'3�9)Q�"f�b�5��&d�Eq�z����<󁎆�R2�F��t�F[.�"
�F
wju���(*���L�"`�&�;i�8u6G$�Ug���$	�:��P�z*Ղ�dnd��Qε��Y06ul�	�	�{�C�Gk�oF�As�-��ذ<DԜ#j��1�~�PD�/�تs��Ugn������B9j��&��Nަ|Qn�M���ܞ����G�x�y�Y/p�u�I����l`ݬ �/\5�s1c���a��醆��l�����*���1D����_��'����Mqך���}'��!M���(Y�����c�J�a,���	��K���}�q������9.�(\mNr��`9�ZNX;akFw{]-�ۚ�DֻN����hǶ�/��*��a)���Q�zm�y�Ԝg�� ��y�C�����n�(�w�k��f�5uj�h���~
*?���`~��^�^4�D;�X�?������������T|>�N' ''�q�i(��#Z�hr[�h���2��a��#�����O�����L�����8�}΅3?&IM1��3�=�0�S�m���ѥoB���6��,` M6���>���3��'�������z�v����
��u�X�ڝ��c���ѻ];��T�	����ޏ��1e�L�F���ӳ�7������0����rA�ϐ~�����{���D�͎��o��C���g1t��ɓ�E�fsS�&Թ/L(]�xGd�Z�;S��������w}��V�6k��+�snL^�{6���8%3�0G iؼ�8�)�d�I�eZ��x�	�U�b����v��`x�Hd|޻���:���	��:�`*"h[б��B��rE��[6UP!H�·&V���4}���7/�s��Y.�1H.f�u��/h�-:@�-@)SMA��!�1̀!�]s8'�Gv:s���ڬMN�ރt�27:��9R=��N�D'��(f�A [�>E�r�u�!�-�
�W��ݎ:�4��2�X��"(�)0���:������:bJ9�#��r*�O�<�.�.ש@P)�#��^��#(��VeDE ��N�
���lx�:]7�ј:�I�@{�<9gy-��P�����#�@����rD��9���z�	��=Χ�L�:�8� b�̓ZtD�B��y�kn���]P�"�����u,����B�+��g��P\�|�7��5\޼�	���u5c.��ʨ�V��m�d�,�Ϝ�~@���O?�g�>nJ=�F�g~]�hO�HI��N[Ic���s�(`����	爴}y_������'

>�ƽD���`�<��ݬݬæ��$#r��Vp��H�H�1���^�nW�^��}�1ZW�ϯ�u�z}��x_3cky#P2�!A2���7�p����ޞjrI�@��Q=ڧj�[Þ0a���g���h� �N؆�}��o��8��M��}�5`{�5,�� �`�c�>uUl�{�T�T*V�% `��M-m{i���
�킫nX��r�"2���M*��:)r^6� �g��U�=� [���yn*H��vW`l�"Q<4+��%ۍ��ݻNQ(Ie���ܶ��nx^��J%�Z,��<GF���ɸ�;YL��'V�^��`�
wDME�:'�9"�@��~xr����RG����[�E�K��k�Hv����h4�1P���h5�U���7��3J=y{����(%&�m��HV@����@����Aj`��	���c��ڤsxR���_��b�U3 ���������pB��޵�Я.S�^�����B����ր�!W`�z��]�,`|��_�}�7�^���m}ݬ�:�IfN�"W��Ϻ N�q�F1�Q�{�)0��h2�����fyJ�>��αWL����������~��m�4�TZ����#-u��)�V�i��i�#�3��_RH�l&�`���'���F�:ə�\�pFb �TjoA|E[?��7�D����M+.�'+��x��� �?�� L8N�&�g�^,v4��q�q���!�ʱ��ا�}���d�!�&
�s�C��?�!�?kD=\K�	`�Ć��+V��j��

0�d)C� 6�.T�Dq��U�EM��8B׎���'yT�o>K�ɀx����'�ݱ��_1��Y[�qs�\�@_�_zL�S�ۖF{���@9G���{������%��;����
<oƿ0Ё���u4� *�xA�hG�M�w��x���<�@���C��H�lǡqE����c�K��u��J��i������70X7�� Z���؜IU�bI�{��=���b3�9W9&C���Mz4c*�P��T��EU�,��ͨ�H�"=셭����%�猼Y� �*'�,6.v��pwN'dk�q�H$�LA�ۆ���7�V
J�3���z��u�mE׎u-�����5�����3Dt�>%Z���
T3���=���θ�;������]|B����D7�zE4������D�ܝ(����@��9.�y���<��`���H�Y�:��p�	lY�E��*�+�������A�#F��l++�ШCP���7�U�/op}���4J)�}�z�ڻ���؛��hIF �t&�6+r�ۚ���ꕂN�p��gwrǫU�w�gm��� � �8�gH��y�q�$��#��-����ݣ����l�\��3?�ay�C=�B�mOX7E�ŋt4�@��)p�+6l�����.];�V�����#�oO�dÎ����S�n9s�d^˺�"*�*�h"ن��E�|$/�MhR�;�fhZ��6��H��+	�>{��u�xz^q��{�a8k��$w<Q	v`�Z���:Z��fc�;���E�P�Aey��`߶&�A�C�����2����@:���
J$����8���(�kcE���
���m.�g����[t<i���h��Qt�̷H���{���֢(����E/i��J�',>hMF)�N��X��Ƚ��^��>R'� ����ʶA��f�K�6(f#i�9SNy�`�^wk���36�Ƭp;c]:�n%W�z\>�׷oPT�ʸ�}�δ���zE�]P����x����l�뛊ys�b�&�#��؍v�Dt�i�<���>(�]F�7��ؾ�������\v��uk�N6�r�Ń���]2�+i�1��8����裳mS ��R�#�Ք3�;WOqG�^�{�u�&��U֯����h�ety���7���uE�T��]!X-R��#��BHN�*�#��'CRޛ�Xe�Y�>)���-�O��� #��I��)"�ؙy�G����"�_'/|�@i��*B���T�E��}�*V]�;p�
����>j}g��~�ju�l��:�l&4:_��8$�s�+mt�.�O����kG�l@�/�w�Q�TGof^�P��;�v�<gJ��D��M�% ��OnZ*�)eC4�e�_�+bk�ѵ���-�0�#�q����V�aU��wl]�MQH��F>�+��3�מ7��o�%���8�*��N���\���Ly�"�X�#�:.�h(�����U�éKm��ϥ����hs��.`}kH�����X	��RFR/�2��ΣݿW��l�3�_@��ܖOT��O=��ߕ�6��|��F���,b�C�1(V��%�hf�\���(��Jg�#G�ԞQ���Ԋ�H+����ס�(���b�aU�`������ \Q�(/V��l���>�m+��NX��uC��|��i��m��z���2��=�O:9�:4�>���{Ę&��Y���9}f��iD iT���II����<�	V�GD�q?�:�~5٭�ŋ;&A�Rk�C1<�L�&���M�� ����H���P��}�m���ذ�5��-�&Q#q2N@� U����'@�"���=�}
Yӎ��Vo0#M����3�-����VF3}h-SԚ �k4�S�<���.��qB��=p�9t��Y�����Q��ݼ&Q5K���tM�v���.����*'\�׾Z�I ؊����s�J2�G�~h�Cx3"��Z�t�[.��V�:%�,(�9 ����ek��̧����I�����z���S��lQ���o�B6`@Ĥ�����ņ�(l�r���&�歞�h��Ώ'ŧ�~�x��R�)��]͔�a�������ԛ��E��^�s�$��k�p��@:�љhR����Q1������֙�0C�N�h�ܽ�ɹ�<r����[�����7ٶ�M�3�����cT�?�+a~f�i�B�ר�>�ң������3��gyu�C�uK�j�q�VX)I�R������m]Q�G����Ӳ`SB_W����Y}r�)z�O���h���'�v5^�-�F v��q���*�}�7�8��p�"�KcJ�HŎ��k�G����9�p�kc��n�|x"f!�|��a�H���Qw(F�v �R�)����
�gڜ���W3��l�z1�<F�`��R���;c�>cY�Z	��h���W�2��kBS=�|�g�VD$��צ��N(��0Uj���X�r�w^����E���Ǩ��T����j�Y���ȧ0k�hF����������g(VcC"��D��'�4���sdv��S�s�s7v|�~�6�<�c�6��k<�Sz8���-��y�zBG���G^��*��=2:Ӂ�ZA\�1z�dd0��p%�R�z\� ���r���,
?����W�K)�L֢e���;���"�ދڝ����;_e�g�]�{A�C�U�ZpN[*-�Gz�X��
b�͘aC{'�Ԣ�;���[ݜJ3�An���UB��;e����3��Y~v�iʢ�렰3���>A`d-���\��o�yK��p�l����k����{�ضRB��\�u3Z���#h[�Z|1*Z,Z�1�Y�n�j�i}���
)ya��S� �w�9�k�N�~"��Y��I�K��#9�=�B$I��Yu{�y�+�=A�ã������������d��5;!��U;��\u",KM�4����fr�ά�Pg5k�J�?�瓳c]��Q�!R�)��p��
$$!v2>r�79����:�C4���}�i�U3B
\w����������;zX''H��/�߾��v��p����qe�צ�X�_�L�TP���{�p��**�ӹ��0 ε,݇�(;ч��|��!w���G/	�⛟��܃�b�9��/��(k��&�s�8�k=}�D;ۻ:{t��Ϭ6uM"kI�����b�GN���Ƕ�'�w>|�x���0:���_; ��}�2`$�y�宋���<�
�\�8�X��[��~��	�V��*����f�[uv�T�����yad�R]�K�S!�1`�qpn4��=�[9�c=0����i�1��4����hO����[t1΅������K�?�
S�_��]��?��f�Sx1jYe����p]ַ�D!q�Z_S%�T�3 "ض��̸-N���N�N�;�`�O�3�e�kh�42L����b���,��`��{�.�����Df�O�32}��A���N{!�h(��:�r ��XĈn���B��ƀ����<��T1)1�?k����	�Bu9��/+�u�i�ц}k���xof#�E	�����+�ً,���X�#{so׀\^vv�abЍ��%όm���ΌzF�:��X���=�2�+`��eF�kְ�O�C�@��\*�r�Xk[�xLAZ5'#�a����v/�2��{kY7��G7y�I�������	FSĉ�[履#��)꜍ݽ��D���q��b֐���F���}�ӁOc���fk y!f�X�U�{Yp����
�טߧ1�B�X�;�z���5�!�8�G�E ��=�EyF��9��8+(
ubN7�bx������$E[aF�q�������^g�]'���ܸ?�=����@9��@�lW���͉.���@��}dlpB�MJd��J��qǪw���io�ڶB�b�v�@a9p�h�:��y �l�[C��Ō�f���d�-z� h��H�Gn�����0�٠��u���b�N�����G�QgS���=�b}8	�:�;�p$�H#-�4;���kĲ�R���:�|P��Y�\^`�Ҁ�#����cumDT��tA�6<>��ȓ�FX�{#�����ʾ��!a�>�������(v�zG�-�_��j�9?O��!�����[>�/�������ތ��E�6 %zh}�l��*��x�+
*��Q�@u�G\�)����$6��]'�A��E~S~Ky�)����3;6-�{R��Os?#�Q������#);X���'urVH���'u熺�ִS��=|�58ѣ�"�N�X���(Ҩd����DбΑ7��Ý�6S%��6�ܽ��2�mj(Σj���g��(�	��`D��v��ՋWI�n�'NŐU[s�h3�mFZ������cu���e3Z���T���^"��D����
*>���0T�����������2�)qA�շT6�ZAUP���X퇰b�}�ذGY,�V@A��Y�7hW_J��	G-��YާDtzɹ��M(�I��Q��lu,}$Ӛ�2 ��0hZ�]�?���o�srgh��=��!SZ0{j����7���m��Y��EE]1~��ʗ�)GG�Fu�v<=]QJ���ds���� l�7-%6�V1R}G��(���	�|˹�������$�6e��gR��ְ�`����c��_�pA ym�*��*gŎ�!���J�y��3��jᵙ,�
1�\7�J�/<���39��􊮴�jB��HD��J.����D��,���dq�=�0�\ϑ�9@d�P��K�s���ư�]p��>W�(�n
��e�2J�2j{ѓ���� a��h"�?�΍kC��3�y����G���(�ʳ�^1������;3���-T:���q�~�Dge~{`�-���ɻ2B��P/Њ����w:oq�ُ��U��S��+8̤KȽu�������z��5��ȿ6T���@�̤#�.θ#���jS��DֱAu׺X�T�S*
��}}F#�e��tr�Y�h]aL�+̰Oŀ;�gBG�3!�߫��Y�7�ى�����|��%�c��ĵ�:M������H�#��\vNǄ��^�uN�Kbסǥ�3��O�km�b���r��G%�R�4��,"��Ya��] �?� �����+D�?�QСX�8�"Yճ{��:Ȟ�E �9���z���v�غqZ'x&�!��"�}� ��Ө�r�3������Ɏ����ع|c|��F��+ht��)��	%��lchO�~FEEe���!��Y�����k�h�{�U��&���� ��z�#Y�]*pf|��l�=�x�2c���Y��ӛ�T_�ݑ�Q�������0�>�n�.X������]RaĴݮPqs�/.��Po��?Ԭ6z���E��U�y�DôKP�F�-��BvSu�vKE8�5�2u����2W�n�GXgB�Y����V��A�)}<��P� v�(i�BV��yĮ��J�w�qԭj^��f_6� �v���3�T$��!9�0�V=��x~N�aLR�a�_����߈ '��ƹ���O���q��{��3�����ڬW���=�b��\�@�X:��Sk���mPK�:�1����h�!CβX��4E@���n�/v'Ҁ��p*Tu�%l7�io��N0tM��Ri���H��e�_�S<�p����b*7'?^�;eb����n\c�.{7�@���`tP�:6����g��W(*�U ��j]Ћm:�a�>�&�	~��kh-K�ة��ܴ;?�S�ŰG� ���Jӽ$CɌ/V��[�/"=���O�"q{C�peJ�_�v�L@!Q�9�A�����C�c�|m!�D�aRm$l��EpXA���&��`��?ZG(ׁ\i�lnuN�b�2�!�k�@�:�BW�4�W"�}�����`����9E�~��制��{䮆Θ�7x�a�a�VKZ�L) -��&����M]��3�A��[��-�����)�0.
�&�������)[���&��P9�sm4*��4����zEi��0���r' �G�""{��
vN=D0��l}���zH���J�]j+(u]2l�Y�=el�����7�k"���K��h)����o��?�t֦6�� əR�eM�3Yx'�B���A!��TA��T�x~�n7���ޡ�c���{1�5K�$��@E���S���6�x>��G���Sƽ������B���tDZ�%a|�������3*�U�r(��@M��r��4x9Bv��m������Q,2L͵��X}�|N�ޣL�Z���* �i཈a�&R��Z���64�C=�������lR��hq����?`���iᮩ�~��_�]��ʬ�&���Q�p�sgOt��p�\� ��s7ex��������|��&��T� =���hS�1�1h��n�]����!�a�"s��ØZQF\�-��7Fc���K:���h}/��������ޙ���"����H�
Y��"Fܐ��a�S,���tϣ��xTw��<B )��q88&�p�������:9eq=Z��¥���vSR�	�*��C��b�������xE8WO�	��N��$����V�fb�؏{����{�{��`_=�	�� L4�ҚFoO���X�]��+Ԩ�/%X��!rsV�~E�(���\,�'>a]7\�+��+��y�fuA=��HpI�2�=�w�3{#{�u����3�����QX���榰�et0P�|KhE�+TW(�DHc����8[�P�M��Z楓]z�a&�1�׾��kN����G�z��� fF)D
Q��EP�BE����EQ£p�c�t��_A���L6�!��@z�T*v�uN��d�(�+�	�@�pw��+���犃�4��0N�!�`�CT4)�]!��w������ �� �v���
�QyA�j�l*F��FF~�̷�X��Ƹ�y�݉Rd�X��(�����J06Xq���;�k�W�ɎG��?���;����r2g\'{Q\x�ܒb�b�����"KR����h��w��|�|�At$#��;kp[��1����y�4�/�-_K@2��2�|��u�.(W0�u����]1:�U�A���P�ކ!>Th_e@���oPF�f�T��5[D�\ݓK+���1G8`���N@ɴc�Ƿ���Nn�C��e�{&��Z|���IϿwtti>�h�TF�6�vу��oX�뺡7A�n��'���3`-�u'g�\$<��u_���$������ڞ3P�q68�3�~dN��
�>��
hAg^��\���q���F9�����A�~t+�w��?��khl�KJ)#�6uT�ʐ&�m�E�bJ���9]bV=¢�d�i	;�S����kG���qgto����B
M|/�!*�'c��^�/>'���� #r����Q>u��x��
i�\v������XE*/(��|oX�������N�9X>(S@��Hr�A@����ɻ�K���e�s�	��N�P�ݪ��G ��d�B�H�P�
��s�5P%�t/C�ja,�`�֝����ZfJw�f�Q<�ֺ��I������{��#�?�H�?�C1xǮ�ńL�=��p��ו�TPJ�p����@���(�6��t2(u]�PS����}TFߒ��DL���-`w�>٨cB�w����f��q�;��RHS �ņ{*�Y�����H����+3����j�~{� 5����k�P���i98��;��z6G�Q {���O�����}���2�hu�4���B��,td�y-Q��f$_�, ��lG�H9	��,�cچ�ܑ��G{��i��U�V�~ھ,��$0�� �]�ć�
zj~���0�à"�ao��W�3G�s��8�)�;d�n����ў$q8�u�q���u�T=R@��F��J$�(�	�q�&%cn"N�C��Rt��(�o!���m�S�*�����C�Js ug|n���z���u�#�#�L� �~Un�B�WE�������	(�r������O��.}��U�/�ϐ�ŉ���w(�c�=Z�cY<;�q=�Fw=S�����Q�P.P&h'��oA�Q��yޝ���D㔎�gx2Q�<;�v�]jfT ��dw�S>:�G9����2��'>#qCF Q��^�}ެ%R`P�.o�v����ӂ�*����e�[Jźٽ�N�Ey�u��zu��,��6�o�Tx��60���uO����������x~��u��۞t�di�m�l6Q��+d[� 3Z*��ܖ�� <R�ש��&\LoG������G�z��t��!�rZY�f=�vY�=�E�Iޭ�,������	�U���b�����|DV�zz��Et��U	���-E�˃9wpq�ˉY�B��5TI��Ü�F���hB5�3&���K����p��{ւ�DN��G$` [�� A��٪�_É�������E�E]�U�yY2��8x��=x��_�ϛ�d�o�ҳ"�?ؽ	f�
�ޞgU� ���e�1p����o��WhF7�KG*�����j��{�D��޼b��(�ؙ���J��k���#6��)�d w��ą�6�e=�b�0N0��c{�c5�,i��a/}�j�=M��ٺ[� `F�D��m�Y�����=�!���"�����@ղN&
��ȏ�����cT8;s���o1��U�^��gU�R*��Y�0���+r��Sj��5��s?#�i�H��T�Щ\���f��
B�>\��1DH-c<�X0N>�mr��Y����i	��S�O)��gبy�>y���)���HTP���X!��l���B��:W/:у�<9�f^����(��)�>G� ,�t��ѓ�us�2Ⱦ�S��+TGaBx��U`�(�@in'�{׻�Ez�b��A�#�M�%��/ZMjDV���ǁ*T�Z� BJ�9%�ݞ'�G�ad ���}N~�j�,?_I��T!�h�u��'��5�e�>�2֏�{����#��$J���B�=9�uc<�y?23V��Qٔ�Am�y J���,ŤS'����B�.`�!�׽IG㫡l�����ȇ��hɋ�#��L���¨ѐ�{/�Q��U�S�j;�����
'��R���������vM�ɗe����^�U��b��"Ppj)4"	�yB�����!�G�yr��3?���n�i�\�$U������;���8�w��v�?�T��r�'�}�ea��6z����b�z������r�(����Ʊƴ�ӂ���j�]�E�ur('����K�ND�z1���q�P]��snU�c���~�D���c�p�%[��
��sC{#��%�.��>Z���A��Tv����fX}��d�-�r�H�t�*JN�BǞ����Z�n�n����-��0"�o��E�PVtCl �A�������!����E9���-��ux6����aΛ��="˱�aPF+�0�(�4�Q3�H)�`��R��=�l��E���sX��m#J4"t,b� �	_ǭ�G3X���
 �V��)�H�1b���g(G��u`bp3U���É��}��C�9����Y'��>ϕU���^�;�؞[w¤M=��M�2�zw���\�@�l��ȹCt�`OV�(6u"���5O)��8ס�2*�<z�;^z�3�)&�]c��@�o��o��b��ENЙ3j'�j_{]��
�5��q�
�A��@ݠ�`Tu��1�;��L��g��C���D�GO$��Q>��vK��/^4G^�a�3-t����{�]K�� ���u�tA���O�6��Y�2>C(}Ak�m 7P'ȲX�{]@T��.'�[4�����̎�]��U=�GE�X3�[c8� �w���	�sK��s�P�^�F���;lV	�i{F.�K�[Ѹ3I���vvhx���l�ehiP�Zlt���G�o�X�d3����6P���A�ѣh�l�������`��//�P��D/Wb��I#7��m��u�Q�8A#��|�c�L���1����;��/j�0o�+���)�����|�AP�$ƿ.`e'�]d��`��E����N�)0�N����G�kc���-f�V���6g�� ��!
�j��co�:2_�Q�'.�|b�!"#:�mI�%�(�Q�}�o[�'ӹ<[L��jI��B���2��?;-\VurJs���;O�B����U����fY��{ħ�t
��3�#S3nh�t�|h�
q?r:_�~F����Zv��LU����Bϼn���C�=���ƝR���#�����+My��5>'΁�)�#R��3��k�^��'kY3���u�)/��
�܉(�X��;{�ɶ��m��(˂�,�Z!��bw��/W��e"��3�c�ݎ��r�����@���;>lZm��A��� �~�T�?$��Fٜs�w�v�ns�{:f�'�GF���(�E��1�9���>����I���f�IFU�$���((*�WP����w4(��0���l��B���8�܉Bo����q̥�Wl����yq�n,]~s;�sˌ��l��f�΃L��;���3��g�1D�CW8gT��I�/�F_R�?�<��~E���m\��UD�/%��&f�:�o�q'�6�� b>#�*_w���vg&���?"��7Г(���)���ǣ
9qdn�P��w_��0��ş�N٫�Έ���s�&�q��`�8:���f���s�i�i� S[������m�D#}ـ���,�P7�T��
��E딒s} L���N�QR���q���4��=������	����I�f�!�w���*��ED�t�S>Q��Wmv���b/�c\�6�3:Qje�n ���jƜKF}��=��0������C��:�[Co��a�#H��]_���h������%6�A��@��E٬�,��k�A�T7��6� F��İ@���X8�%��sDO�l@�73@PU�kSH3X���ZE�K��s�5;�S�� �VvBI��`���ts3-/D>�����=��X6�r����i1E�C%��G��qwo�;D�=��M���Ӑ�@�B
���������ܔ����W�����r�a\�uν�;����Տ\�-���9�KQ���D����`D��}�T�NF�&�r���$'��dF�a�ZԸ�}78X�BG�HU��'&��P\'��䓓EJ��b������5���e�>�|�`�06�p�,R��8c�t���H�&yn5�J(���A�6�Ċ��8��ts��,R�W�i�t�*�3Й�}�p��3�p��#�r�NU�;���p����E �,���	�V�ɀ ��-��Գ�������[[Q��. .���[��s�I}�'��!����㬏����ry)B���y�7��7F=́�Pv���o�Na��N���B⻗c)8k����S��-κ}5���oH9r��$pn�-�6eY��u��2 l#�I�,����Ñ�(9U�*�����T�8ˊ��[,8�dy��c�n�+G�oB��K� {��dnQv�����^���^�;���ѣ�?N��".ಀ�Z^�#D"��U1D�C����_�������չ¥wE����K�Y�g�F�7(�z�9��T���ڑp��A4���ܻE:ꟛ�9*���^�Y�Q�@:�&��(�Č�uW['����bѢ�D٤����-RB�P�ec�"��F���D�;	Ԯ<��n��o�q�xN��i�?/]�H�JG�x�^�JΏ�GG��g�5!�ѻ�#���.�@�4%Y��ᡝ.�qYܙ�;ڎP�q���]Nh��Gbb�7ϛ���X�1)%D�����F�{�A�B��
mV�ޛ)�bP?�x�y��z~�r:;����ఇ�����9��o9��CP��Š�NjU����zءk5ϔN�N������I��91��@�w�=96�ԣF��,d��+H�,pc�ͳ4t���es hx�tA�v~H���}��o� %�o+D#/hp/���?�}E�y2%��8dcJ�p`�;A��j��~3f������;����#�sO0~��t@�G������g��Xȶ�)߷��]����+�bdEkB�F#p`E��H\	�s��P�����fnQh<z�؀��)�,�=p HrwMn+����,�A����Y�!
�s��(<)#�d\�00�R�� "r���	1j@��;�NםĂhǴ��B��Vɬ(k�#�n؉��0�@CXZ �6���)w�X�w!K�.����_4N�8����
��p������P�kz"�	_
6����3Nft�HGۤ��^��c��^� ��ޯ��yt8G��v��$g�N{�*�%��2�)Nxޛ�ZP�*��NtO��^�Q��ԡ��y���D6b�{�Fyx@=�@�SI�=�_jd���F������@t�z��)l9���'Ο��EpH��n:=f��3�-4��M�T� ������"=;������d�o�Da��'FA�CdF!��:`k6�k X����_�I��Q��n,�ЮoѯO 4s��xn���r.��Y+h�x5B����&�s�5ȸ7�v٪cy��͜=�/#����z� W����|�^��	���<A��b0C���h����1=�\ׄ�y5�� ���`t�:5�O b{�D�&G-
)B'G;a!q4!T���
h�iX��k{���tV��{��$��\�xF�7va��+t��Z�ڤQ}�8U�IG*-S�j���y=��-b�id��%�b}s��XW.2�E�3W��s���$�PBF�U��SC��}�0���	�-FD1$qj+T�)9�=
�
A+��*tWh�>������
����VW��N�fA�z�C9O���]p���e���|�fԧ����tgT���9���;M���<(N�G�55	��
��]-�Ĉ^�&1�)EL�Dњڷ�l�Wo��HS*(KO�yt��ڝ��wH���<�Q��&'�z+�&>)�ߟ�#���ǽϛ���(�w#M�@.s4Gؓ������py|��z���l� RP������k!
8�rPq����RS�s �U�
��hJ����j}��?���*Z�W�.�O��o�.O߷>}�(׏�킢�	d]���@OڄP����s�ݠ�r���<G�V������g��2�q B)%����{>�q|�[ͯL8s��Ul�<�4�À���yiFO��D�q�}��Du��f���"A����r�n��H�[���fs��@!Ik� 44t]mp�Ѣ��u�]�MȨ����!�<&e*�z>��i����P�4"р�vxʹ�,���I�aMF[K��;���P��E���W�w�����,��<#R�VPF$������1ʾ�
�T���ۄP�t��07���DԻ�2M��=e��]��5A�������C�"
[ZD<�o�_Nk:��z
�^�ItP�N�a�lvH�>뽓5�Z�t��K��:�x��p�:�Ml�촻(Ӳ����cG:�lq����>)T���Z�M/��8h2��b]4�^g=��2�~[4O�+|Џ�1N:���m��D�����P�޻��/j]tvcT]+���9I"���VR����Q��y��'�����z���F���9�j�5��DG���r~�������J�������
п�v������/���|���#Oo>�O��{��\��1]ߞt{���!?o��ʽ����	e����JC;A}��d3��l���1'�߇[����`H�,o{�Ȁ��������.7��mD�?MCvR9|�Ip#�D�uD
t!�"4)7$��B�S,Άf=�Pꝵx��3��#?���ל��.�:��P.<��g����x�#SᏑM�$@��F�*c����pnsf"6�X�P(����!.{��e�t�7�XC~f��x)Z�����M��Em�n�X�9E=��n[��@��&���J�����1ǟ��,Pm&�����
*}@���-p����9��v�������[���_FE�+�À�]����g�d3�:)�"���y��^#����0�Z�Z3���\R1��d.�j�E߼�4�ra)�����o��^b����9���wA�|����Y�3}<��=s�ߥ�i��DRc�)z�U�I����M
�U(���RO�`׷����_h���'P�`��?�����^���?�]�K�~��#���~Z#|�aŶ��?�_�[��7��������^�>���?��$_���p��(g[t�JW-:dT�igz�j��P-?`�K\s:D:%J�~�� @s�Y�=	�,x���=��.%��Z|!��Z:@شwʪ��4os��qx}	��!�b9�%��Ӂ����pbn!�o�5kj��2�PU�����\�^kb�1$����J�2?���
w��� e����	�D�����JQPͰ����/��>9�QB��?�������qRV��m�''���K�3�{_��!w1��>vM,:�8:	��w.�`f�zZ���(�1'�@��߼����%|���i7�V
��l�:�/�>^3��<H���w�}����uaAAcڳdb0N��HT!N�j�����y���T�r��ۿD������3R]����P��	�vW�����t�}��x��HV��4�-��<G���B�dQ<��� C�T�ڌ���O�zF==��G�ԟ�֪��
c9�!T�i������_�����<~�Ͼz�����?����+��?���կ�4������K?�7��ͯ}ܶ�����ۼ<�~��ў>�q}��UY���+�zV=�v���#y��R۫�{%uFRb�.S|qPǩ���L�(���R�7x'EGo\�3��Ľ',)^��A�4������?��0#����'�><ę�j {��k�ZYJ�yTmK8G����#��_R�dO�s.ܓ��>v�vݝyE�&A�؝�a�͞�DCJ9�9� !B�ځցnSkuR�N�6�e�������g4�w*�1��:���s��FP�mP0��1B�?o��I�I_P�Ӗ�$t/�p���<�����;��);�r�ɀ�:	���>rYC��wN�S�0���d@���,C/��;�=䥵8f���N���������X*�3��QWq*b���hR"����r� U(�	�t�����g�j��7r��h3l�Nr�c�rf�ˆt�uLR�i�{�R��a�u�_��O2���	�d�p�5���Ƙ���h=2L����IQ���R�����$�QR
e��c��T�����>���_����/�?�����?���|�+);7����#� �ſ�����_�����O��/����^�w[9���>����+X	�W���b5̉5����������z#�7��~􂻇˪�GE��D�����1��~��vH�ה����<�^��=�r�w�E�!��$�
t��	K��N4"t�KAQ/|ӽl�!Mo_=R�� ��qs:�PC�h�fg�%�~�8���N��1H��r�y	3�-�ށ�['�ݢJ�A�*�l�h�!@CF��Sňt�q�7�g��
���& ��4�����������'�3�^����2��=�]�m�IRd�S�V<\|N�`ϑa�aIMݟ3��mSq�F���#��_��:ݿ�[߿�������Y�����[f���t��QjEe���8�1��
F����vl���z:�>,(�RC�qJ�L9��{�1�#苑
Ǻ1����9�#�	�߳=G�!��|G��K{�x���Π���.RǄPN�G����z6�}yQM?��68��I��� ?���ß{x��\�����?����s?�����!P|� _/��z�����	|�w��_���+�o�r+��=���w^��+t�@H�	mӺ!*��<mB��#��iCW5�[tp/��ţUo���A2��������U�����=?z�zI�T����9�Y�~�D=BG@�{2�8����k��c�D1��#:�< 7��6�x��X;}�1�P���L�]Q�x����`lL������v�ݻX5/x�hV��a�l��vJD��T� >�G�cIk�h��O�R <ߋ��d/Ϸr��}q�������^2F�Z�k�6�m��H�v>���=�4VJ���HE���b�tPPa��7�oQCA��Hόvɻ�à�\D�<>�Z��c�{����0��ϰ����;�\����E��pH���-�T|0P�`��������"��(��z�R�sJ��C���Ngи�X��71��ɩ��O�+��h�=Y���Vd�&��S����X��;��Y��H�I�(�lQ���=����јhSV���a=?��W����?��_����ӫ������F|�t�t�h�?�=?Uŵ5|���6�����>���~G�X�w���կĶ�d�C�LΛ�����:S٪� ����*�A׌����#�q[ݗr�A�q��T�z�."�D��������g{љ�`%77�! ��g*��@M�N1a2V.2o�ݴ��ˉD��p�V�V�A�d;A�nS�`����!��Z�_O{�y��c^j^�DFQ�H���2W7\�w�</����I����&m]�6��AA�^͂�;�TLn5�$�S! ��1�jjSqGGG�����ar�g��m�F%���D�><7+�w$��#���9
��@�wV�6�]@�ԛU�������耘�,�ؔ@�Iǉlx�*l���a�����(��{���ؚ4���iy)ʞ��^>���P�{	���QkHf�[�>.ڊt��Jݜ���Ή����h� ��S=���H�`3$���J�6�E ���U!?,#�iݰ�!ϒN�4��f�?κ�^ڎ���{~�^�A����(�?�t<�!r�g��R� m�Z�^�zBYΞ)٩Hb�D�E��@B����������|��_�G��~�7�r}�^��}�/��~���M|��}<��gN�����imu�=�#��U�\�a0*l�}�T���!��G�0Ըɡ���xV����S�%����g�i���}�����͓��&6���!�=�Y�� ���FPAǆ�q(��S4�����+� mP���Qu���tX�H@���M�S��^�/�qWF�T��k�6ѯ�.F��;;6���#�04��fp)˾�ɨ���)�|��� ]��"�ֽ`�L
铧̓gޢ?tLY$Uk%��*@&�R����U3P��$^�T¡�z�D�w��"	�EgErV��x��;�{oc�-��c�Pp_�r�A@��>nq�� �'C�O�r��6�3�f �d["I�:l����P���m��MD7G��r�sQ�X�{2zgÑ�P��Nʔ�E���\_�\o�z�A2�"h�H�1�Z@�T���t����`ش̲�.g+]�j�iT�q�Q �BNe�����6��Q?�U�F6�w�o6&�����nF/&�7������I��j2":�Bs$��#C�d���*�:�Ƞ��drp�����M�^���(�>�X��>>sy�3�S���4z�S��s?��O�N���������x��=��c�W��~����O���\��W���r�����y�j������
�
mH�ԃ3zuJ��F���3���guzg ��}��~^͕�Tޥ�0�;>Q�z"��X���z�ҧL�� ��3΂,��{��� ��I��	�n�P��5�<N�r��i�������Jґ[rJ�=Vrxw��dx.{�~�y?y��c�^��έ_�R�������hTk'gDa\!��;=�˳�Agi�K^�;d�Nt��h�`��뽧LmNw+�����)g��Ϯ�5 Z��Q��S�;�4�F���Ƶ���]^�������V�Qйo���:�����c�%Ekf8���:0�Z��UQj�
�@�@��6���v���zGa��m��X+T�M^�3;�KIG���ڼ��b�^Xs�ĬD�ǹدW~���@��ⵌ=$/��;!�x�ՑU��F�b]I��Ǜ�Z�r��j���>l�-2G�������3��������}"����o�������2�-�x|ϯ�!|��� ������WUdٸ�����#6Q��bסh}��	�ä\@� j4��͌�X�{0����ctH�����f�Q����i�C�@�(�N0��_��"t=ٷ�����;�����KE�� uQi,P#��37��(��n�tB(�Nc�q����a�윪���)O���Sۣ����@X�U������
��XUU��)�9�V�*���v ���1a�����r��1R���	��c6�#�^4�p}�Kk�N�Df���zWE��[��JD`�AHs�QM|�ji�@��@�����%'�@�cO4O�y�x��������I��M��ұ��]4�b�,�H>\J�_b�;--'�DQ����k  {�IDAT8�)�R�S#��Cl�+��ST���/��h�q�bOj����9ǥ�Ss�z"�'�4ޕϹ���7` �w4���8G�8�� �re;W�bRr&f�*��F/vV����N��<6������?�����k������mt�r�_��?@߮_xx�ST7��V�'��p䛍9Ǽ��R�%�bԆ��)⽩]�Ź�i_��z��W\�{���qϻ���a=K��6����@�"7:���1�wy�c�v�#���&�3��Wv�u/�Q�wQt	%�)���ب�B�J��ή}�qǺL`��JhΔv�&ϯ��cjRBw��U�*��x
%j(L2ܥ�<�Maμ_���@Wc ��0h2�S"�I�Q�%t/זb�t�EI�@��|qW��䱘c��ˆ9�mޓ����	�4t�
��$�ĊW���%�G�~��ü�H�O���/�GBn0^�,��|�
H��L�R��^�� r��·w=���_��@�	����G'��='�G.(������|P�U�;�S��hC���lNz��/�����ebv2�{Mg����%�ِ�8�i����^�(�=ݞ�@����J�U��4lV\H�-�DF�����j������������|u�����
������xz|�p��t�~͏�ķ$����6��/���/�g?�����&��j�簾)��,���
���c���b��4�0�+ȩ?4�Jx`��|w���<F�d���� �[{4u��߇�C�d;4q��q7帱�*Niy�yVA����ޕlֽ ],Ci̠3�AL���o����ۜԢ:_����d�W��*�{51[E�k���H�n%�J8~�
��ٽ�euF-���;<�SC�<�C���f7�6'R%�,|�k0.�r�i����������;<�q���A��=��\H�U���p��D���I��=:'���b��Ɂ����V�E��`C����隍�|��*����,�Ѱ�2F��ɽ����l��B�ڣE�@(5�A�Xo�9U�K1�7��Ҭ�X��f�
pq�ݲ��s�{Z{t���<�[��T~+Ծ���:�*��)z��0�]��<�G0���L����cׇ��	�щD�R*J9���@��zYD9�����[ey���������g������5����: h|ק��?�������"�A~�n0���
1:��; �������ӌ��Zl�o摂�{��+na������`�o�1U;�Ӝ���=e/Գj���A7�(#�.^d����o��
�(^�G> ]�Ό�f�}b�QL#��.0x�&�tvL�6�ca�U��W������{J�4��R�U":1�k�쎟&��8�e�͊����[�N�] ���3i9���F�` ;�y�q�#"�=�̕D��f85��ǘ�(���Qr�q�*J%&�IՊ�^|L��=�3�אq�7�ywgX�����p�a�c�8���E�����7f����,�WW����[9�/�ɼ{Q�;�;cp���D�y{�:�f����ާ*��]�Jo��r#V�JN�$-)[}��5а���IF�]�e܋��2q�8GGv��;�:˰��n�MQ����$"�`�0�׎.�;��ہDEJT��#���c�ƭOlF��+�<������?����/������2���;6���_���ÿ��g�y����/����/��� ��[���n���;�
)S���O�WOաMσ���S�ӵ$�o�ncX|
>�[�v����4���k�홆3��}�0�&�ɫ���A��D�M�)G�&��� � �^R6#���͍	[4�<r�0c� ���R�ESTu@�3����r[�*�m�@̎��E�J����/� ���{��S5�
�ym��z�X7�eSl�8�Elڔ�s�>�`�t�P��Lh
d�vvx��1�]~g������(��HQ�v'�H��{zN�Z3�9���c'�N�t+�$o�;����[b��YC�l
]!w|�o���Ao����Qp_OS�_P9�5's������*�'�5
̣�h�+�!�8�����hZ�:����#��Uw`C�H����츼q)�,�H�:���,�Z�@�	���������"ք�����HA�� ��i��ApG6��ɩO1p���/a�o���>��|�����F�μ�=:�����~�ٿF�0� �G�LՌy�Pf(��� �������x9�������������oů��t ���u��O�5�3�������|��������i�=]�������w�^�X+B����"om3�늫#��ywod��n����6�n>襛�`�1db��,U�}��w;�<[#x(�P�0�,������Z�`!RXn��qH|`��7��1����y�~������aW�E*��
M�k��(����S�,��o
��U} ��}�<�x�PW������]Ѥ�ڀ��X�b�ag��9ڔ����V�nF*����g%�:9�Fu,�L�0�2�~�4)�5�Cs��(��i�]i�<b�| ��UG@ҽ���p����;��m��~~U�����BLA�������X��n������	Zރ�����,}�M9|�������򏜴)�a��m���Q�����WdUQ/3�C��ԋ��za����R@��h�B)F�-�љ|��*qw��9��V]L�ȟ���%Qk�"�E�a��aTp�!}N� L;YO��|sDC�C2h��ٹGd��=��I�x"�ʌk��Ȁ�i�*o���T�����&tdgj������\�d�I�sDK�
*g���W����㯽y�������S?��ߚ޻��t ����I���/��_��^_}��U�~�_�����~-�3( @�%��P�[�3d�=g�\��3
�o�������s��O,��zs�[O	��{��0�?
����P��#<� 3�1(��p�`���I��X�&O���,D6Ioҝ��P�}�G��1m�]�
fk$�N��v��0��\��
q�|#�V��Q���5!Wx2�k��L9l,YQk���l�"�BCfW���5vG-��l�Ս(ᥢ���A��Ĩ@]�rXP0s�W������Bچ�6������98�Ű��M��DS�v��d|���U¹p4ϨO]n��6G/<SzG�4��	�6n�!��3��.X��9�r��y��9�Jٙ���s�����_�d�����LPf�m�n��$�N�n=r'���L�i�;�2�,�����PD�/�^�og������g}.�-��D�3u/�6 ��\�_�������8p��r�B8��s
4	�KB�\�����@��BkW|�=~%�_�A�����i�>>�z�~���ڷ�E*�hW�r|�C�p�[�l-]�S�4ra�M��%�� �����_��ѻ�'ŋJ��1G���hg2��pX�]�4a�-:+����d�[S���ם��G.6�;����fo�b��x�*�l4�4w|F N���1Q�qM#g�{Cv�i�9uq#u�a���Ju���s� �֦�4�&�8-+[�%MF�����9�4���`�{�d3���c�(����>�W�v��9��c��hh�d&��7��"5!IC��K&�Q�x��{�����WH_}���]�Ќ�(y$b͐g���
��Օ|����2Ҍv� ��?���O�i���|)Ĳs��u����ñ�~alw�{�|^8uq��z�y�u�̗��N4e�32(�w�sv]Y��������dp{q��T�Ӻ�3�)����n�C١g��s}  L�䨲�C���c��=��j=�=����3W���r�����hCگ��5i%O��,B�ji�@/�<UPY@��%�ğ�������?��}������Wl�����	�����u�ׇ?V��GD�?�}��RVXn�X����
g�S��@�����2�\a�1HV�1�b2�����f8e�!_��'/�F��3�/�r�����0�{��q�C:���+��tj�ϝ�$�1�{��V|r�PA��K�{���s-w��M��)��v(T��鵻H��7 �{�A\3���W1�T<�#�hB�n��*X{8#�7�7 p�0R�ժ��͝5F���Z��6�@La�$����|�Sq20z�w
K��x��/&��[B��Q0����:����E�w���A�
��q��������<:K�;hθ �������':���n�#�Y��Ζ�I����$RK������
=����qxtȧ�o���N�6!u4Г�+�>�<.x_�0���*�Y�>S�:�SD�:r� �3��u\�/F��pz�d�k\�����B �(�0���V�N㭺S�g��wQ񌀌b9�qu�`���X*��<��l�K)V��S(_jI>:/A�GC}SH���L�1�l��r�3���d�{��4q=e1����zz�7���w���*n+���ǯ�A����o�~��տ���U�?ޅ~-�P"��&�/hޝ�r������&43V4��!�՝�=�$�6yn���/F(�{��7��S�������!�IHTSk4�;���t}@v�?�Z`2�Sn��L���W�P��8Eͨ����ɘ'�8�k0I������&�0b����o����Ús�1�Ȯ�5+��lk�h�6�"�+�� K:�F���x�G�~�UCl;u&I����k�0)���0\�p ����0���㛭P����E�� +{��ۮ^���.9=�&�m6��2-|߅r9L$��fA��ơP T�T����؛���4�Y�u�L�q*�B8��i�fu����M L�_�C���ʜk�`,3���X��k���
P27-6��{����H^�y�F�Z�bC����v���G,���+1���{6DT\�u��=C[�st8���r�3Z
	�N.���ʭ�����M������K�D;��{/��C>]�a�r�	J6�	��i�+�h9	��_ZN��'*�&賟ů��Wՠ�����.�-��C�����(~����R�ђ��&��w̥���/���z�ɽ�c$"�㩴�@2�x���杇IJ<.9`�Y�)'�vR��0��#
�C$ޮ�0r�$�D-��3�N,b�U�H{4~�O�"�%�n4��Eq�\�q��~U��ppr�o}��aBe��?����؋+����(������ڰ�-&V��r1Gd)x��qk�W�ϝ���$�]��m�������}d��es}����!�{e�;9
���'��f�U���]G���b�c*�$=2��>�H��n�
�hv5ǈ�#^r�tΜ�J6�$`q�������~��ŴV��LeZ*����ϔ��\��>g�u������~�F��n��A� ˺T:zQHS�1�ǝʜe��<U`yx���3tk�ۆm���,��U]�D�&�B$�Hh�Y6�Ο�p�����0���a����i'>:㳃�x_d�_�{�{�a�{��Q}��x�?�ʲ���.��A/���߹���?\N�oן����oů��Wݠ���������Y��]P�$��D�?g�1M�a���8հ�.��{���J�lƬǴ��]KD�M�"��#e�	��1M�{����&%�Gh��w���(�1}���# .3�6��&s)Ōs�9݅&�k�H����gT�֬&DV.��.�E:-hq�B��P����Ǵ�4��k2T����fx=����鸏��4gu�$��m?} �	P�S�^g���	�W@�2�
+����=#�
����yDP�R
ά`w�p�3�	�GdtB��l�D���\���A���1�>R���ϕ:�jr��̋&�к4wX:������tt:�8���D�u��FDsxJ���ȏ��N�i`ҹ���D3�����!ս1pٍ�m��@���J�o �N1j-�`k���H=΃�cbdt�E�O7d=}L�����e2�2�"JE}�^�`���a]W�m��A���;�j�iL�.���6��C��G�2��LE�CC����ռM�t�3ՙ�{s�s����`�p̵N�3~T4�h����X��\+J=��
.%i����s� ��-���x�������~ ��R~��_u� �����������k��_����?�x�qR��k��Gi�*�2/�Dl�='�f��ȹ�\9kU
���{��vo66/<�1�2({
i��̚q�S&��( �)�3 ��Ǜ��W4 �h��52R��iE*��V�,��x�|����v�*CdC#�(^�U�bɫ�TT<�{��%��3m|��Ӄ|�Bw�aIX."]�[��k��R�F�!9U��*[YA��nX�׉!ڰu`�*��@��nO�������(�8~�Lv����פ�8-��2�Hh�ް@_�p�$��#X���L���hҊ���{��:��3�RW�:�^=K �v�`m�.��P�(*0s� 2N�
��6�� ���ZI ���/ � ��3P�"͇	�!DP-���Kq�:E��@]�~�#�:���Oy�TA8{���ADܐ�jB�����������9l�AM����m-�샙l��2N,�4�|ƹT@�*ضo`�Zh�X�:d�D���r��a���t��1|�����";*?f�a���49y�m��&v�Y&�<��0�k�0�i\��/o5 ��h�>Ӝ�*g�ogCP�,8�k���Љ�"P��]���������~��X: ����C���_�y�c�友�E;��唹F��� e��q1���DKC� �Vc�#~�a���|���O_E�FD��VJ�N��d�%Z��]W)�B?�4X�|��G�Qe�H����[F^Z::8�EYD�u�C�ڰ�����xd1R9�a�#q��Zs싺�{Qّ��P
7�.p�3�#k���X�>9zc���`��Fh�]���J�B|r.uW�$t�*������XQ����<H~Vb���
�m���;B�{��X����n�ۺO����A����ށ��n��)v w�B�
�qD���O��2�)1�����y�d�����`�(��4u��[.�-{�����{��i���	Q��A΢���>�&�;�x]�� -Y ��y�Ul��9�x
ʉp~�@ߜ �P"�z�Њ�4gtv�ޱ^�^ϗd�d,�ps�����)9����mi6DՈ�DB�vw�x�:`�ӵ���A��NS*��I��T��՟g����W��|�������[}�c3���G�o~[oW>=�;��O�<��.`�@ڲb��\\�,�I1
T
bXTl^���{�I��}�}�j�W<\�	uŉ>4+M��<�'�NcL�����[�����Üǁ	UESͶg��t�ϡ֘�dF����}F�k۰��E,LL���$�{��"��%z�^���zג�R��,��w���7�7F�7Ի#(��fQP�CiT��]
Val=R4
5u�ϙ��nl>%pF\c�S�hI�����A,5��&Y�:�w����g4�_rA���&��)c#
(j���~B�BnU �'}��+h�5�ϛ�C�=�h����8�2v[62a��됋H��C7�dv��|�;������t��}D�"á�b7�m�cFa�h�ʔ
`z����j�2��V=�T���S��a���l&K1��A�ay� }�F�$�e���
�*�&��l�~�!/K��3�я"w��J�o��_H@�df�AȊ8M'�H�x��dDȔ����`^��Xu;U�؋s>?QY��e9��'�y=��[�����͠������[���|��_��?����h򛣚�,�H&�y|�8�������mT9{!���a�^z����5�>
M�OR��ÃӃڑ0�4$� ��wJ�	���!��5����hD��������n�& !�ްiCG�
�P��h�
P�y@����[z쭝+@�e������N���~��P*�A�ɫ�cm�`E�5�����4��	:�D4��{�<�%���C�����m��@��;>���V|(�a����A{eA�3�'�'�L�b"r���ioZ�����!�{�F��i��qo�-}���_/����� l�p�>.�f�,mAP$q܍�X@.�RЉ�!�)b��О}��m���8lf%��sFn+F@�H��j{8ڨy�(�L1����pPF��B�` zoh���0�8���[CW-'�v�b��+zP��|^�u��8[qQ{�>,�;�������!�����R#����SR:Dn�sd�dx�z'ӝ�|9� "�2p��?�/��G�\O����p�ys��'����[�/�D���_y̻���x>�}�����|�+�+Z���B L�ژUt��L�����OPr�.�|�DD��c6�s�����D��y�!�Js.*%���V�^\6yʉ���3v/Sqe�0Y�Td-�/����sLe�v�N6{%:�����������=��ð�2��:�Oާ�̊0�b2�|�~?����1c�P��l]�|��(����1��i��S��O5;��Q��t��r�n8#��2��fx��9����-u/Y�]�����Um���~ؕ|�l�$1��C�Y	��nn��}�jv��\/���6��G�
ι�|���v�����ɨz?�,v5���-�߀9'>x�<�Ǿ�\�Y>��ǽ����f��^������3Mn8#_?��TQ,@�(ݣ\G���G!͌��	��n��;�Q����'uQl��m�W�$�(��Tf��<NAԋ��^�i �K^i����`6��{�(�& ��YS̓O�@*���{�x
�E&Ƽ, -P��ǝ��ᖿS��������o������oK���?v�N����i\���v~x�����.��$Ҡ�-g�N!�YU��b�ȹ�(�k�����!�����t��A�ȫ��j��T1���A�|`:�r����3^E�k���.����95#�(��n����Ѐ�=�ǀ��4/�i@o�l��t3Ӥ��+��PeT����Z���En�q�V��,�^5�mJW��������v9�a�
��veFA�O�o/�u[ �ص��W�(�Xv�R���N]�n��V�DL(T�(J`�1��=m�\X�S�^x����*���eT��
j�6�C�(h���u�O���Y�w���Wˡ���[)!��A��¹�1�ƴ���>�=�Z�M�M�֗)!�8;S�|�U�Wh�o9$�gG���丅�G^����"룎�}2��@+�,�
��7HkPQp	G�u�s�
��q�ܮ!	�X*N$t*���7x{�#u����N!�����{<��#'՘6�h@�����h�c��	.��֙�uǣŞK��}ܷ�Ǎ����l޹}���R߂�O=��}��	[�~[r��<�����#?U�?�����l�[A�G՛��Y��A@L��,֩Vй@�8k
AVC�Lw�N�&{�b��ｲ���D���}z���y��!ǎ�v�lv �Хa��U�F��Ū��U���A#���A��|bu~o"g5�@EA�>w36_}@��f4��K
��`�e84�:�Z_��G��'PTG@��%VQ`mT�O�v�(�4��U�u�7��u$7h0.t�&7���\��O�/���o���{��l��B�ʊ�4ǅ�>X��^N�I�$"��HC$R/�SD�ٹl��G����������k��bmˮ��9��{�s�[-�"�H�D�UC�ɆaAz�yȋ���!yH� ���(q�8�b;Aذ��U9��P��I�H�b'���朽ךs�<�1�Z��[
`K��<>�X��=g��ךk���#yj��$�$�@�:���z�A�·�ȑ�B�y�E{�k�ܷ%OpB�m@�w�.��F�o���p�V���3���	�պ��F�ͯO��٢k���S��v5f򜮨~>$g[#0����� $���D�}A���A���A>g�{���1VD�{~�x͊=�{�����܈b�8h=B����o�C�U`۬o_�~-����jΞ[�]o��X�y+����ސR�hO^���������`\���ɔ�8�Q�)�;��	H�o����{�ӧ�o��]���|St ��7����3 �oӜ�
R��H�(�S��Y�蕚�b� � ��T�+G�d�z�����=���V��z������jk�ppxԶ�0�ȫo��G��Ͻ������w@e�,3N����$�W�A�c��X���z��+��
ؼy�H��!�[En;&ɦ@��gߝ׼��X���#$�֚���RoTo# �@�R����t�����r���㄄Rp�ͨ�!�����w}u�n��:+�C9`H��f�k3C ��isŔ*v%!�l&��6�m���ka;4®`�yd]�����i��{����f5�lMW�Yĵ��lb�$�*6^9ۺ;)�xBZ���Pb2�%���#]��=���"���z�a�x{ UF��q��+t}���ovK���%qփ��f�0��QN�V���f*�O��x�{m���	�#�� ���
���~�����Gћ��=�f�(�h��RF��(�6^C�" mH�.*eE��K�ǹ�:^�E�y�<�=�/�ނ�̣R^�У�ϟE*]gk��)�g��j��P�:�ڈ�wAu���̄�9�~�j��kZ�,h�lmg�3BU�{��Ϙ=gkQD�He�i�\~���'�����w>�g�}��i���>�/��G@��w���P����.���z�S��Y����u=�H6�ΊX�0�vV\u�}����<?�e�w6^� �J�uz�6�z3\�Tp�`�����-3
���e[DK���n،��o0�/t��c,vX�C-؜-����0�����*�9��}ޣ!�P�t���(��F8�-�ko_�ń#���s]�k(UsS����r�ن��D��K]���_��[r�(9��q���ѥD�P����F�i�;z���|�*X[nVw{=�5Jg�~nܗǴP����9��nc+.,#>$��Q��d�&���0[�^��0�.����Z���z{�z$B7+���{?��}��v�z�o<�}�=FNx�����e�_���>�U�~v=��Y�Y��X��u��ݼ����
²4�f������V�Zdu�d�9��mޢ��kŸ*ԣ}ԍ醡O��̍��j��k@�w�U���ԪEs�߭׼?����w��FPO�l?��_�fx�{�������Y��\���v?��5���r�4��i`�sB�T���rE\����3��^A�w�,�i: ��=«_�,T��'�?)ҾhO[Q�چ,��7��g�<E�Y��U��C]�4vcn���l-��}}�R������(W�X�]��������;�y�ɍ|��y�U�4,*�;���O[�<���������V=��&���Ekn^-���H�ҲjcCoN���_,��ݾ0ڒ t�|D4ܪ�n�9v/�z���Y%�����Bk����o���I�T��T��^������HDP&h�=8B�q���=�%+JR��:�=i�д�Z�u}���Sg:c���\�՛ܬS=�����ޓ�C��{Y��Mz���6�³]裙�7_�����ڸXxT�,"▛�3?�ܘ	�@��Wj���q����^�g�7���5�H��;7��Y��lk_n@m�W�V�st���[��lv�8X�c�B�E� eF{M�JFJӴ�߿��m��*���<f,}~b�״{���o����.(�'���c�����v�G~�����V#���Z+�#\]5o�Lv�����o�O�<����Fa�����ϕ�U������a�y�C�'��G��l��c���x�\�8.)��!�ݟ���r�Dx����7�o� ��Kb�)�ť��B�M���KJ��b�m]25 ���=n��ᦛ<2%h�X;7�{����z�ga��p�ж2`�������g���o'M�}�\a���ϓV}O�uS%W�S�!�	��u�3?[�*
ۃ��{*`�OC4�_y����Ln�Kkr��Mα�m�Ms	SHm��,Xj���ൄ&��ӱ��0"��X�p=/ :��t�ߡ�5�	#wj��ke�v}�C���A���{c} �����%�b��}z�iW]\0����#x>���8YΝ�W����_�
uc̨�H��R�Y��RJ�G�W�
�q���n��|^-���5���Y-C_���nK����@��F�˳N�B�aw��~�i9a96��K���r��M�K��!�P�I̦��Ƙ"/2�բ-�V��Ix����MM�#������~zc♉��h��������g��r�#�����CΞ�.=@�3M����<LV߰F����)�a�t�"m�P.P.@��\�Ly��D�"��/~�L���s�~/���W..���|/(�����]��f�Y=���*��@#�8���	�=�)��B}�w���r�k�n|��}@ȣ}���gS�zhY�Ko66�����7ӋlN�{�je���N�Q��g>ސ/d5˔i��>�9<��_�{M�����u���h���m��!H���������W&_)J���$����1�<mk�r�f�������6,�۠ɼI"/ SZ7]d��Z?pv��3	_�{V7#���k��L]o�Y��_�.Ȅ��EX7G����K��u-'P��z�^�LxUIܖH�z�����t���=�n����m�����=�k����'^�@���0�G��|�v����������	*e�[�����E���H���њ��\��׼������X�_	�d��"�Z+겠-ER����,�ݣtM\�P��2_��l"�g_�\�>��Pd�c"q끎��nu���o���)o�k�M�M��`�������|�l�7j�!YtJ�s�f|vA�Jy�4�/���SϽ�C�����|�t ���_��G�A�����(�zഘ"\J�Ruo|-8�n3�(���77����c�<��^�&\���<~jͷ��Ϛ
�)������f�=yȳ���U]�%lg�w���ga%�l�=mb���j���3dcWW/�7勈��9��=���������3��[�g5:��7�����&�������P\����4����I�&�j��
[�Xl΃E:�0ڼ�-9@M#���X`sK*�0�i�R�z��PzT�_��d�w��7�n
v#�~�V�C���M�ϥ�V�<���C�쇆w$���<c�W[�q}:6�v/"�?�̣m
C��("hU�se���M�E�?���r�����A|�N��ͪ�a\oWjԺ
ed����3d�|6�EE��N�,f�]a������۸
_��kDz����D梣���@��'BK�^�]W�j�ٵy$}#�ؿ��n�i���3}ܬm���&�cݳ���g`Ѝ��Jgn�*�k����f�|m�I/R4�=G�NR��5ev�JY���1󟑺,x�xCt x��n�W��֝�_l�?B���Ԓ}�J�jT=d�'J�����x3e�B��V��|�&��_��^
�}H������i� ������"7s�����p-�9�|{��Z��Y%_J#�:z@�?$��0�����f����>�	�L��>Jz>���B���M��>�_�q�}
��ʞ�2�M��[n�}F^�?��@�!>DVA���6<8Uk�iu��矂{�m��Ms�uH�Zn�y�O�d1O!%7~�`Y��%�A�庯Q� ������#}6A/�qf��C��=��HX�Fī(�y�D���tow�3t���&lFC����Ev4fh���u��ߪ�m�3�?0�זM��Q=��~hml��8������0Z6ѡGX��7���)�G�k��v��+֐��>� N
i3>|t�̋�f9����Sf{����Jƴ+���n�c�įA����z�R��lv'���t8E��&����$o����u��{��u����M�v�e�Wt�@m��9�F��>vw�l����ꐽ#�[��7�Mjek��1�}
�$�dav�l9���ze.����OL��J}C�s�<��r�í8��+m��?���-�Ia���B6�O���ΐ�M��%��@h��5�|�w[�لf�-����X�HCLHc���o������r���s�Y��7� �'����������SF/��;��=�N}������-z��ՠ;*��%��9�6 ����6*N������~h�5���	��W�ԧV��GkU�a�+k�lc��#2� -�tif��x����z���!%F&��8�A03�ZaS�D�B�s6A��@MAd��T�\UܛOk��<�m�t�����J�m*s����2dh��h��6�:�B%{'�goS�T�*ZO>1-C�$s���5�	=F�%������6
�Z�Z)�SF˄�Pջ�� q�skuYX�ad���=q�#�	
~P�z��3b���:[���{;�y2��+Z�F��$���X�Ao��{]�� �vrJ�=�������z�5���x��x<b>�����+�8y�G��� �12��`=�b����5�2j~d�Dg��x��Nz���gz�C�i�fk���b�]������������筱�N������d�̉2ɟ儔
R�����"����o<��|����;Пx����_���~A��~��OQ*,O��U�BR>�F�@�!vb��	D �E���܆47��o���t�����ۙg?5o�0��C�����zcaZ�N�j_��H`ZC�}ZQ����=�&�<f}k���N���ڇ���TLrec���C��/����ԕ˺��zЯy��
^�`���x�����͙�ޅ��U@X@X�z�-�i��it�{���[x��'p���W_�7�/��M%7�T�z��4�HlmhW��hk����GPl�L;��k�m�%�s����d\�����c�;7s�7�)�����:"c=}3fx{=��;�{h*eU�+�k�0u��`�(�'CϿ7bHJ.����5��Eic8Co�Y���q���7��*{��z�;{�d��ߌv��H�l-z��GkЍo�����l3�N�������e�jg.�i���=/��`'3��b��p%QL%Ck#ےim���0��n�9=���y�wQ���=�M%r��O?����
���f��MQܸ�����{���#l���*Z���\0�(����iw�}Ⱦ�O+�ߎ/߿8<����F�� ���| ����g�_TF�K��!�4MUN@+X{
=t�d��zA�`���3o��{�#F�����d=T=�=���F�{l� l�@x�E�CD^#�	麐��&^�m����(���7���rֽ��N�,n��fL(�bX���ׁ�z��9�ǉv�m���u�m;�u��%ll���5������긯��Ud�[�j����iͼ�:�q-�)����	/��9|�ޅ{��z>���0��t̨}^u��~��nMVcbՕ�Ȕ�{�
u�YU���VX�f�?K�=�F�_�q��_������D��&xr�zJ^p�Ѵ9���u���:�!xb�iy���:&�	u�u��:�_�M���2���o���#i��g���腐�P��AX�[���	�m�7֪���0�Q�&��Q��8��pA�i��eF[��lW��g��(��
"Eʄ��F�21���*r����tkA�mRghc �_�GS�ۃp���p�t6��fG����it���/n`f�Ƽi�>nO��ɏ���ޒ�t�b�����wNy���@y��g��O���'��[߃E+�}���z���_~
ZT��A������x�Q�
4�9n��U�wk�&����dV*�-����8��G���x�`�/��w?�W\�eUA�}74ȨF�����t�Y�~5r� �������2�V�V���V5 �
�K��bu�B7�9�<w�#�:��6E�g`h�����	����^=�ؔ����j��^��@85�q!4u�X��	kH�H*�:���{����k���]3ж�-5`C�Z7�2�*�&x���\CQ۬��IHv=�m��-kps�b�_3�'�z�lDf��������g���}s뽒�>�+e�J��{�����R�{�j��ŕ��3*%T�ژ��کG䚎��z|�.����c����a,���9��YMVCDקWim�R��@a�x�W|[��M��B� ��6S�Li1�ͷhc��GJDP]��9L���vhˌ��R�s���Aٞ�B7X����u�G���q�Ekg��fxG��yx�-ճ��f����\����T<t�7�~D�3%8�l�R��3(O�����4���|�o_?�C==���{�F��o�Ї��_�9d0���禩�WJ���w/����n%r�m��H�~���J�����5�C��|�M��������}��S{�����џ_�L=L?���44,RQ��I3Fz�ݦ�<�m���S�=D�����2��k��l������::
6�a��<���ڶ��P�m�Mׇy��4�+�[*���Hl.UQxQW}ځnm�T�cePb$m�m�	��V=|�T|�׿���������H���	=�C˶^z��I��g-X�"&��k�u��]|�&1r1��Z+j]�JM���ȑ�����vM�������=rn���u	S�"B3��o5e7%���H+���U��q'+2��`�O�j�N�	���M]�Jb�)eԥA�j�^ϱ���<Ғt���t����p����X��mn��Fȹ�i��=� �E�"k1dJ�a?d^A ������󔐧r�[ſ�Y�����q�����P1����� #��#����������Cfd<N�K72S�Tv`&����/x��|�bv�5��^�{nz�ݠ����"M0�`�j�����c���34����Tn�O�<�-���?�7�7�@�����  ����駾������C�s���N)x���e�2R��̩�=�ښ4p^���V[���<M�[�*�y�f�g?��2��0V��x�iC�f:���E�s�.�L����)������@��w��{n�<��D�^K6�md�c�pcs��yN���I]�$�����i�!�����9�x��=���b��ko@�[��E�S��y�a1�F�bf���W|��	�64졻V�#���޵_���d���є\[���0�h��9N�	���N�!�2�}���2c��?�ߝ��
���{��HI��z$��W}����7S��o=�|ֶ�����]b4�3R. f$ʠ̠\@egJ��%�Ȼ=�T�4�h��]�8T7�1�j�{ȷ#�i���f^���=�d�w=ܲ
	�1Hg�|_��O�Zb#��cE-cm����>AXj��T M�Z�iF��3ي{o�GE�z�E�8c�v�7�n�6��e��I-����#qs��F{J��w`f,�y+ �׽S��=Ӵ���Í�����WV��H7h�!�kO��6վT�#��N�l�N�E��O�2��e9~-�����!�xS�U�׾�19��?W��NH�w�ȥ�"��x{a�p����Zĺn���|r�j������!,}��}cu��o�2�T�6�;�n���1tKY�&�!{��1��]�}zߺ�F��t�*���ER;�H�t����ǯ����z��d�a��x��iW��Hcx��-`�*c�&�b�ns�z$�o�g�{/E$\#>����ЅQ��HIM����+$'�4AZ2O~� ��yM]#�ߌxn���%���L�ځ��ہ�̣��c @�b^�l��1.��cch��}=��&4��ƒD+oB�#��G=t�b��O�Jid�m������>uʫ��C��i�&�T+n%+n圁��){4���g�$��J��kB����ͥ��V�ƃ;�:�J]]w��{�X�?�:�&���=��������O�m�j���*V�����*C�=,�!���*č{��UD��������ݣ��q�=M�\���58.ɚw�iY{���tG����U�-��~���7�O�o~�e���� �il0�C��Ъ��m-r�� {�sB*;P�~�S���� ����x��:П}�{���9 ���r~+��H�X��ԭ4���}�o�@j�#]�^�*$ [KR+�#��W���s�Ƭqtݱ��m�|�6�]�ݲ$�|zYh[=�=��{zQ���f`�{CX��]cX=
�եz�e��i* 5�¾Ag"$����LDA}L����vA��!�Vo��t�2vۤ�o����j���ĭ>�s�����Jk��\,fqO:5+�Y@�����`�083L��&1���e0+r��guU(ߚ=�/��N(d1���WG�1!� �wX��̽���z�ͷ�kߓ�XQ�d�:x����I�H#W޽Y#)���:M̢���t�܈+�$K�d�f�]��D&I^�h9��� M٢>�w-���ugQ��������[�˼`�ŵ��ͫ��}{{���F?n����%��m�4����>��	�s귕��WHպt K���S����TPe��Ċ�#�ہ�Z3!g��tlW}k�Մ,�c��xh^Dp��Hy�Ϙ�)\ER-Z'	@�>Q�ڣ5↳�BU��?��7�������a����^{3D��m#�2ڂ\�������$"�w��;��9�8A�
��r��\ (�N`ڻQ[@y��Ȼ?��?�7�����?�7Ձ �����_�9,K��n�JOr��ip��0���P��NԚ�x!ء�:*K{���G�������c����_���pc����YĲ	k�Yi�L��M�0i�>�O7�77������ɼ,�l{H�7�Q�L�F&��5ܷ�R��0�> �c}����5�%��� 6���m8�/�Nv�j�$~	��A]<a�:s#\WEU=������hJ��-R��y�x>�Ɋ���p�4N���*�f�kǆ��q�'�:G˩E⑏��5�QJ��E��k;������0<�/tv�ֲ�"�PuHޓ��i�l�����'���f�71�:�^��)!!�Y�F�i��^��̮�X.���R�.��*VX^�6�Zl�^X��t�Ϭ�$C}r�n�I-��g�����]��^�W����X�����ӫ\k`�f
p̌R\��>�4�h�v�UR��5ۏjkX*0�Z{V6�͕dG� �_�{���P�u9�I��E���5r3��#�Q���-b7�"]���=j�Q�d��^6��SF*djp�<d�X�4y�������t����w�Agq�����~��K���7~���NzE~�HY���h2�7���rZ=��a�]�o�2�����,k���m�cV9�߬�'76Y�hm.pϫ��Pݶ*�o`�y>���r��e%�y�͐t%� �V�:B�6�I|��9#�y���@N	3^T}x��i; ų�ÓD����5�{�!�l��彘,�^$�)2Ī�uV�M�M� r[<�A�J��`��ŕK������J������@�N	�^��
4��Sww��3�^[/���ӄ=�8��I���Z�:�����������>+�X�����:�^�u[���՝t�+�48�b�/��	>�N���SO�)�&9�5�~h+e0'��m��R�C1��ٌͨ0���z��A��g�y��������@"t��q���z�7�\\��Ū��Vḧ́�ך�_l{�=�$�ު���j\�J���r7������f`8@�V�	)OÐ�V��d3�ن�����u]�P<m)^i,zlp]��v��{Iלޮ�n�l��gA�m+���Kߺt��"������ϻ<��2��	x% R�(�<�ly#�I=�)!BJ�א��s����2�^���A��xS� P���o{���?��~�����|K%��M~W�̓���0��F�Эƞ�j��e{�����@�l��l����]e<�}'H.[�19{xh�gW�z_���
�0�y1��؄�Z�W�ZG����f.���X7��X3#b҂ H�$s�x�i&{���3k��!^?K�ٔi��@���u���:�6a��#^6�x[�sU y�V`n ��y�P������h��=�f���\�b���m��	˲@!�rBNdS����̣*��|�K��]$�W�����f׍y�z�c�S&�������خ_���[���ӱ��f=�����}� aW��e1/�<$��{�잒��!�Ecm�׾�\���@+�2��<	��$���,�v_�쨧��K�6�MX�/����ֵ�][�_;����@�/k�}���~��x�ǟ��vcٌ�_����o�=K e��6�~Y��� MpCI��n͢�Sbp���^Y,(@"F���ڈ��LP�H �)��M�3�،G�{(6?\1�q[�G�H��U�p��9ҿ�h�����8�8��=j�w����!�c��E� W��8O�#�8'(gP��T�<�R�0=��~2��+ǫ{�=���Q�y����~��﨟�9�����Ͽ��?�����"G4,X����C���IA ��۵J�ԇ���R�^/���O�6w��鮘�mB�:�D-�	�.�V>�sQ�Jzh+���R�2]�!�ILloߋglZP?_��IU��b��EO*�����t �4r��mU�g�{}�ȉ�h۞���?��26�5f�!Cү
�MR�Q�Rd�3��n��{���K2V�,��V\^6<)�L��Vۨ�ruh�S �U�d�3 ���խg�!e3D̨i,:��յ���޻�cܧ�g���ՙ��z�F�9��SztC��9z����~���M�A ͞̳�1r�������WkU�|4e@���zw�}-[�;�-���}
��]�2�Ț 9����ģX�0���y�\�|���q�����#i��n?-g��=6�k=��n�z��X��kU���4��"�%'L�	9%;�`�L
挤�T9	@�l�Fk�4r��CY��
z���M�B܈�\�H٣~�������zQ�p��������7�����zU�Yn����n���zU���{�*m�ל���@��(Д�����7�\��mJ{ ����ɟh��}���aqޤ�it"�~����Ư��q�����OO	��1�H��֦�^A����e�B�aH����#T�k�]M���C�7��ƚ�G��.[WF�yzŪ=�ݳ{�_�(Z��Z�V��Y�_���'Q�VJ�D��Z����3�0��t�6v�����"����)ﯕ֜��ٕ�n�9n����X�g�W�ۡ�s�.w+�:Q�M��s���e��+\���-S�n�qy!x��@� R=�n��j/SL)#1#�Aa�2RS�g��L4[;���抔3���L�\@<�6����h��q2���zR�b���M�j�7����Gd���{�CZe�EٚK6.b�֘�(2sF��BW[ߍ�
2�L�T��y���!����sF+tqt�.��y��@/�Z��wz�Q<�]O���zM����Y@���U6��d�{�Q�p��l�x3 s:o�!o����{�Z��li��~�4M`2�k��b�dbO�JV1�'�ͧ�l�*���*cؑ�v9EWEi���O���Q5�e��`|@�����ݯ�*�D7��X�vO��,cF�f�z=Ł�ߏܻ/w.�^�z:]�L}w6c���{p��yO{����0s��e������ `�(~���ެ�it CB�s�(�|]./~��<x����0��ݽ�q�k7�M!��湨����z��u������X���æ�lv�&44���%��t�9��#��4<�ѿO�屛��L�������y�Խi �40��v��`$O(��K��;�m�%v��IM>��=3*(�9�++	�������ٟ{� �:Q�W�JU���QEէn	�������Z�
hJ�1-G\��oy�Ɗ��ZQ[C�L���PB.�zf��y����&X��V@����ē`i���PJ��eƝ�~���W��&�9�f�mk�p�)*�zlN{t	MҪ7��w�Ev������aHٌoej���v;�a�r�l:�P�6��&���N;H���A@*;�i�@��'s�tq	=��.�8����Ji�n��a3�'7�ӣo�`$�\9��#���l���#2�kH�+���p�ѝ��Þ+��I�^���}�Wd��[=���m���b��n����N>��B�x��-��V/n�����G�9m���\�\zAl�
jd����å�>i�H�!��G��,����U~�������H�)Rqs�~�	�ŏk�EG�f��;@��kDJ��C��Ɣ����2퐦�T&�r���i�������S�����7���M�M}�w����s�(>����������K*�	Q����˧���9���e�ՕP��=r`�ʔ,TBCAZ�^�Yվ S?�W�����z�h-�R�ԳC
O���Gچ�\�]�F�����Ⱦ �(�a��B��@�)���j���[�	9�0Q�!gܚv��.pQ�8�=&-��9!��vJ�>'�Z��ۃ��d�ѣ��MW�z���am�{# *r�P�̌&�|D�'���l��{��	g���A����V.�Z��ǓU�i��3�
�Q���a���	mO(��e^���b��dnD*NMq���'2���t+cAc=�t1��}3|��^�E���t�Ve�*���E�x��;��}^wJ}F��NH��9���=\��&{b��кN�y<�i�`KM`�ВВ��!*�߃�'!w��g0JbdΞN�ϚR�y�<��7d��(�ի����U�&��[����Nڣ?�Ag uY0��=?SA��K��郡l*[�N�
�� M7��6�<��#�,H�L�`ڡ���&�,�V�'IR�tEj{��p<][$*O�i�z��CS,�tid�r;��?�z�9���"M�������[Ov�)�S�Z��E�v��6y�.��3aҸX#�}��+Fl_�}��
'���#�����-��:X��D�+�?��2A��\,���`���:�>ޖk��G����S�7�o��C�3�0n������^~��9ܯi��+𣤺K������|�%՞�@nM{ۅ􇗺����V����V�@�W��X���K��m����xo9a��Dmآ�E���ƿ�W;���	9��5�o]�@2#%�BJ�����[�`���T�����3i�e������%v(v%SvO P����=����U��>%�BA���H�_o�̬Tv�DBDJ�oӴS����'䴳��4�ݑ[���Z��¢�V�dJzJl=����`�k(�C��&�s<����&03��Ќ�)�J.���-|�Kh�Q���D6��� �	�+�d��'2�'�����б�������Ƴ�j����ѾǤ;����/xލa߽)����?�+T��n#]6�\lP���*H:���(B"�5���R&P�x�M�4�����m*����S�˧�r@&'�V��o&���5ZU��`���Ƭ AM�A�H9�%e&eb]�E[�*M�*n����������N|�����M�D���'�UIDIUHd�Jċܴ��}��.��0�X�R�)_�̱��� ��?y;��3)Ӕ��_@�p�X�()�	cވ�Z_����dެx�@�!���RaKM�}��M$��IU��u5�!d�(�5�;F��(���F��7������7�S'=`�=#��h��SA�%���r�;�:��ns�3���j�������\��|Ͽ�����?1�2: ����_�ٟ��˸������{�=��$���酪���k��+���q�����f�KI���ja\/"���zC8b�=4z��r{@������G����xiKtE'�zPTm85A�#�d�c����>)I�"��gMH�(^�iyfFJJ9`��\pk���t�|�|@!k� '$0)Zv�>�����������S#JU�-��DG"����> ½�t���!�'�{<pՓ�^K[qF������
9��*�*�T�lҞiwU���v��}-�:�'ngpR�Xt�@p�GiIN��2��e�t\x8N[D��v�D�����E#B*��pk���-­���.����yL��X r��k�ivD�2���MWA���vf����^�E���Y�U@�!��. d*����
��Ҿ��4%�\4��!�"������3v���O@�L��K��'�O�佧��̤��&�ĩ1s#BUEm�.�<SJs���r:��� >NJ�>щ���隠G �rﵓ��"h'-j�,`���W��(���p��C�])�n�����>�|	�U=�&��-mr)��փjۋ�I[+R[��L��$���"�T��HZPX�XG�\���).��)��@�KL��Φ�ժh�J��Ac�>TB����H��nl,��&P����=� �
�V�Aɮ��;�ױH����}���I5��u�g���)#�؝��*S�g���X�H��{��}�E)�K��7��v~��,�Q���w�9���G?���
~���=�f��˷ԁ ������+��q���_hy����m���<1��k�/Q�"%ki�&Hb�0i�N�:���*&X�ܛ��x=��hxI8������V7�U�C&`l �U`Q�PSA&��V�'�W ~�0)R�P�ȔL�L2�0�f1QA��r��i�;�ܙ�`���<!���VA[`�ښ��Y����T���<�Ӄ������5f�� }�2^d�<����h͉+���ݾ*s��n���ҔX.�����2��r��Sʍ�y.Rk���&�eB]
8=U�߯����wcW���������T�E�ITx�j���P�'n)�4/x���Ǚ�JΦ���	9eH3)K&����S�>+n���pkG�mFW"D���+����}��6̨��m�.o�J]ꛣ�^�lm�Ex���~��Z�.���. �Z�����	uf�(�H�V��݄S�q:	��)���gԚ���%��ٕJ�n/|�����S��#_3�Cb<,�����_�į xE��,*ߨN/��[.��[ޕ�)7�,�rc��D¹4"m��kd�e�&Mx7)�De�k�,�jEz�Qr��m�@��r}dL�y*iJ�K�Xu�mn	@Zj˵�,�%�9Km���V淋���R���|�H}mym~B��Vkˡ-ׅuIB�mAʌ�����q��i�����B�N��]ɸ�`\��КE2
d)�vB����hb:]��HPP]Еۈ H��u�Ż+]�����dE�"����Q�;��'�#u�BDS�;oM�{爌Z�q&�a>�@0{�>���>xe�R�#O{�2]q�-�������������R�9�-x�v���Ox���_�{��Oѯ�ҿ���A^�E�� -&�)&<Cb櫶il��R����D��dZ��\���lz�{��f����!���&N��@2AQA3�넂v���z�����+de
��M�1MH�=�N9{�3�JW�c���].pw�w����z*C9!��Ҥ�,Dt��&ί���Μ��S�\N�O	��*��9O'N��ʇ%]ޞ?�3?]�|��r��R3���֟Ih�J���n(������-���Vlr�js�L��'���������9\\�5��Y�q}��YQ�KD�[k���i>��c��[A*Y/��P8=��J��e��yλ]�23@���5��ä�ĉh_wD�/3������?����²]KοNە�9���D�`P���F�1Е�[�pV(�GE�B��:V��� �MՆt:i�_B�	����Δ���K�Zv;�ۇ��R�I��x�s�j��P%���y��SO�r��xI�o�i�Uʻ_W�/���
PK�%���VJie�qj<q�����7e��[,�"��y+��v��	�fc�T2���tЗ#�X��'kgj3P��5�S�L�z���Pv�L��Ί4�EZ�5H���P����"�a������u��Xj�3Z�2�_��m^^���h�۲�g��nk�����T��z(:CeA[ԥ�-���e9��#)���.�*{Bk��:5��m� ���־�D6��SS��' $Ӽ��l�J�#��vng�k)��0A��}��1 h����n<EYi7587"<%��Z,�;��R��xJ;K#��W����^*��J���.>��[�����-w��K���>���4�˸n����?$*���/u~{�si���fH�!��0���n۵b-�=�
�<�����L7��^ �ʱb���߱�l	�W�pya��������+�
����`E6jU��.�֐S�R2�2!sƄl����1+ Ta�
�|�C����%����gO�6����v�2	8w�_Ki����/�gSΟL)����IR�s޵��V=<�T��'>����z[3CiBK�' �g�y�o�z��W�
 �ZѤbYf���=�����^�ƽ|��5?|�Wi̜H[�Z+��L�-;�tGTo�����E�u߄wJ�������rI�3Cs��I�LXTY]S��'��Ki��T�%����z,,`�jR�["�*-��GA��L{�`�-�z/�C�T�R��fPv�RR�uG�}k=�ѓ�Px�&�U�[U�U����Y��ki���R[b�K[�R�)�:/u��~��ݾ�P3�ք_���|Yr������?�z�g����4?q[�p!�ť�|K ��}�SH�ۨ8y����l5����5���?���x~���  �IK���eF���!��m/����y��Nz���г�������;�����<�xWP��@��Y󤏧X�+d�RL�XeW��Rk*��tD=^��%��i����������R���f7�Y�t���A�0N��st���6C��P<r�3�X�\� `��X���/�6ʀ���ƞ���P&Fd��N6��],���H��i�������N����������Oķ� ���G��w��~	iaҧ����.˿�d����&�TZ;B<N*�y7��f�M���G�X��+?Yŧƞ]�.�^A�!�⣴�͏Tتe��ײ�ի������z}�Wu����
h"̲`>��Dؗɫ��r�dNإ	S*&/��g�j�(�w8L�qQ.q�p�������S�Ň��ʴ�r�ʧ	��=�_�����WN��i*{-��|���~���r�0��	���	w��^�w�RI8=8�x\p}\���}������Z�ڽ{�ݿ�w�S��,���=,�	��D��,hMH�uB�ɋM�D�o\1e��.�rb�2A�k�+Q����c�i��~�wW�ֻ���-�N��d�x޷$i�95��Ě�sK��wAV��&a�=0�o�{�M�7\!�*)TD�6�(�q�nr�n�r�ׯ<���8����^�_k�
�gk��.tw�6P��2��O��/t~�{��S�[O���3�[���ew@��HE��}�F��7z������~�+XN�X���f`>bz�I��5˼�\�$e��I�i�z�b�E}7P���4�ҔT�����j|k�C�j}�&�,G���ꅔq<U\_/&*����4pݴ��6�c�F}*�����T� �#&��Z�u��Zunqs[|C
ٍK�Q�H�����5�m��
ǽ��vS!T�^�m�ZJ�۾�T.>���.��?�����C�,���#o�R�'�[�@���/�P2�_��SU����j�ai�;[��&kaZ���R����pk5�9Ϗ�$x.�+m?��O���#޾����6�ի�{�+|���k�W���Ҁ�r�um�>�S�������*6PD�]���p�i��~qUP+ �q��;�{�$��}Wn_�zpk��������y7}\���~��_�}��اtwH�����l��t���^���Ջ#ꬸ���)�N`͠�P�x��5�EЈQ�RFk%��u�_b�9����6L��z���X��^~���p��C���ⷿ�{s�U��g>j��`��p�O?�=}j��km~?D_$�}����\?�;�F�|��x�,f8���"g�����Ԅ�i�i^��+�
���r��;>&�%&y\=�]�pm{��u-�+�P�yʜ���M�Ȥ/{�ڏ�o�~��P8%3+��J�B����bG)#s��8�\v���)���xˋ|���?5���Η>�1(	��5�O?��?�aY�����I����iE�I[��XߢV�0�}h�o�ӽ���X#U" �/���i�-��ke�"�
WU������#��W��'�bC)���QR���(�$L����!>�b`�&ȑӄ[��ؕ���jŔn#c�D	�/���~�ٯ=y��������n�����ҧ_���$4��sϾѷ4��B?�a���{
����an3Z[px�����{���%Ǉ/��J��K��Z�k���bAkC&��^�M	�
�B8͋�N'@��i3/W�Zsx�����F%\�I���+���'�9#%B���d����)���pLލB��Z�l#Y}��	 2��4ٰ�4������k9��J�WA����>���8��-��7�������@�/|�ؽ�i\��h�G�y�����^�N��wf�ߩ�h�����Ui{�Z �Td��^��G��7mܫ��#��f���a�
}������J׆������,*�#� jC|��I��WhRQ�u�K���%d6�f���i���U����\���w��;O�}�c��̻>��/}�ݓ�s����p���7�6A ��_�E �VA�3�y��镯���t�.>Ȍ�6ײ���{ҖI*�r�2� ���s�>m�P���ٔ7��@��xS����]�>�
U�b5�UKIu�����e�i�GǞ�2��qA�x��y+RE`���{ΩW��(/�r?O��r��/Q��H��r��;���/E����=�;��O���`y������SO�vz[m�gAx*ߣ��Է�ջ"� �C2IUXUX��h��d5�㒮��R���Ůq4%+a����{�}�EM`B\���� �����MLPb7MP.>�E-4�4�\�����������������O��,������e���[Z��?��O �^�����>�j~��[o� <xG=]�u��
�>��{���і;m^��T8^�Z5u����54��mmV5�&�'o
�v�k�z#�����3!�U���(q#2��ܵ!o(��p�˔�g��I�.�,̩��2_'N��k����?���?���^�� ��}��F���t~��[��?�ҳ��P��׸x�S}����[h�Ro�N"����P}Z���[*8a�������խ����c_q��
���7�.?IB�,�m��*����>�0��וf�����m���5-˂��Jɨb�1S.Z�W%O��������px�s���/�{�ٷ�-�<�����o�� �g�ԧ���x�|��� rxn�,�����6�<S8�J�U��o"z��o�N�Ts���(��yO
�jz6O���"������
�6C����ܭ-nk�$))aۤ>�i�2"��2%%NB����J�f%>�
����K�ӗ�����qY꧙���F�^|I_��R�L�Uo{���ѷﷄfw�/|�v�j5��@� /����#K]�&�h�Y[M�IRQ6�g"�邈n�-�iOL;UL
ͤH`Ndc���X��J�d�G�*T�`�FB��5���B}�+��De�8-3��#�*�2�~�'�V�J�����<����������O������/�u�4��|��ѷ"�JT�}�8�M����p��~�N��p:ͻZka���:�D�ۙ���������nI�Q�h�k�y^��T91133)"�b��f��@�Y�Z�\r΀���W��X))1	@ں�-�1QQc�
�
�3���9�gN���U��N���,���>+���S�S^��N������¯��'�
�����w?�Y�؏��}�� � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ��1�Ӓ������   %tEXtdate:create 2019-08-11T01:25:28+00:00�d�B   %tEXtdate:modify 2019-07-26T05:04:57+00:00�_�X    IEND�B`�PK
     )u�[d��   �   /   images/a262aa33-74c4-460b-b0ad-c746896f6744.png�PNG

   IHDR   d   d   p�T   gAMA  ���a   	pHYs     ��   %tEXtdate:create 2019-08-11T01:25:28+00:00�d�B   %tEXtdate:modify 2019-07-26T05:04:57+00:00�_�X  �IDATx��{y���u׹���Z�j��ez�����L�b'������2�eH$BaJ�@�dC��`�@��![G6NlϒqO{2��=��RU]{��ۿ�����1�'��n�u�{�[�=�s~�w��ʥ��1d���1@�lL �1d���1@�lL �1d���1@�lL �1d���1@�lL �1d���1@�lL �1d���1@�lL �1d���1@�lL �1d���1@�l�c@�a�z��Ti�R��)�|�H)����]ǧ0�Vg�¸K�F�Z���=:0��y��8L^a�&����4�"ϨH32ʐv4������>Y��6����=�n� ��w�H��)�~�����t�g��!�<T~V�Yz`�����j����ר�����Z�:@N�NF�ޢ���,S�ޠ��NY<�Zk��J��� m
& ̡T�nW���]����{}*f��>s���m�ݽ㯐[����u��)h~�����>�����R����h_�М�NݴC͠���ޘ�g>�?���g�~��P�R8葉ڤ+�T�O�8�,�`�UZ�	!�n�6�a���y6O"ǭVk��D o�D9~G��[�m���^�u�'^"�[^���O�N����+ DF�u
��v�����/M2�P���&���8\��
\��w�z��V�K3�K3���h㇟|������~ݟ����W���f�ȉCD�M"�!Y֕�.���n�Sf�	ch��G�&�q�H5���*o/��%�ݼIj��KI�Z����.J[�(�\ׇGk2�j�4���X:
A�tԿ�M?�Yg����K_����pkC通K�23�*0o�g3�$����0�v�g~�/+�W7��|��ּ�,un_����� I;���\��u��_},�~�n@"��-ob+b�v��X�I��f�L]�Һ^��U�8�E'?vV�x�C�k�;���M�}$�DLi�S����mQ�Ņ�:��(_Ug�����F�����	��ġ`VcrDqf*��q
4SU�NLm&U^�������G��i�8�3�.�۩.tؙ9|fp�[�D����W)�lSg}�����ѡ��0���%�]���pa�[���>PD���~󧢵�� �v���ԡ�����?�j�UZ��ε��@��_
��e���,�=McB�'�pt�&���.���
{^�K�zst���t��I��#���\N������r���4a�8&:��i�M����fS޻�0�*N�� ��%
V^��'B�%���w�1�@��Yuh$L�wQ&�0�3��	B8f��e�wA���Hi��%�?�p-,$|M^�0$ln���ÃN��'���S���;u���}���~g�| ��eP�>Gӧ>�����)3���I�+Q$d���򼴍�*ձ�aѣ�x�M�"D�ܤ,=E��Cdẝ��HKb�=~���kur��0!�-�)���!��D��)�px0D!�`����!��YҞ+sU9��x�T�J�,�OR@do6v�"�J��:������gB�K���E�����Ԡ?±��� ����s�Kh���+��7^mn����&]
wV�:{���i��u�Z�|�I��'��&��=�{��֠}m�r�<�r � ��c%ED��*�	���8k�0�Z��5�׃S�w����i@�g�ׅ�âz��w[�D'��I�Ar<��a�L*�އ\M����G�+�+��߰s[�����
��T�l1�z��=��.� �v+r�v��[�D�KO��c�	�K�N����[_|���S\�m#$ł��y��s��~)�oR�"�qm�ߵU�/�ԃpw��
"��U��2��Nڦ�<���w]B�^�X�U�F�ozZ�3d��(w�m����&�ҳɂ�d^J��)$��D� ]��X0�*\KIy,`Z�S�oا\G�څ��k�ԫ����G(4ED�+�i8���\r;Y_�Fa�bn���V�`���܉'�n��z �}G����#7��{�B���/ga�`:��v!{�%Z�A�q�P�w���~CYT�UM@u�C�D&�����m�O���KY`��Cs5�e@Q�f�\Z�m��-�%*$4�H`ٟ�i2WD�L]VCq�)�~�dQE�:�)IX˵喝
��O=E>U�)��:[[��Bβ�saȜF3�`H)E1��>>CN�?оs������=��;k�.�$�ҩ��x�~���p��_Α7�p�&q�@NTNu����	yф���ά�K���	]�WQ�6���p^S7����N�z��7e�WY��G�95�F��+�ÁBሚ�t�D�,UX�/��p $o�T(M{5�ր�2�gBrNa��r����
�7_׃s̟z���S��\!3X#߳�7��0��p�3��<��D4��Y���b4~�:��˝�7^�H,P��J�ܰ�K핛tv�y��'�w���y�����a2UNQ��8���/#z��!X�4Ee�w�.���9��� �ޙш���.U�5rI?��H�>��!���~�
S%6Y!
F��[ͪJ�亢�"PNтĚ�Ҿ��\�*Ȫ"�윬c�*#��%j��}���y�����﵌r+���Q����5��#w�<� o`Nٰ]M�꿞=��3������i#$�z,�Sm��}ݕ��}�{���ޑ(P���̄ZP^U<P��7�E�)s��p� �Jg�"L��s���8=�8�&Q&	�A@����d��U��Z%p@ e�w�C�� jT���xbn�[惟^��.�ӶxmhI�R�8��X[;��Dn�E~�^��WR# j.�5�RX�_�r�+��]�ʜ-��"���^�t늬դ^��G� x�s�⿸���ԉ?��Q���:�o��� j���g㝫���8��/�(���E�a���r��j�Tܻa/k8S�PY$����I:9s��;��1�M��0RE��<�Rھ��DR�y�2���D�*��$�ETdF�(�8*4�uD)1{6G�����@]-��=F���r��q����0��؜(y�s����@onm/;1�y�&�'����YH��.�KT]xP���SY2�A9qE���	r��������������έ����{>�����@S��/�c��eu��ʘ���	9%�Qڪ��x�"�4a�$ۡN�o��t���"��Z�m�O�ȉ�/SmΞ���%���b[�Ap�����29?gi�IH+�� p"��� xH_�\U�#�8 �=���� �Ʈ��Π�P|9�G�ex����)ݥT�$��5����)L��H��=�c-9Q��3�C���"��BS��4�=w9Z~j;�~����i�ě�}Ű"a��$�ڝ{<��X�1x;"g U.�*Y-���$�0��=��FG*��wi�f���zK�l^���~M��!t`����E�ޗ��5@���R�3�7(T�rl��<��T��;D5�PD��ѹ���d����\�p�!ё�I�#&��Hn=�Afa������[�M�����ox(�}��jߑ5*8�ҷ��D]�kduƵX���E��e��g���s5��w: +�KaS��q��0Y*rc�dZR��+J�*�G�Zc���"4A30��7���ޯ�Q�/�޸D���xs��D�p���.a����6�9%�3ա��XYn�"L[�˭"� �� 1��MR��(a�F��Pcs�6���w�UD#�ƴ�k�:&g�ɻ��P����]^[U��գ�W�s�%���@X���f�S�?��:	���.�B�r8�魐��57�ڛ'�G�͢�k�$�\.�Ӳ3�������|�R�|�|�܁�ڴ���P-���ץ�+Qhlo�)�^��˹!;�S��1C'�aT����Uz+�t�$½�;j�9�d(t��x����m�0H�Հ�"�Yi��BT������5���8R��/6�̽L�FKn�M_r;4��<�\�؊K�E~�%ut���ص;�2��e�@4�����*kY4S���X/���9������
�Y
p=���8�8,Xp��ͽʶ,�{F�>Q�H�Q�Ĩ�SCsnF���g���T���胁őX���}d�$PJR�_Ξ)�
���֠�hGh[���j����'M1��'�>�Hd�D5��8R��,
k"�Y!���C��\Ŕ�AqY�(7��=�b�H�Kr6���e�Nو+_2Kc�����]9ڪ�£���a�Y)@+[3N���?�u@Y�I��2�a^I
��a�|&R��e/Ki�Y����������<}8���$i��{{*2m��"��ZjF�R9\ c�YZ���V�#�j)y�*j�Pj�T))6�����Q�Ƥq��(؟���Z�K�כ�ό��bЃ�l%"w6�s9j�k^\	�m��J� ą�|�(�MҜ[_$9��.e�h5e��ؾ�eJ�F�M0>ߵ�����C���W��4n�&8A�{�^�U,|^x[]��~{�/ۓ��S���r�*��VM:�Ibh*,J2�{`PY��-s�&BU�S��!b%f6zx�"(���u��_NM��ϯ�]	p���[ِ�������C(A��ʚ�&V�%n��Ҳ��m��XZ)�77�lH>�~X���w>�ⴇ�P8Y��e�z��>�!,�S�}%�[��˕�P$+!g�0��Qd�F��-¬��X5�@�iPE�vٟa�T�r7����hޅme���-�a�����Ɣ��;GМ��`��?��{��~�ɿ��'�������C�r.r��Hf@�޾�ѹ���J�ƲЛ�J8����1��� B.N0���=6ۈ3ei��0����E+<÷�V�sI���ϋ{=)�[Q�����#�Ap$�r��q�a(�`�FQО�Y��jî1��X�~�ʍ����C��V!��e���z�3�r�[)W�`�'��?�%��_x���gg�~�Gk�7l>�UH��E�ǡ.J!�dv��:�Ք&�6N���&�1�Ri3צ��=#*�!>�
�mI��P�{�0$j����쵲�ABf�Y֒#����j�����K+GDA�iy_dv�Q��M��T�b���xm.��P�vű|����g�e�X:�JP�W�})B����qQ���H��=���t{��?;�U2�1�	���`���'�~?l.���!Q�w+gD��w��<F��8� ��#$�I�G^�Aa)�un��-O!
c�	����ԋ
�	i(6;��R��	�����|#M�RJd�sRa��
VO^'ANL��Y�k���PY��6��Z��<mMf7�4�t&{,E)�*v�t$F[��1!,�Y�y�s������}2;7YW�����c�q�u�x��T_,.y�}?}�y��,�Ӱc���Z��团�`����)&��|,Q�%�3�Z�T���OD�R����M�όy����|DJ�s�<���O(]��Yx�L�|��X�ǀ�ANY�ؘ 2��H0/n]��z�̍�s�B$+D���"Ys3�T�
Z9?�`NY�h$�(ͲQj�cIQe�_�)��T�~.�t�̳�z�U:�����!�����(��+/�����_s���n�E}��P�{o�����\P���r���J*@S)GG����Ae!ȋ�G\^���P4l�ݞO��+�;�,�}!<��F�R�L���=T`��v������[C�����8/QV�I��@�[�%���-s"� d����uH2��<�P1��:h��gI>�b��I�ѯ�Ch5�������7���st�]��\�v�~7-_x�K��c����YtH��O�-��:�F�"iK�\Ŀ�׏���4�ϐ�x��
�d���Y���Oi+���V���!���h�w�e
 Ң)�;�YِR;@nom��@O���#&���V��UBq���ͯE�.E��4�΂+�5YO�{�F��`d�mp_>��A�Q/���t���h�(��;�_�Ï�|���|����k����W�n�u�1��H꿡������H1��;�^�[��dQ!G��Ȇ2�@qN��A!)�k�ҶVE�V��u2��f�u�k$xn��(0p��]6�F�DSFF!^���+
��l��?W�yn��\Ԡ)v(�6�r�u$��k�
PEO!���$c��'�,]
�Q=�st�t�\���ׇ^�������yo����G����!�v@fg��k/����?���������S�ҡbЅ��e�~i+e%BVG��b�f�n��Cb,�N�w���Ƚ �T�k\�K��'���V��h���]�B�� ^�>]�����lM+�wJ�2u������5)Ly�2�MR�UI5�}��L��k1����k�	oN9Vy�߇�#Y1a;T�&�.����í�~��c������c��i���?0��e|�)�u�T���[itď��FC��'�Oūx��i�\�s����3Μ�-���'���*��jו�6$���-��4��"k����z��J�Z��sը�Pvo]B5��\Q�{߳5�[%g��ٽ)8�eC��0�,~F�_�J��@t�4U�*(�R��#��>�M-�hQ�3�܀�t�m�e�l�a=^s��������~�wx�̇�w�������K��|�vV.��}�?���?b��;����"�e��=�f/.��kT_���En��u:��!j֏H����V��|W;^�K���MD���*��4���AUy���Ss)�f������|��#;���.�u ɎHw���.!��#К��BZG�����8�%��N5O�zGSY�u'�}����O\B� ��Ȯ�H�N���a�'.j�.Ҝ�g)�#p+Ti-Qe��E����a{c��n.�������ճF��w6�S'�������:���H�}R�sn)���>���z�&�3�Uϣ�?M3�����Go�V�3����W_s+��&��N/�G�+���Q���Yz���k۝f�f�����@{��㙄�"����Ju��9�r�i�v������������X��� �:��LT��N{�/)<L����l߭;�f�y�5����ߗ{�<r����.��y/��^"�@�ZI=�F?s �<8^0��U�s���t�s;���H�}oJ��y�V_y�q�����d�����~�v>��n�%G GS+]A1��4��x*�������D�ۊW�=W��k�>��/]�򯷛G���	��P�_'�*�.kqgv{��RoQ7�d�*qR
}EQ��0�і���|�>9Bൕ�e2�-�i��,�bؕ=>'K�w6h8�KG��� `<PRvP<�)���y���?�ɠw��G%�:��=SSt�0Eu�婙�H�Z��S�z��M�yם��?[�N����s�<E5�X�����w3���}ȁG�CwΝ�J����is��*4������V��6}���ȼ���T+�����ڌ)	w�9�_����W~��W.�C��%ZlP-h������}/^�L?N/|�b`|P��֚l�nܜ��U�y�ؗ��ڇ2�[��}�[����<t9`@K���w:�W_���BՇ�{典H�o�4�f��2-��_���[�p�C��
��9.'u!\1���tz�5|�|��>t���W�9��D<����Auߙ'�~�s�"�?�7i��D�����G~��_{)�]D�D��.
ɵΦ��j[Mz��ץg�͆t����q����r�N<�m�W.~���CTi�݋�%�W�ƉluKu�P����FS��5����� ~i�~��wt�?�}�w�����O��O���wf��c�W�c6&��٘ 2fcȘ�	 c6&��٘ 2fcȘ�	 c6&��٘ 2fcȘ�	 c6&��٘ 2fcȘ�	 c6&��٘ 2fcȘ�	 c6&��٘ 2fcȘ�	 c6&��٘ 2fcȘ�	 c6&��٘ 2f�D�{��w��    IEND�B`�PK
     )u�[�c��f  �f  /   images/c88b2895-5e8b-4a57-9f9a-b80dd50058b1.png�PNG

   IHDR  �  �   ��ߊ  TiCCPICC Profile  x�c``RI,(�aa``��+)
rwR���R`����b
����>@%0|����/��:%5�I�^��b��Ջ�D������d ��S��JS�l����):
Ȟb�C�@�$�XMH�3�}�VH�H�����IBOGbC�n��ₜ�J� c���Ԋ�_PY���Q���Tϼd=#CsP�CT�%���X�}�����ߍ�������k'BLÂ�A�����΂ĢD�33��10|Z����� |�'�8��,������z����j��N��������.j���p  !e�2���   	pHYs  %  %IR$�   xeXIfII*            (           J       R   i�    Z       %     %      �    o  �           a���  �zTXtRaw profile type icc  x��S[n�0��)z^�8~$R��b;^eW�J�ё"�@`H�n-|DI�D��@ȴ�v=L�"�	�s,`�ۮ��z����"H����pz����3�ͬ,9&�h'�tN9#���(���d>CQ�h�|q�k��R�R����mOi�q�6�Z�ܶ=���C�>hrK$>���U`�͚t3�s;����%�S�T�c��\���~�y§b�_"%�G"a=}J�H����|)�Ni����2��yl�c���r�E��|�7$��8��s���.PJ����
��wq�8��P'��j����[ܞ�c2����g�+��|����RM�=�c2gҥl��ϞauTh���҈�\�z���줡㜥   %tEXtdate:create 2020-01-31T21:31:09+00:00��y{   %tEXtdate:modify 2020-01-31T21:31:00+00:00	�   tEXtexif:ExifOffset 90Y�ޛ   tEXtexif:PixelXDimension 1391c�   tEXtexif:PixelYDimension 800�요   (tEXticc:copyright Copyright Apple Inc., 2017���   tEXticc:description Display P3�y��  a�IDATx���|SU���M�M��ޣ {��Dq�����~�V*�~���(���(�"{�Q6-�-�M�{�'I�M������K��{onn���cU{�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!@��-[a츱�aC�5?�q8�^ݺ"���0�
�"���l�a���>C��p���Oo��vn����"��mE�9F�1\���?ۛ�����(:���c�X���_wlP(�ʔ{���=��|+��#}�Y��mo�w��k��]�o�������?�O�0�?���'�Q���W?s��3��"Sڶo�dՊ�}�I���i�f����gf^�t8Z������^d�g`���>�n�q�0K���k|=Ϗ���5�1��}���I0�p]�y��U��'3r��~'_{���G���ߢ��h������1o��v�#�����޵{�I��z�}Պ�ged��x0'""��!;;�߁�������t8�ADDDՎ��4���N����E�l4"""��L�����QQ���ԿTP�UK���	���sn������BDDDՓ}����{�������H/�=��|!'""�c�4a��sh׮ݔ�#F���u�}�?_+.q��p8PPP��o�O���m+�p���DDDG�}ǎ툯0;+k����C���PA܉��\��+z��I#<r䑓�\y���O5�Q�?�^D��R]�]R<�5k����q֦=11Q�s�*Yǖ�Ull,���0�C�Y6'"�`V|֠g�HKKS�o����T���Ύr���������GXd$���(T�:����=3+Y*��D�~2+3K��H�h#"���sx���_����`:͈�����O��;r��"""
f����6.��p�)�ggg��oDDD�����R�7Mgx�'�����"""
n�Cii����p:M{�'��]��QP3��SSѼE�8���,�3�:gOݟ�F��:�������y�
�DDD���";+;ơzI2�kff&���(��j����H�4�L��at""�`&��:���K@/3�^�a�Љ����nC����E��J膻��0���(���*w�^���(@VV���(���*����:��D^^>���(����p�Yo`� ��;w@/;�����FDDD�Mr�0��mPP�ϵЉ����iB��'ԭiՆ.������Q�V�%""�Qt/w���^J�&�΀NDD����m6È𶁴�{+�Qp�/^�T���t""��g߾m�*���6�Q𲧤�H������]��1�'���i��*w""��g����m*`��r���/��Ä�m�����NDD���3��G@g�;Q�S%�Æ����˝��(��3�����G����ΐNDD�Lس23��i�I��S��)U�ge���'{�3{NN�
����%�;Ճ������zdDD�i��K�DDDA�T=&&Ff��Н*�;Y�NDD�L{xD�t�S�:M�~Q��l6;|T�;�&L�Љ����=L��*w�Su"""
^v�a�ax�&�܉�����0�QN	�U�DDDA�T�\J�׉e���U�DDD��.K�|tV�3�|�i�̽t�U�DDDA��%���F��8tV��rK��U�DDDǀ�����t�K���˝��(���K�z���X���(��E�{	��7���t�,��ʝ��(�ٝO	�:��:űʝ��(hI����4�r��YB'""
fv��a�iz	�n?7�)���(�ٝ�sm��NDD��r���SQ�n��^�n��GDD�쐕�L��T07Љ����)U�J8|�r�Nq�DDDA�n+/�K�g@����<����@=?""�F��0;�*��乸ҵ033ii��k�.$'�@jj*>�����9	�QQ��S�ѨQC4k��6���\���1%>�|��%rpq��+�*3��?V�Y�?���Eb��-طo/<���<W�C=��,|��\`�!6&u��C�V�ЫWO0 }��A�&�f�1�Qȑ��i[�I@���p�{�W�܌���X�z5���;�:��V�ޯJ��(��Q�w�{�>)ͧ�Ė���/s0i�$t8�#�=�\|���ܹ��v��D$<�����pU���Ʉi7`��r��s�C��\�U�^�x1�����n�n٬��E�ۆ�)����`�E���Oq��W���GR���yv"��\�g.~��w|��g���;п_?�i`7нN��¹�}�\�-[�b����Gcǎ�p�W�����=轢������i�O��P\p���������O���u����拓�'�S��o�T!����>���2>�͘����3������_��p���T�Y���tf������ذq#��nԉ�cP'��'������ix뭷�|�2]�Y�^�z���'��2���V�{!�Pz^�0���*RS�µ��Gݷg��g'a��Mw���������{���#R�۟���#G���x䑇Ѡ~}u"
Zy���7o&��f͚���8��yHo���;�1��&��ޔ�y~&M�\�f��`�
���hܸZ�h�:�E˖z8Z�*UGGG#7'�z8ۆ�n�:lݲU�TU�[�Z�QV�a����HOKǨQ#� 1�A������K�,��߁�����Qi�tn��lC�C�����g�><����!??�oF׵kԸ1����3���&M��v�ڈ�{o���b�ʕ�a�:�~�:w���Gf ?/~�$��'�@LT�:�Ca�^��,���eʐ�0���or�gf��_�G*��`���9Q'>�>n��V=��v�Z�ϖ�|/C:�5i�H?�~n��L�<S>�\��S�5��s���[h׮n��z�~Y�(�2+&K�"��n�f9U��W\�Á�U	x���s���Űa�p�9�v\-�_+Ƴ�L�׭Kg�;��|2��֮�ù�J������ѱc�ؿ?K�DD!Nt�s����!�{Μ_���~�2�M�!����#г[7�_+O���/�	u�b��aX�l)�36�6��ѥK�� "�P�c�i7���*w]-̀^�n�ꫯb�d�z��L����p�Wb���hռy�Kƞ��u�@����~�H޶�����{�	�_xK�DD!ɕ�۝�i���q����0��)���_Q����p�����FTI0/N�}�Yg�����ǟ@���(�/3p�@*�y�m�4` ��cP'"
9�����rg��#���,F�9Y�.;ѵ[�G�M�VG%p��,2����/�L񲕁?���?���%]""
I�L�곛�k�Ԛ]B����i_c�jo��L������ރ^=z�R�'�N݃~�os�o�X��3��0s�L�{�DFDT��y�"X�X���x�����X]��:Ne��.��� ״������͞�}���[8�2{�u@|�ٸ��K�ɲ'8�w�{���O��������m=�c���xbP�p�ٟrss�����f��u&"B=�ߞ��y�v����y���Cn^���OV}���a+���N�[�8r��!�1�(ǲ��V�Nq�|����EFxȹʵ)p�>[u�rm��ץ���u}]�����OC��:����9�?���"��\}��ˌ���^��Пc�{�hU��)}>޶�R�5RT�y�s�C~J�@~�V�,�[9C�����57"��_@��U�?ϙ��+V�ۭ%cͯ��zԍ�?�7�/&:�^v	�M��C�0���-lطo�-_���Y"v���X�vV�Y��6`��]f��S�P�,�B�Z�ШQ#�n��:u�q�uD�����JZF233��]ۺ		:�*�>��)�f���X�x֩��s�N�I�##"�{hѲ:v�^�{����k�}^ŏ�r�*,Z�k�5۵k���t@����36o��{�@��]о];Ԋ�����u�8��W�3K��t�	�H��r��!���Q�X������u���lչ5m��}ջW/���u�9��a��5X�p�>Ύ;�q$C�����M�4E��ѭ[7$%��k U��{2��3-=[�l�K!�9n۶�))�����C��(�OL�3A��E�ΝѦMk�V���~�:��.�����MIJ�)���+T���6mB�>y��zK�D��f͛��,�u���㐘X��ZT��gVvv���}<p����_�X�����)�T��21g�(��t���k�8t�(���S_om�&���O<�R�>}�]}�������֊����m����ޭ{w�P��螛�J|���f̘����[�nEzz�����u^��t ���x�s�98��S�P%���w���x���٧��U8r%���5l�/��2ڵiS���C�o������
+T�g��>އ�";4h����õ�^�A�����8;U��n�����/�l�2���w/�k����(u�p�)����N>�$�R�ؑ^�/���<iR��r]d��_��*Hz����ᇙ��/�x�b��>>_�͎z�����5�\�s�g[O��J��`��F�ܰdrd�$���q�#T�T�9���u�	�$xUU��\�M���5�'���X�d����Hp�uT�.�6P�]O�ё"��*�W6�{�U�~1#G�ҁ�0��j�L�#�<Rbd�<������ս>Uw�MNNF���zoR����Z�.�1�sp��#�}{���� ���'��o��H׌2*��ґ��,X6�����?��v��#����.�С�)��^��C�`�l�R������;�ޱ�A.ǭ���*�4h�=z�K1�tP���>��U�ɫ3U[����{����z�g����t��.��c�JXd:ܛo�Y�ʮ'� ��%�ϕ�X��$�9[�
y���N��r��z�8�ޭ2�|��~��^v)U�gR�ve�]�b���ٳ����:���q�*w{�6|���0�Ǚ�Zɇ�J�͎��T%���_��u���<�+�ȿ����_�sGvv�_�+�lʾ��5�����y��ǟxݺv-���I�����B��Z�'_�.w�ځi_}�9?��ŗ\��{I����'g�k�|���z9ϕ+W�i���-�����nՏg�T���p�������KGb�*����?�{���K���Uk���̾R�����'[[��>'�dIAa����G��o֙)��L��M�����Z[j�֬^�u��T&��ge�ԯ���(g�pKU0߽[� �=�%~�q�I�������5�گ�GZ����[=�m؀�^{��9N;{$�6%������/�E]�r�Z����5�m��֩��,ǘz� ^U��7����}(���\�;=���}lٲ�����]J������7'��^��=�ܯ��5sm�?5o���ά���:v���)푆V*4u��p����N����|���f�?c�u�!�_L�[�n����|��"�>� /���]ŏ��VJx�n�\��cǢo�^��r&�9�UeXe�sU�-//��<{s][ɠIFsŊ�駟�裏�_����2��-�S�-��⟩��]x��gT@��&��̊ٵ�̮Z��?���H,���>��I����6��x���r�#����D�Х�2���>���:wB��m�Ӗ���[*J>�9*Q{z���믿�^�)��2�J(2���ч�R�J�H<�!C�v'T�%���'�x����d�k����~����@?���B����3�{5j��4dee��2?E�q80��oUf-�Ox�<�$�*�9
o��ffT�|ſ���Gzo�3�up��8���J�/�_R���>������O���$}�+S%57�F���Ƕ-��f�x��r��0��iذ~=�}�\tᅺ�_�SXO���/�£�<Zl�)��m[6]��������۶n�NjA@�����:lM.��t�t�2[�зO�׉�:�\jf���C����໻����m���WJ�Y��d��bX�w��_�h!��^�����_���*ڋ�	Z�1�w����a�B^���t|߁�'U
�4q�Q��-,���1a�J�=U�9�����NJ��= �r]���1��W0��	�ζʼ�������yx�����K/�Nco��^;i(��?��@���u�ȑ#�h�#!����F����9�[f��zH��������|���ū��s��z�
���zg㪫�
�gYڌ�3K�b�c���+�������Ǚ?⥗�cܸ�������eR:����ǝ�Tk��g��Ѝ�bz͹xť��`Ϟ�^����B�.]t5o(]!OR4��Y:t6o� ��ê ^�~��8ӻw4k�u���UT�h��]z���˖��]	��=gö����Ï�k{�E��T�ק�~��%���#"Ѵi3�B]Su���7';�R��Ҕ�n���VS�JЎ||�ɧ8���|�
_/�]	hLl��h��m�"11QG����uo�;v�;�Yg|�T�H��E_�.�W����=u�4LU%9W{y���D�=M�4Vץ�>o�$��RSS�a�l޴I��[_W�2L�:_r�
��0�L0w]���u�4G����u��n2�Jz��]�V]�dx_�X����(��N8�_�������ȑ��v� ���N��B��I��K�.�3�����Qڵ7oެ۶�'|��C�.Fq6=���=�;�^�I�$��t�2L�<����\ރ|O۴i�{�K�HG�C��r�򹦧�y9w��LӁ��}s���c��A>�G���}��/��\=�7mܨ�[�d��%�ף�t�S�֭[6+��)s���2>�����ak2�H!�ک��H 5��_�|9�?5��`�Db���T%�W^y��#פtu���ԗW��M�:����k�Nx�;�oÓO<�F�h�8Ce�Ru tu�+
�R��ۯ/���J�v�ih�����̈;)q�P�9����oM�R�1�f�Ϟ{n֫���]7�
�u0��3p�:N�޽Ѥq#=��s9���6�k\�����}{���#Ìf��:��^��"�>R�s�v.
�a*A�ޣ7�P���[�j�;W���W�dΤcۤI�����e�	�34t�x̘�طgRS���v":�N9�\}�U�qӦMu	�s]dH�֭��ݷ�����W`���"C�O���}zW����3�ǘ����yp'��o�駝����,���!�1�S��߅�����Y�,2K�s�{]VN����y"����}��ΕΠի� g�u&.��b=�q�ƺ7���zA~>RTfm��%�����H�Qِ�o�}�]�pB=����m곸��{p�-7���]���;u������gj��Q#1��u?�Lɐİ��?��kf@�R�+���D6Х�P������*p_Ub'�|*~�a�q�@Ĩ���'9��x��W�������6g�l��X��mX�z%�W	�۪�Ѩa�J't�P�\��T%���;q뭷��JPQ�L�p))�҅<������>V��t�Q%�����[���x��Gq�E��P��8R"�ݳ�w�'��?��*SeyUR��N�m\�а�8T`�*�G��"�*�ȃ�Եi�Jp�+c�\��-[��u-q�
�R��
�e��B�u��l�kޢ�=4LW97�_��K�jת���ҹ���N�ñ��?��IUb���{�͚4���^֬߀ѣ�ww����'�n��s�mh�2c��:��&������Izʿ8�E/�(ٰr�r�S�O|�Mԫ�P�{]�냅�Q������O�Ї���멈s�m�y2��|�q��aʔ)5r�:�����$C�j�9��nE�Bf��Gq��Յ���2����4��>A�I	��zg�'�q��ϬH�Zž�b���u���1}��qc�}˻C<��&g<�[��c�=�i_M��8B�)�|�ɧx���T�V�6j�Q�G��7�Ꜽ���R%����믿�vxz���T��^��K�DwZ�VaoǑ`0d�`]���۱g�.��lܸIWG׫�$.֊�K|ݺ��8����I����[Ǥ$<���X�n}���H&�ƽ8�{��1ͅ-���?U�1c���nƖ�-�c`��d=#�t���a�ĉX��[�թJ��1b�H]����ɞ�V_]O�II��V�	V��3f`�*9ߦ2��Q��J��u�_��T�3�9?o��!�Ho��]Z��~oSKK��|��:��^��X锸��Zzj|j^�9bz.w��멚�)N:rI��+�['P2�HL%&�6�i�ܵ��.2K5�u7p� =L+�]�#z�����J��t5���H{�|�ǨK/��\gW{�C���]����ݯl'��I�ᤷ�*wk�.=��`^ѡ���:^t�:�D�g=6X�z�J�+��;�w�q��ů"ץW������1F�t}��H�[O<�.8�����{��N��T`�>��C�aݺu8EmW���]���-��V�e��O>����+0��g���L{����t�{�+6��hˬ��z(��g֥〥)�|��a�葅����h*�I��K/�K�,յVs�H��c��	�N���Ց]���g��m�vM_d�p/SfVWs~��ŋ�[0�j��숃���V�ǞxLw[�'�([)�l~��ttx�� u��8��tӍ�ڸ��A�L�������mE��ύ7݄s�����9IIpР���O�x���1t�=iK'��֝�RʖL�ۓ�Fj�>x���J\~�e>k,���*�O�4��C("7JG+����S�#S�Ju�Ν�U���|�M�A�n+̋�Ƌ/�Pw}a����$C}��1�����Nt�p�Zb���W^#�j�G�)S�m�U��y�f�?p $k,��Ͱ�۳�&��KG���l[�V��P�i)��~��7�Y��~i�'�T.��SN�|;�����}�}�a���k�������s7�p�n���qM=%�u�]W���:w�&M���`��G'Z�l��.��2:$�~b}��f���A]�&"#�����)�Oj�V�Z�:�y�xm�>C�u�Ǒ���w�5)P����蒤�NS�*	����2��:wŭ�ݪ�D��.���o���f��.�+K��e:��^�\���0��$��a�k׮���B�{��]��Cꚻ:�ѱbJ��M&a.GMkC�_:Qe����B�+�ۄ�y���$\q���L��OI�.��=��?�:�X�b��5hr�9�<����uĀJ�엨J;�u@_�u�SO;�U��� �p��z���L��U-��V�[a���+���ؼE/S|��s��ǣg��*�JB����m�uQ��^�s��Uj+�2�aa�ͼC��z\�ަuk�{޹z� ��ҿ�.�M���[�5h�Hw@�L�kO@�*yw��	�M�n����̬��б�>k��]/�jb�db��[J�6�`�=D���3�:�[�
h��Kz��w�y�c�UU����0�!�^}UB)=g+P"UF�a��^����r�#��.N����72C��- �>=z�@�J���u��$��ye�лO�J��/���KH��uY�C:�z��(���3o�<����^v��F���,u��x�	i�8p &�5�G��ۇ*�"�Kf�c����(�;YAN'���*s��"1tL�v���u9�����M�>f��ܵL�*�W�L�b���:2ɔ���B�F�4i}�7\�c,XY�K�}9���B:]�t��{��_�׶BSO��1 �Ԇ���qb�>/A+�g��IV�mV�5�ef�U������U+Cw2S׿V-�m��zQ_v�ك��Vx}�k�nh߾j�Hr7M<����J&ϑ9�s�n��^r�ש�������"B���VMcNgH��Ւ����yU��n��sTt�ϭ$G*������٧�`)Î��z�Y���j��ڷw���n٪�l.=����� �+KWT��{�ԓ�4k��e�����H:�1u"ݮ]�J��}]t3���A�?�l��%ǩlgTڶ�ː@���;�`0���I����K[7o�|�y�w53+���m�Fe
7O�d�$3lU�.�Ռot4�_˫r����$ш�Yb1��4W�Ȕ���ɬ�i�u}TsV��]R�����<�b�0��;v�eJ��(qq�t'�ʒ�k�')=���y?�u*�픡��&ޛD\%t9Ve�U��쨌M�7##����=\��[Uj�_��d`�e|v�ڭgᓀ~dLDFE�q��Nz%�*ڼ-��b��/�$t���g���3�I�!���*s�I[]%�Ƃ��͝��Y��4C��I�oU�	��!+�Ig$�6:�t����W+N=j��IЊ�=�Z��k\�V2TU-Zer�t��*S)&	�nݢ�}�H&j��=���_�HaS��L�*�Y��?x�S�W�8��A�@L:TD������YCg&~U���JJ2��M�����۷O�U�w��`���4�eɼ޲�CU/BӴi]��(�8��;��[��.�?G��X�(U:�N�H���Q��H�������܇�}޷G��YO�����Ǐ�믿T�o��ѽ��z�����d�1�F��(8I	�^4o�L��]KJ����MWz]=��i�suj);�7�����/�yJ�99e�2�:Oα2w�T�JG��&�;F5J�$�v42 R"=��M��R�&��x#�k2��q6e�&5��؏�d����j�k�#�\m�5�m�Q�ƈ�]���:�i{�w��`&��[�M�*>
U��1���Idsr+7,�nS�+�����]M��W���e<���X�����z�Uѩ��jH	���n����dLm�zu�o���.;�Ɂ������O���V��G��*@Ib���C���l5s��J.�J�*��<�f"W]HG���e��@u�*��d�;Y����r{��jh@o�X퓒�F�3^�kv$Y6P��7o�3e5o��u�`>?��>�P`��+\��U���Q�*��SNUC�1G9��qk%�Nӽ�0���pk���a��򎥚�gϞ�V�;���˗/׳N�`��ʒ�F^}�5|��7�бz��޽{��%�KOfo3_IU��`)�hf��0HR��g=9�!c��5>�'
��L���C�v�\�3G�f3u���@T1�Yn���5��^*�K`?�a=fu��eض-�:f��#%g�/%EO��c�6����l��ZĐ�3z��K/����)�N�p"	��(�H�`)�W5�s����OT͝Oǎs��
M�?��$&�?f��:U0��8ӟznC�u:N�n[`��(�mHNކ�9�]�]��7�B<�*=Ʒmݬ���ڷo�zi����A�p~PzȘ*�gdT}�_��Z+�و���Ы��`^+�{'O�0J�\h�8��TT�Mu�H�ʽRU}'�zY����?���_�e��]	؇���%����t򓕮�ԫ[O�Ѷ��(��Ν;u�۪v�59���v��1̍f63�٤������Y����mT�:1������]޵Ls������U���v���_�d�R8�rF[�nÌ߫�J�̭>RS�v*���� Q�������*K:ffe!.6�J����]�N�L*Svq9������m�2��Uږ����۷��~�]���R����ft���;�-^��k���Æ�;vbʔ/зO�c6C��gb����|�z���#q֠Az-i�O�^�zhּ6m�^�e�Mz�}\_s-������6��u2;�$x�����BNN�I�d�����K.�Z�%yd^�#��n�Ն^3'��%k�r�U)}���^��u��]vN9i�Q�b��yr2>��s���d6�����mZ���O�܇gq����1��_,�"��u�֣e��
[�n�ƍ��mXY�֭u��(ڨ�^�nv�*��|#d	S�z������H���.���R� 'AIa�������������t�m6\~�e��/�q�:��ٰ=y^z�%t萄���G�)�L@1y��X��?�7��s���0{;�������`�1�Х��Qe
N+LtE�i�쟱{��>���٫�^~��ߊ �y���T@�a񬁕+WaŊ�8픓z\��������s�~��*cQ6@�&MФqc�h���:�����N~3u�	[yU�5��]�}�Νqɥ�`��qz&'+�&M������ȣ�e�i�l���{((��L&�hּ��'A��9���[q۱}�f�*���]wމvm����ٻ3�NG>���ckšO�����}'R �=$�����s����>uON�2����.\�_���Ԕ�أ�d/:��]�>�p�'�se6s����巽BL��:/l�
�W]}��6�[��e����+HHH��s"�ë얔m�*�?�̳ػ�[�z"��.��{�*w�R��ۯ�;��f����0u�T64`S�����|K/���ŤI��úw>ё����3�w��S8�����^ݗ�^���k ��r�ÙY���U0���;��2�UI=�S]�h�����z�I�YN�l2����~�m�a�S��p���؟��}N_��o����W�|�^�/��,^���dNt��7�|�.e�:ݎ^��?�|UZ����&m�'N���N9�J�/9�e+V���^Cf�� ({+JO�s�=͛5�B
$��ڧo�4�GX�1�=9/�8mޜ����W|e�Q���o�nW;g�uV��i��ЭÏ4�y�d����Ə:sJ"\݀7� ��*O��+/��6]���O�^<p?ڵi��	D ����3Ĩ��x��`����E�.]�>�Yg���y�υU_��[6���c�L%rmZ�:���j߇^��*�[�V�hѪ.��|]�
���O��UW_�y��!+Ӻs܌�CR�x��'sd�Lxz��^�cǎՙ~o��N���5ADd�^��j1���<�Kܒ%�ωe@p�v�����ª���n�{�X6d��a�oa��ŸM��SZ������6�I]6mقw�yWW��L���NJ�W_}���
�۞eY
��oT���*�;�����J4�0t�0�ya:�kW�DN��c�.<��p|�ŗ��l�$,,�^{-�w��`NU��s��_���V�z~~�|��G������n|���ҫ�ɧ��?{�j�v��|��hP�~���ccbi�?��}���3rM����t�SB7ٖQ��XRU7��0l�CؽSz�Z}A}����O=���'�����y��'�u�V��c^r9��,lܸ�~����5V�Ҭ����X�W<s }����}���~��3>��S��e%��_���}��GqҀ�^�&��Zi..Z�J*���7��/�p��	'���E�������{J��}��WGw��.:s�����q�
�����"G%_��Q����g��Y::{�ٺ�����w����<k�̾t�����z�T��n_���N�e�U�Zn	ݕ蒇L6q�嗫l�	��jއ��Ds~�	���;Z�j�~���G�����84i�1��:�K)\������{�`ٲ�X�d�.�oS9��Y�|��LO��1ϣm����}݄x�Y�իWc��%�J䤏��ٳ�f�\}�5�����!)Ig ��N:mڼ	ӿ��>�[6m.�WYN�l��?��^�`NUi����{���#��]z���eMM����q���~-[�@���}f��`��ǧ�->��l\���8ѵ{<��Cz\zM����j�ɢ֭�z���];q�}`��i�ԩ���9����ߥ�q�1��+�ak�r���6`�ZD����_�uz���F`�~�+odC��v�����٧vĨĠN|��)�H@�ǲT@Vw�����}�߳|�I'�ŗơO�^���ӫWO�5��s�^��[-Į�;0�����T/5+��e<�L#����g��)Y�p!�'o��᫆����`��0���@T��b-*(�y�ر};�y�/C@��z���xRe�'O���w��4j�	ut'���=m�r����زe�*I�.��{�F���SO���WMIg�}Ʃz+U��s�^�ru2���4���as��2q�i������G��T@/�#�蚢*\����$��z��c\r�˗-��Jg�[��d!�Çӽl��J���0���{�y1�Yt��9 7�9C�F���裏b��M�ԥ��k�v��~�=�UxD�c����<��Ư��M�5�SÇ��T����hеR*0H&2?� ���C�v�m�#遽i�z���˯��uהφ������3#��y�&x��q�X���d������u2
���X|�\������{�a���HP����z�Q^���ß�Rsx��e�^�6mZc��Q�q��ɖ��\+o�:W�L�ÿ��[q��w�I�FKdH��a�����ß��E���^)z����I���ʕ[�ҵ�J܆�63���&%ntlɽ�X}wF??J��ߞ�6�I/k�Mi�W��*�+�[^F���mݦ-�����
�\�����G��X����f
�))ػo��Ŧj�
��k����={b�ĉ��������H�|=�ze��W��SO;��s7�W���$��;g�^Fv�8���-2����U�9�s��:�	���K����ݺu�Čp�3���^��:�=��Ӻ���W^����aZ� X�E�ʻ���=22��q�}�����DU�]N_�#�=���{?v�H��A����HNN>f+\)���ˣ�����?��ުґCf�[�j5������G���!O�[OO[y�5W��s��OH�۽kL��:��x������,l.�H�M���O���O9�]w�^�F&�����^!N����5Z��W�������@�S�Z4���q��^��z�Ksp�	�>����*�e���G~y]lt4n��z=c�dοV���7��~?3��C���
�Q1�ر��Tw���6jРR���Ɏ�{��^�Z���bu<��qD��Is�|��F��}\(oi���9nӦ��=Opv�A�Н�����Ti����õ�K�L���m.���lݲUw�������HH�G�vmq�	'b��A�ӻ7��M�[�*Ty_҃]ޓ�������3�`�?ر}������К�fG�
�mU�\f�2dN:i �={+}��^�[�e�v:�zᜰ��Wmʾ���t�ֽ�LWr��I�V�!5r���֭[�kWu���Ǒ��S�Jur��=�d�%�v��!`��ʔ��{�,�w9���� ̋.׿Es�믎Ӷm�A�Hy�:��2r�sz����9?��ʕ+�����ɽe\
Oa���Eb�D����w.NS%r����Vi�٣�
n9% ��e��/=���tb릮yZڡ��/Sjk���W�\i^�fK��|���i�Oزy3���c��B��Zj3dTP||�����K����]],�J���մNG�s��gC�t�8�3t�;v"y{�^&TƖ������Y���HH�ڵ�PO���5k�\y�W]�fw���[�9��&w���ur�v�Y�F�N�e��Y%#=]�Ws�$*�j��^f��ر:w�W��#d����׫�	Z2���$�뮻���V"""W��+�I���>����QQQ~�ŕ��qϊ]�#>@���S�/�r�p��}e�#������-7�d��|b��+}lԵ�N����6m�ڵk�z��}�����lnn���bս.�=˒��ڵC'��v�{�Z�Z�
��s;��S��w�-kO�\�����S�|��/-�%� _��C�:�����Sqݮ

�����~%'�:u�ѨQC4i�T��1�2�S�
Ԭr�"�W݌�*ˣg����ِ\���5���@$��A)J%J2�Qj�����_��%�o��>�]� C��2w�zߒ ��� ��Ë����}�u�Dӓp�:�ʪ���qU{�o�VD�=��������"�LU}��qq�Q��)�/�I���&=ⳳ���ס�}��$�(:yHf˰�O�H/����r�;P�7��aUu<O�Tc��Q�9��k������΀^)f�K)C�\����b?�w,��#��L�im/��;�hݥ��8��|��8ގ)�ňp�z�����<��58��0K���0�~L��6�@;�\{u�yy�PM����Ni��f7����YB'""
f�S\�[y:�Q�ѝ8�)������^����3�-ӯ6�|v�#""
b���������(�ٝN��ֈ���7=S\�[�,HN�Љ������W~	]�9:����T:v���3M�r'"":�����,�Tn�7+�O"""
�K�ݯ8-%tFt""��d��m�::QPR1����DDDAKW��UBg�8""��e��˝Et""��U�:#:QP���U��8t""�`&U�~lU�?"""
F��ΈNDD�̊��3�)݆ι܉���;��~e/w""�����,�NDD�L��YB'""
jXm�m�DDD��"���������r�z�DDD՞S�r�5""����U*�}�k�r'""
ZR���VN�f,'""
fz�5?7eX'""
V�ߋ�0�'��,�U{�˧2�5?�r�܉�����m�r'""
b��U��DDDA��Nq�����(��~W�Q�b�;Q�Ǚ∈�B g�#""
~�C�˧2�+��^��DDDA���2DDD�ʏ�\�L��NDD���ΨNDD�����*w""���*w""�`�ʝ��(p�8""����kb=S+'�܉��B ;�U\m������K�p.w""�����\�DDD���X�U�DDDA��Q��LqDDD!����,DDD�*�˝m�DDDA�ɉe�������CgX'""
R�
T�Q�͉e���B��m�&�܉������6t"""
F�U��Gk��DDD����܉����
t�#""�`���WЉ����Dh�m��(񃈈���aT$��UBw8�HKK�!�p���� �`PS
Q���c�=�l����j���둓��ז�n��0l�C��Wæ�5�������]8
�������p����*�&6���e��-�8\yS~U��^�t1����h2�g�.��6��sDDDt�I��f4��&��� ""��JJ�:�烈���+UB7��͖n:�� ""��Hfsأ��ege�U;6�-3:::�^�n��������{�g��0=""�I&������K���;w$�Өqӻ<�t^^^/�4cTD��u�ƪ�3*8���c:1ϑ��g�#|���g��OF��x���$�����jժ�y�����W�<l��k�ŧ�O����;v����LP�F��]mn�G���E��l6�&m�v��0�æ�`ap�4�����rd��ϫXf��Ta���
�+����ſ�F�_JoWl����l�	�Q�k1׉x����󇢿B�8*�g�J����b{/���}����(:f��Qxn(���.u��{�`[�~���0T�.b�ҥ�{v�
/���G���NC�&M�T�^n7TWr�֬Y����[f�������=��ILl�o�Nɟ�f��MX�<[Q��}y�~����1�\4%�Y�wϮ�����,�{������vW��3K���yxv�c?%�l�Kb�R��\��W���)|q9��,q%��[����ĮK��}���n�a���{��_�]�r)�'�z_/)���N�l�b+��(�-6-�Y�b����J�-��ڨ�9��G�}{ΧԖ����t��pJ�e���%���-:�b�G�J�JM����.rџ�ݠ��:IϹ��\�������0̘�hg|BvIIs�����Saw���ʇ���G4�΅�Ϡ ?W?j"�gY"P������Ӑ@�p��ÐB�l�S�t8W pr�����T$u:�Õ��p?����w���&���\]$�b��$�o�^ܙ���kѾ����m6�����u�]o�ٽ�ً\t�Ÿ��[Bnn�;z��͸�λt"Q���N���on���'�<�������OOL�<O�EyUw�g��&�%�f�L������õ�Y�I�?\���u����hY<u���	S�,�;u):/��s�]6
ӛb�r�����
_��G���R�����̰�^����kc��4�ͦs�6Wy��-5�0�\�����6�]^cs[�e�._�CA��o��0RB�zHٿo��>�S?�� O�l٪UH��7�

���Vtx�is8t��4��J4�m�j��m�w��/�(5�_�O!_ega2�J%J��#��X�]<�g�إ{�i�'6�^�٧�Lexb�Y��Z�;�'���|��������Jl��2y�.�-�܌Ȉ��Zu#WD ��x���\���j�ژ��~̯s~Y߿}���E���[_a��p�2�mW|�ҥ�R��(�P�F�s+��(��/��(]�*��2�M��x�k�9��?ós�t�<�t�B�{��#�?=�Og^�{Tx6�k��F��'�����ܙ��r����w��=��M\�C���x�y0e[��|�}������vU��2��pU"R��Ɂ�
��c8�Զ��r���گ�S������r�Jt�ܹ�ug����e�,���o��� ����W;����"�#

�eF���e���سgZ6o�/S�T婌���o�c��-]:�mҬ�ks�u���'`��u���+AD,Щ���T<�$$$����J��ʬWr[�l���kt@�`.�;���*CS���f�^��?�>��t��6��{�Q0a@�2ڷh�ǞxR�����v��V&����a�?�`��A�>������_<��sػG��R���Jn߱ø���vh�] "
F�d�q�&�ݧw�_|�^�ڵ����������:��m;����x�駱j�
������f͚���/s�~y��6�w�� "
6�d)-��p|n���V���]*�J[�j5�nۊݺ�:ҝ���1f��y�l�i80ԫW��O>��/��Lꐄ�cǂ�(1���N�#:&f�
�y*�G��¦;�-Y��������λ����(�	N����h׾ݘO?�$%'�0���:Y�6�6m�ʔ���#���5*�M^n6����\s"��Q����{���K���@��0�=�Q��o��}�'�?�fM��;�"�`ŀN�.��b\{��6�#""|Wf��Ȫ/���K����^�jӎ.�bي�1b$��މ��\�����g��w�;��>�Y'>�G<"�`ƀN^����۴9�����U��Uv[�n����t@�$������ѣ�d�b�	�JtTTr��-�L�655/;DD�:y����`r�ڴi�Ff�*;ͫ��b�e8���Q���㭉1��o`5���W��k�.���� �n��O?"�`ǀN^}�~.����j���s�yyQ��q8�p�"���"*22��g��oLx��ٰ*�׊��ѭG��Np�����޻o���:`@'��M�ݺ�@TT�&e~^nS�v�U+Wb_J
Z4k�`�i75r����`��y���ϛ�����C��޻Љ��`@'��z�\vŕ��Ď�QQ۳27-���m۶bÆ�A�u��~w��b�vs�ݞݰA��+W,[8��G�Գ;n��jU��S߾}p�ק�<{�Z〭�%�:tK�.����`$����˒�����|�)�ߓ���mxi� "�N�ɧ����
���e�Ͷ��뻗�t`ѢE��ɑ�AՎ.'+��'�h7���]ٮ}����-c��� "���ɧ_�͚�D�:�W���g��^�j;iG߻oZ�h�`�״����p���n7���hܴ�����)_}��K�aԨ "�n�ɧ��.B�=l˚ի����Xt��۱~���	��SRS1z��^Ǜ6�,����\�պ�k0�|���K "��Щ\	uиq�ݪ�%=-�M�-����y��y�5�fϓv�I����v��:uz��/�ʱ���)�����b@�ru��I��9�U�a�Q�c�t`������Flt�1oG�v�7&L���[��#���7o�r�/?��y���ؽsN?�tUW�T.w�8�{�^�򚣠� �j�U+Wa�޽hӪ��x�#Gc��vsy6���s�͜�����O��3O���:c@�r͚5]��@|B����������e���ؾ�֭?f��<�`�E���_{�����/���w'OQuǀN�:��q�7�t:��/]�+++�n٭����v��:��(���y�EtL̎�mڌ�����0 ��Qv;"����_�z����/��?x�`�mLӡ�S���BlL�QoG�����7����`n���7i������3#����`ND!���Ҹi�rӍ��:���l��]y�e���ػwڴnu��MB�Ju\�j߻w,�����P��'�<��AC�1۶m��oL Q�`@'�<��Ø��iG_�J�9y+�Ihݹs'�o�p��������`���n��]�v�g�������q��_3�QHa@'�HǸ�I���Y����J,�v�e˖��AgU�9I0�/(��＋iS�I�?����#�7i����[2���ѳ[Q#��ÀN~��q=��t"۵�߅�2�3,�V3��ѳ��sƣ�4�g���k��΄U����s/�`J��]�v�Z<x߽ "
5���m����n94��S��`5��X�z��KA�U3�g��u6�y�w��˪vUX��]��Ν;��釙Y���� "
E����Cҹ�ٳW��av�� ?�2��x�M7VY@��JO�ر�������n�ڢeˑsf��)�a��_����Q(b@'�=8t(>��+ԩS{UDDxFA~^�	f��Ұt�2�y��*9��~�?|���0M'���e6���Mz��W�r�x���0⹧AD���o���Z�i���M��ѻ�23�Xm�׽*�G����ܹxy����̀uU���s���Mxz�3�5�[��ND!���ֿ�?^Ƥ����/������m�5�Wc_J
Z6o��K0߲u+F��m[7���m�ڷ����{�r���_���?Q(c@�
9����1))�s�n+m6���Hޖ�M�6,�K0����K/��彩�-�����4m�t��?��9���дi\q� "
u�T!��ɨ];			K#""rsrr"�n�jG_�l�vj@��0M|��g���>���U��a��~�ĩ���K/3���1�Y��Q���N2��3q�"22r}dT�����&V������%K�������J������k>^�"2��[���ۻ��*�<��?�����n4$kBGMk׭�bv�r�s'k7��f�v�Y�j^Rlk�Uh3#l[��dE!0�&"��*'8��e7��s�[�<|?3g8����w��9���L����ܶ�3� ���~�>*J���k������%��8m�F�Y�Dz򃴘מ���5k��\���G�|}[Ǎ�� ���T�|~�3y��' ���~�6�f��ҥm�3�t��_`�Kjj���ٳ
����Z:;e}F��������zWxDĎ�~����
� ?_�n� �pB��oK�zJ[`ƞp�m%��e����A�%-�-RRR"���;�jQ��y_v��]v�����	:���cGW@@���1��v:��Ç%.>ABCCK||}�m6k�����V)*:!]6�x�}:��W���Xa��MY+��f�����	�����Z�N��M*{��:�m������gŠ7T;v��J{{���_�|%M�&�w����74HRR��*+�^Q���ᆌ=|��W^����አc@�B�d��Sr?ʭ���0�Ӹ��*����	z_h1���ƍ�$���<��
�?w�?����/�k� W29�$��ϲ.%��*�~���p3J�su^ZZ*�Ϝ��s�ݷW�l�"6�U<͛�Un���o�ަ��RXX(��� �pE�1 ?��DG��M�'����X-���q6[�?^$֧�b4��禥�Dq�$'�H���t�����=>�Ճ���; �.\���x�ጠc@���f�~��������k�X:�=]Mk����-�q];��,)�k�d�	����N'QQQ{�WO�?c��v����+ �;��������L1u�
�k/{�$?w��������&[�n�?�#�}��Z!�!E3�e���hjn�m��  A� ����c�>bޙ�uZ���{ڨ���(��e2c�t���ҝ��'37HW�7ڢ�r�K�Z~:yrʮ���t�3R[^..  A� DDE�,0��_�Sl��~�����(/���EEb�Q����{W���%yM����Iϭv7��Fo׍��;�צ~x�;��Ȋ�� �_6w�,���Hxxx�ȑ#-�W�~�o�����XZ��亠����F6��Jj�:���/�Ӽ���ZdT�;�ߙ�>����%9�� �w:L�"uz\����-��dn�����R[S��o����)ٻ����i��%A����3��^{�g5���*� �C�1`�G����>Ѿ^��Ω����t��_� {��S�Iz}O���]��.�X����s����s�bc7�d��ߕ�P�1���y� ��:eF|��
h	)3��6���8m]��۷K��Y2g�,�8wN��$u_�WK/��i���_�Т7W�|�.�,~H  �"���ks��y��t����ߔNj��%=-]���$c}�=rD<=��]�GFF��=gv�ƍ�N����
 �cP^߲E��#gΜ)�;엺�����򤪲J*����Ԗ�u?o8j��֙�fnX���g�!�>yR  �t��%�n�Nʻ�|\z��t~�)�'��MR�e���i�L�]���훶lq���ɯ�<)  �:�d2ɒ����������ں��tz�~���w'L�X}Ͻ��ݺu���ݻD�d;A��tZ��J�:m��/>q����ā��%�GZܽ s�����j��u�̝@t�'��˧G���;�x�iʦ���X�V����`0J\|\ުU�v,8䊈���� �aC��?��{\Ǝ���?���b}�.�K��`4��W�Ǜ��j����pF�1$��^��:f츎�G������q���>��K:�n[xT��i�ؤ���[� �Cf�Ν��ޮm�r�������T����C�i�+��<�����-�  ����2˖,��/���s�J�ط���w���-���*<!!��]wߕ|������� }G�1���ِ������l�X��m�I=��������3>m�^9��ŕ���*/���  ���cH͙3Gv��-oeeɁ��"_�$�ݑ�]�Qn���z�;f�y��g�9��ӈ9 Aǐ[�x��d2���D����t:&8�UN���|�����`4�1��Eǋ���ʤ��V  C��8UZ*:�QBCB�'LL375�X::��lA:�����'wtp��u��wZ,�z�j1M�$ ��!���86ih��^��������dn�:V: `�:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
�O��Ր���    IEND�B`�PK
     )u�[��EM  M  /   images/d3694a2e-5bba-40c3-8069-8db85c4c9209.png�PNG

   IHDR   d   d   p�T  TiCCPICC Profile  x�c``RI,(�aa``��+)
rwR���R`����b
����>@%0|����/��:%5�I�^��b��Ջ�D������d ��S��JS�l����):
Ȟb�C�@�$�XMH�3�}�VH�H�����IBOGbC�n��ₜ�J� c���Ԋ�_PY���Q���Tϼd=#CsP�CT�%���X�}�����ߍ�������k'BLÂ�A�����΂ĢD�33��10|Z����� |�'�8��,������z����j��N��������.j���p  !e�2���   	pHYs  %  %IR$�   xeXIfII*            (           J       R   i�    Z       %     %      �    o  �           a���  �zTXtRaw profile type icc  x��S[n�0��)z^�8~$R��b;^eW�J�ё"�@`H�n-|DI�D��@ȴ�v=L�"�	�s,`�ۮ��z����"H����pz����3�ͬ,9&�h'�tN9#���(���d>CQ�h�|q�k��R�R����mOi�q�6�Z�ܶ=���C�>hrK$>���U`�͚t3�s;����%�S�T�c��\���~�y§b�_"%�G"a=}J�H����|)�Ni����2��yl�c���r�E��|�7$��8��s���.PJ����
��wq�8��P'��j����[ܞ�c2����g�+��|����RM�=�c2gҥl��ϞauTh���҈�\�z���줡㜥   %tEXtdate:create 2020-01-31T21:31:09+00:00��y{   %tEXtdate:modify 2020-01-31T21:31:00+00:00	�   tEXtexif:ExifOffset 90Y�ޛ   tEXtexif:PixelXDimension 1391c�   tEXtexif:PixelYDimension 800�요   (tEXticc:copyright Copyright Apple Inc., 2017���   tEXticc:description Display P3�y��  cIDATx��]	xLW~��d�(%�J"��}�%(�Z���B��_[y~R�R[u�E[[����J����ҿZ��j��B)��'s��;��Ĉ����>���=��s�s��-�37:�PTB��A%DaP	QTB��A%DaP	QTB��A%DaP	QTB��A%DaP	QTB��AW÷&��z\I���7�)I*�Ev�Z�:d;iJ�3mtRɲ�������V�$IY6��"a[�d��$}/����~�l���99��t.��$u0Z��d�M��(��5D��a�}0�*�
��?���h��dY~�`ȫq+��L��yY���@���[���������ƍ����0��`�Aк�C��"�|<B&�������r����t�PQ:�;w'N�{˧����a)y���3�t>���ʂ
E@fB\yyP� �f�3b�1�(p�3!�<ÃY=��䫄(�d���?0��&1A3vH�JIi�	�YCd��c,�p?��0���g�Ж���lqtws���%b�G��ɒ�2d'jaxR�v�Zl߈s��S�����_C���2Js;�i���8�f�ɒM>�Q.]�����С�x�g/�5J<����зO̚=�g����f6.:6lX�t]������B��5�D��;ѽ[7���s�p�0g�,�n�=_x��(���E��~/���u{���F�m�6�2�h��!����v����;����dX�i5�7�}�����ٿ�2~޳?��#n������1p�@xV�$��u˖�Ѳe��H�zi��|��u��,�Ν'�����ԩ3�/�5PP��7o���,�_���C�޽ѵK���ǚ5k�t�:>�,^|q 4�XȺ����7!&&�+{�_�~��d��ǎ	SԥkW�o؀������A��n��B�p2�7n����Na��>$3��ARLN�G��&����~�� �����QQ��wq�������Тe+xU�ºu_ lQ������͐�լ�K�.����ԙK�.��9����(�QN4|���X�p&M|�����5�OLLDu��x�"�.Y�9o��&�l7ww7�b�rD�c�)��?��޽E��jO����[���a�0�?B��ۿr6n����o�Y�}��E�E�:uh@lAZZ*�i`5]�ر�u�9Ǻ��<s�4�V���ի۽��1�Q�n�:AƢ����D�?O�F�g:b����a� i4puuÑ�#������W��u� ̜�iL8^<H�Ȏ��ʕ+Bui������®�v�u�zS����u>l�ФΝ�P�U�@.��+��������^M�5c�L�L��S��nW",�Y��e��'""#�|���'B�B�FMТœ8���	�R��ӓC��w��t�b�_G�R׿ƛG߭~=L�6U��?���קў��ݻ[��Z���\�rLd0�q�	��o@Ey.D<kI��
2^U��~�zB�!C^65V�E�6m�W���$!-^�j� ��溃��������͂�٤������m׮j׮����{��l"��e����G�fg�AQ�%{ΫbM�6��F�흚6m"�.\@�ƍD���]P��	��g�ΕG���e?h�V��\��ӊ�����ٳq"m���`1i.�[8c:fd��Y����<P��6���׻�2�sq�{dDG2kd'j	h�͛��)2;U�jW��%�=z|j���)�b~b����!JcӁ�L��+$3�i��ߪ[�Fc�8����2�F����~~���dG��?��%\�9���ɡ���3lw[wGDD���Ç�6�V�Z8AQ?��6U_"���YԢq�0��$��_M�i������W[P��@�nns+�F*Z��@'����!����ǤI��`�<a�CI�>��p������<*T�[�Cɩ�1K�,>�>}�/�h�M�vhD�*��89�-�aq�֭�M0m�t�jQt������5k?C��M�ۻ�Mk5���Z�e����ZSVY'�����L���������'����F����g(4�Ŷ��P�^G�>|<(��p������_�R�VUDK</`9rr��WhI�6��E^��9��~��΁�ʧ(��K�c��K�^���}Ѭis<���b�s���J�efp �e
���,���5��<�5o۶oD��h���%.�sab��F��%a�ȑ4I܍��u�Ȗ-�!00�==̤?�9@���������A��"���K�T����J��2
�������r�̋h���C�Шn+���\�t	�i~`�'t�dA�����Ӄ|�'���GEDCQ��z�5{zP�gA`�@��?�h����\�h*��5���]�r^^^pbb(��1��[ޒbo�ػ^8�s4�叽|�4�@����4}�#0(h�my
?A�#����Mg�<��7��?�il���_ �2Eto�����"����j�37-N^��4g��)�8����&��'�*JBCLQ�JH�C���=d��,���}X5D�2`�����0��g窆(&Q#,���!�.o���e�TF��[���9ʲIQ�[�<l�M�V��|/="D�xOR���vG�_G�3˚��7��aj�gE��s�6��ˋk�Q'I����܊�GBEiB���j���QCG�h4Z�D�$ݢY�-R��By%�V+i�T���I|3����4����ĉؙ}���2r����)���Om�fk\]�zH�|�R�iO�l�Mۗ�I6_dْϜf4G��Fk-匷�ݥe�k�\𛍶���V���_�3���X:�-�b(ڴ#ݾ���KĤ����h$�v!VI~}��+s�^����xg��p�h4"�E@�Ӈ$^N������1���	�����ǁ=j��������o��qbZW�?��i�1��wI�t�G��v��e��^3�x޹���k+�t�w��`-;q<3��rJ�r�##���Κr$55G��޶;�a�±c_�ٿΜ�V�{J9�Ԕd��=�(B���}�\�.1�7����׭w�^v�.\�[��"{x<����̣������{�"o���]�|ҵ�"#��[v��n�ٻoޚ>�Mۢ�̛;[�A���(Ks�#�����@�V�s��I������׸��������gn�fV��8\��@�*e	%F��#�n�����8v� �2�Ǎƙ3�2+yV{<6���ܜ����#d9�¡��ȏ ""�z�ז-_�M���^nzjJ�QNk��i�܇��#��~_�Z(_��?���&��2�G9��ɡ�=�gge|�yx�fY$�Q�/R~�'������ll���<����� ~�N�z�����t
s�PVQ��<^�q�s��mOrrJ@�=�t-���K		粲24x6�;�;�%JHJJ
*�|D��-KKMN!p5�olI�x��ݺ�Ge�F��kǏ�H�"A�ռ!i\�xzz�/_�<�R�u�7�u�����U�F��K0��N�rx����̬L�(B���^b���x:y9��}���E������k��%u����QTB��A%DaP	QTB��A%DaP	QTB��A%DaP	QTB��A%DaP	QTB����Blg���    IEND�B`�PK 
     )u�[�G79�  9�                   cirkitFile.jsonPK 
     )u�[                        f�  jsons/PK 
     )u�[�fy�(  �(               ��  jsons/user_defined.jsonPK 
     )u�[                        ��  images/PK 
     )u�[����^� ^� /             ��  images/67df6019-bb76-4308-bacd-6454b246d44a.pngPK 
     )u�[����  �  /             \� images/7de8bea6-aec6-4ad5-83ac-8e47725efc1f.pngPK 
     )u�[�W&��*  �*  /             y� images/b3e67e62-159a-497d-aba3-70fd70f56319.pngPK 
     )u�[�W&��*  �*  /             G� images/ab942d8a-eab6-45a7-8f5a-30ef729b6f10.pngPK 
     )u�[��n GV GV /              images/5a738b76-89aa-4728-b8e5-f09c859dbb14.pngPK 
     )u�[����C   C   /             �b images/ba153158-cccd-4fb1-9320-38bebad1b7f9.pngPK 
     )u�[	��} } /             9� images/bbfae99c-8036-4c5e-89fd-a87441410720.pngPK 
     )u�[d��   �   /             �  images/a262aa33-74c4-460b-b0ad-c746896f6744.pngPK 
     )u�[�c��f  �f  /             p! images/c88b2895-5e8b-4a57-9f9a-b80dd50058b1.pngPK 
     )u�[��EM  M  /             �� images/d3694a2e-5bba-40c3-8069-8db85c4c9209.pngPK      �  8�   